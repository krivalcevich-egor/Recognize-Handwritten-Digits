`timescale 1ns / 1ps 
 
////////////////////////////////////////////////////////////////////////////////// 
// WEIGHT MEMORY (ROM) 
////////////////////////////////////////////////////////////////////////////////// 
module ROM_weights_2 #( 
    parameter int WGHT_INT = 6, // integer part 
    parameter int WGHT_FRC = 16 // fractional part 
)( 
    input logic clk, // clock 
    input logic [9:0] address,
    output [WGHT_INT + WGHT_FRC-1:0] dout 
); 

(* rom_style = "block" *) reg [WGHT_INT + WGHT_FRC-1:0] data;
generate 
  if (WGHT_FRC == 1) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 7'h00; 
        10'b0000000001: data <= 7'h00; 
        10'b0000000010: data <= 7'h00; 
        10'b0000000011: data <= 7'h00; 
        10'b0000000100: data <= 7'h00; 
        10'b0000000101: data <= 7'h00; 
        10'b0000000110: data <= 7'h00; 
        10'b0000000111: data <= 7'h00; 
        10'b0000001000: data <= 7'h00; 
        10'b0000001001: data <= 7'h00; 
        10'b0000001010: data <= 7'h00; 
        10'b0000001011: data <= 7'h00; 
        10'b0000001100: data <= 7'h00; 
        10'b0000001101: data <= 7'h00; 
        10'b0000001110: data <= 7'h00; 
        10'b0000001111: data <= 7'h00; 
        10'b0000010000: data <= 7'h00; 
        10'b0000010001: data <= 7'h00; 
        10'b0000010010: data <= 7'h00; 
        10'b0000010011: data <= 7'h00; 
        10'b0000010100: data <= 7'h00; 
        10'b0000010101: data <= 7'h00; 
        10'b0000010110: data <= 7'h00; 
        10'b0000010111: data <= 7'h00; 
        10'b0000011000: data <= 7'h00; 
        10'b0000011001: data <= 7'h00; 
        10'b0000011010: data <= 7'h00; 
        10'b0000011011: data <= 7'h00; 
        10'b0000011100: data <= 7'h00; 
        10'b0000011101: data <= 7'h00; 
        10'b0000011110: data <= 7'h00; 
        10'b0000011111: data <= 7'h00; 
        10'b0000100000: data <= 7'h00; 
        10'b0000100001: data <= 7'h00; 
        10'b0000100010: data <= 7'h00; 
        10'b0000100011: data <= 7'h00; 
        10'b0000100100: data <= 7'h00; 
        10'b0000100101: data <= 7'h00; 
        10'b0000100110: data <= 7'h00; 
        10'b0000100111: data <= 7'h00; 
        10'b0000101000: data <= 7'h00; 
        10'b0000101001: data <= 7'h00; 
        10'b0000101010: data <= 7'h00; 
        10'b0000101011: data <= 7'h00; 
        10'b0000101100: data <= 7'h00; 
        10'b0000101101: data <= 7'h00; 
        10'b0000101110: data <= 7'h00; 
        10'b0000101111: data <= 7'h00; 
        10'b0000110000: data <= 7'h00; 
        10'b0000110001: data <= 7'h00; 
        10'b0000110010: data <= 7'h00; 
        10'b0000110011: data <= 7'h00; 
        10'b0000110100: data <= 7'h00; 
        10'b0000110101: data <= 7'h00; 
        10'b0000110110: data <= 7'h00; 
        10'b0000110111: data <= 7'h00; 
        10'b0000111000: data <= 7'h00; 
        10'b0000111001: data <= 7'h00; 
        10'b0000111010: data <= 7'h00; 
        10'b0000111011: data <= 7'h00; 
        10'b0000111100: data <= 7'h00; 
        10'b0000111101: data <= 7'h00; 
        10'b0000111110: data <= 7'h00; 
        10'b0000111111: data <= 7'h00; 
        10'b0001000000: data <= 7'h00; 
        10'b0001000001: data <= 7'h00; 
        10'b0001000010: data <= 7'h00; 
        10'b0001000011: data <= 7'h00; 
        10'b0001000100: data <= 7'h00; 
        10'b0001000101: data <= 7'h00; 
        10'b0001000110: data <= 7'h00; 
        10'b0001000111: data <= 7'h00; 
        10'b0001001000: data <= 7'h00; 
        10'b0001001001: data <= 7'h00; 
        10'b0001001010: data <= 7'h00; 
        10'b0001001011: data <= 7'h00; 
        10'b0001001100: data <= 7'h00; 
        10'b0001001101: data <= 7'h00; 
        10'b0001001110: data <= 7'h00; 
        10'b0001001111: data <= 7'h00; 
        10'b0001010000: data <= 7'h00; 
        10'b0001010001: data <= 7'h00; 
        10'b0001010010: data <= 7'h00; 
        10'b0001010011: data <= 7'h00; 
        10'b0001010100: data <= 7'h00; 
        10'b0001010101: data <= 7'h00; 
        10'b0001010110: data <= 7'h00; 
        10'b0001010111: data <= 7'h00; 
        10'b0001011000: data <= 7'h00; 
        10'b0001011001: data <= 7'h00; 
        10'b0001011010: data <= 7'h00; 
        10'b0001011011: data <= 7'h00; 
        10'b0001011100: data <= 7'h00; 
        10'b0001011101: data <= 7'h00; 
        10'b0001011110: data <= 7'h00; 
        10'b0001011111: data <= 7'h00; 
        10'b0001100000: data <= 7'h00; 
        10'b0001100001: data <= 7'h01; 
        10'b0001100010: data <= 7'h00; 
        10'b0001100011: data <= 7'h00; 
        10'b0001100100: data <= 7'h00; 
        10'b0001100101: data <= 7'h00; 
        10'b0001100110: data <= 7'h00; 
        10'b0001100111: data <= 7'h00; 
        10'b0001101000: data <= 7'h00; 
        10'b0001101001: data <= 7'h00; 
        10'b0001101010: data <= 7'h00; 
        10'b0001101011: data <= 7'h00; 
        10'b0001101100: data <= 7'h00; 
        10'b0001101101: data <= 7'h00; 
        10'b0001101110: data <= 7'h00; 
        10'b0001101111: data <= 7'h00; 
        10'b0001110000: data <= 7'h00; 
        10'b0001110001: data <= 7'h00; 
        10'b0001110010: data <= 7'h00; 
        10'b0001110011: data <= 7'h00; 
        10'b0001110100: data <= 7'h00; 
        10'b0001110101: data <= 7'h00; 
        10'b0001110110: data <= 7'h00; 
        10'b0001110111: data <= 7'h00; 
        10'b0001111000: data <= 7'h00; 
        10'b0001111001: data <= 7'h00; 
        10'b0001111010: data <= 7'h00; 
        10'b0001111011: data <= 7'h01; 
        10'b0001111100: data <= 7'h00; 
        10'b0001111101: data <= 7'h00; 
        10'b0001111110: data <= 7'h00; 
        10'b0001111111: data <= 7'h00; 
        10'b0010000000: data <= 7'h00; 
        10'b0010000001: data <= 7'h00; 
        10'b0010000010: data <= 7'h00; 
        10'b0010000011: data <= 7'h00; 
        10'b0010000100: data <= 7'h00; 
        10'b0010000101: data <= 7'h00; 
        10'b0010000110: data <= 7'h00; 
        10'b0010000111: data <= 7'h00; 
        10'b0010001000: data <= 7'h00; 
        10'b0010001001: data <= 7'h00; 
        10'b0010001010: data <= 7'h00; 
        10'b0010001011: data <= 7'h00; 
        10'b0010001100: data <= 7'h00; 
        10'b0010001101: data <= 7'h00; 
        10'b0010001110: data <= 7'h00; 
        10'b0010001111: data <= 7'h00; 
        10'b0010010000: data <= 7'h00; 
        10'b0010010001: data <= 7'h00; 
        10'b0010010010: data <= 7'h00; 
        10'b0010010011: data <= 7'h00; 
        10'b0010010100: data <= 7'h00; 
        10'b0010010101: data <= 7'h01; 
        10'b0010010110: data <= 7'h01; 
        10'b0010010111: data <= 7'h01; 
        10'b0010011000: data <= 7'h01; 
        10'b0010011001: data <= 7'h01; 
        10'b0010011010: data <= 7'h01; 
        10'b0010011011: data <= 7'h01; 
        10'b0010011100: data <= 7'h01; 
        10'b0010011101: data <= 7'h00; 
        10'b0010011110: data <= 7'h00; 
        10'b0010011111: data <= 7'h00; 
        10'b0010100000: data <= 7'h00; 
        10'b0010100001: data <= 7'h00; 
        10'b0010100010: data <= 7'h00; 
        10'b0010100011: data <= 7'h00; 
        10'b0010100100: data <= 7'h00; 
        10'b0010100101: data <= 7'h00; 
        10'b0010100110: data <= 7'h00; 
        10'b0010100111: data <= 7'h00; 
        10'b0010101000: data <= 7'h00; 
        10'b0010101001: data <= 7'h00; 
        10'b0010101010: data <= 7'h00; 
        10'b0010101011: data <= 7'h00; 
        10'b0010101100: data <= 7'h00; 
        10'b0010101101: data <= 7'h00; 
        10'b0010101110: data <= 7'h00; 
        10'b0010101111: data <= 7'h00; 
        10'b0010110000: data <= 7'h00; 
        10'b0010110001: data <= 7'h00; 
        10'b0010110010: data <= 7'h00; 
        10'b0010110011: data <= 7'h00; 
        10'b0010110100: data <= 7'h00; 
        10'b0010110101: data <= 7'h00; 
        10'b0010110110: data <= 7'h00; 
        10'b0010110111: data <= 7'h00; 
        10'b0010111000: data <= 7'h00; 
        10'b0010111001: data <= 7'h00; 
        10'b0010111010: data <= 7'h00; 
        10'b0010111011: data <= 7'h00; 
        10'b0010111100: data <= 7'h00; 
        10'b0010111101: data <= 7'h00; 
        10'b0010111110: data <= 7'h00; 
        10'b0010111111: data <= 7'h00; 
        10'b0011000000: data <= 7'h00; 
        10'b0011000001: data <= 7'h00; 
        10'b0011000010: data <= 7'h00; 
        10'b0011000011: data <= 7'h00; 
        10'b0011000100: data <= 7'h00; 
        10'b0011000101: data <= 7'h00; 
        10'b0011000110: data <= 7'h00; 
        10'b0011000111: data <= 7'h00; 
        10'b0011001000: data <= 7'h00; 
        10'b0011001001: data <= 7'h00; 
        10'b0011001010: data <= 7'h00; 
        10'b0011001011: data <= 7'h00; 
        10'b0011001100: data <= 7'h00; 
        10'b0011001101: data <= 7'h00; 
        10'b0011001110: data <= 7'h00; 
        10'b0011001111: data <= 7'h00; 
        10'b0011010000: data <= 7'h00; 
        10'b0011010001: data <= 7'h00; 
        10'b0011010010: data <= 7'h00; 
        10'b0011010011: data <= 7'h00; 
        10'b0011010100: data <= 7'h00; 
        10'b0011010101: data <= 7'h00; 
        10'b0011010110: data <= 7'h00; 
        10'b0011010111: data <= 7'h00; 
        10'b0011011000: data <= 7'h00; 
        10'b0011011001: data <= 7'h00; 
        10'b0011011010: data <= 7'h00; 
        10'b0011011011: data <= 7'h00; 
        10'b0011011100: data <= 7'h00; 
        10'b0011011101: data <= 7'h00; 
        10'b0011011110: data <= 7'h00; 
        10'b0011011111: data <= 7'h00; 
        10'b0011100000: data <= 7'h00; 
        10'b0011100001: data <= 7'h00; 
        10'b0011100010: data <= 7'h00; 
        10'b0011100011: data <= 7'h00; 
        10'b0011100100: data <= 7'h00; 
        10'b0011100101: data <= 7'h00; 
        10'b0011100110: data <= 7'h00; 
        10'b0011100111: data <= 7'h00; 
        10'b0011101000: data <= 7'h00; 
        10'b0011101001: data <= 7'h00; 
        10'b0011101010: data <= 7'h00; 
        10'b0011101011: data <= 7'h00; 
        10'b0011101100: data <= 7'h00; 
        10'b0011101101: data <= 7'h00; 
        10'b0011101110: data <= 7'h00; 
        10'b0011101111: data <= 7'h00; 
        10'b0011110000: data <= 7'h00; 
        10'b0011110001: data <= 7'h00; 
        10'b0011110010: data <= 7'h00; 
        10'b0011110011: data <= 7'h00; 
        10'b0011110100: data <= 7'h00; 
        10'b0011110101: data <= 7'h00; 
        10'b0011110110: data <= 7'h00; 
        10'b0011110111: data <= 7'h00; 
        10'b0011111000: data <= 7'h00; 
        10'b0011111001: data <= 7'h00; 
        10'b0011111010: data <= 7'h00; 
        10'b0011111011: data <= 7'h00; 
        10'b0011111100: data <= 7'h00; 
        10'b0011111101: data <= 7'h00; 
        10'b0011111110: data <= 7'h00; 
        10'b0011111111: data <= 7'h00; 
        10'b0100000000: data <= 7'h00; 
        10'b0100000001: data <= 7'h00; 
        10'b0100000010: data <= 7'h00; 
        10'b0100000011: data <= 7'h00; 
        10'b0100000100: data <= 7'h00; 
        10'b0100000101: data <= 7'h00; 
        10'b0100000110: data <= 7'h00; 
        10'b0100000111: data <= 7'h00; 
        10'b0100001000: data <= 7'h00; 
        10'b0100001001: data <= 7'h00; 
        10'b0100001010: data <= 7'h00; 
        10'b0100001011: data <= 7'h00; 
        10'b0100001100: data <= 7'h00; 
        10'b0100001101: data <= 7'h00; 
        10'b0100001110: data <= 7'h00; 
        10'b0100001111: data <= 7'h00; 
        10'b0100010000: data <= 7'h00; 
        10'b0100010001: data <= 7'h00; 
        10'b0100010010: data <= 7'h00; 
        10'b0100010011: data <= 7'h00; 
        10'b0100010100: data <= 7'h00; 
        10'b0100010101: data <= 7'h00; 
        10'b0100010110: data <= 7'h00; 
        10'b0100010111: data <= 7'h00; 
        10'b0100011000: data <= 7'h00; 
        10'b0100011001: data <= 7'h00; 
        10'b0100011010: data <= 7'h00; 
        10'b0100011011: data <= 7'h00; 
        10'b0100011100: data <= 7'h00; 
        10'b0100011101: data <= 7'h00; 
        10'b0100011110: data <= 7'h00; 
        10'b0100011111: data <= 7'h00; 
        10'b0100100000: data <= 7'h00; 
        10'b0100100001: data <= 7'h00; 
        10'b0100100010: data <= 7'h7f; 
        10'b0100100011: data <= 7'h7f; 
        10'b0100100100: data <= 7'h7f; 
        10'b0100100101: data <= 7'h7f; 
        10'b0100100110: data <= 7'h00; 
        10'b0100100111: data <= 7'h00; 
        10'b0100101000: data <= 7'h00; 
        10'b0100101001: data <= 7'h00; 
        10'b0100101010: data <= 7'h00; 
        10'b0100101011: data <= 7'h00; 
        10'b0100101100: data <= 7'h00; 
        10'b0100101101: data <= 7'h00; 
        10'b0100101110: data <= 7'h00; 
        10'b0100101111: data <= 7'h00; 
        10'b0100110000: data <= 7'h00; 
        10'b0100110001: data <= 7'h00; 
        10'b0100110010: data <= 7'h00; 
        10'b0100110011: data <= 7'h00; 
        10'b0100110100: data <= 7'h00; 
        10'b0100110101: data <= 7'h00; 
        10'b0100110110: data <= 7'h00; 
        10'b0100110111: data <= 7'h00; 
        10'b0100111000: data <= 7'h00; 
        10'b0100111001: data <= 7'h00; 
        10'b0100111010: data <= 7'h7f; 
        10'b0100111011: data <= 7'h7f; 
        10'b0100111100: data <= 7'h7f; 
        10'b0100111101: data <= 7'h7f; 
        10'b0100111110: data <= 7'h7f; 
        10'b0100111111: data <= 7'h7f; 
        10'b0101000000: data <= 7'h7f; 
        10'b0101000001: data <= 7'h7f; 
        10'b0101000010: data <= 7'h7f; 
        10'b0101000011: data <= 7'h00; 
        10'b0101000100: data <= 7'h00; 
        10'b0101000101: data <= 7'h00; 
        10'b0101000110: data <= 7'h00; 
        10'b0101000111: data <= 7'h00; 
        10'b0101001000: data <= 7'h00; 
        10'b0101001001: data <= 7'h00; 
        10'b0101001010: data <= 7'h00; 
        10'b0101001011: data <= 7'h00; 
        10'b0101001100: data <= 7'h00; 
        10'b0101001101: data <= 7'h00; 
        10'b0101001110: data <= 7'h00; 
        10'b0101001111: data <= 7'h00; 
        10'b0101010000: data <= 7'h00; 
        10'b0101010001: data <= 7'h00; 
        10'b0101010010: data <= 7'h00; 
        10'b0101010011: data <= 7'h00; 
        10'b0101010100: data <= 7'h00; 
        10'b0101010101: data <= 7'h7f; 
        10'b0101010110: data <= 7'h7f; 
        10'b0101010111: data <= 7'h7f; 
        10'b0101011000: data <= 7'h7f; 
        10'b0101011001: data <= 7'h7f; 
        10'b0101011010: data <= 7'h7f; 
        10'b0101011011: data <= 7'h7f; 
        10'b0101011100: data <= 7'h7f; 
        10'b0101011101: data <= 7'h7f; 
        10'b0101011110: data <= 7'h7f; 
        10'b0101011111: data <= 7'h7f; 
        10'b0101100000: data <= 7'h00; 
        10'b0101100001: data <= 7'h00; 
        10'b0101100010: data <= 7'h00; 
        10'b0101100011: data <= 7'h00; 
        10'b0101100100: data <= 7'h00; 
        10'b0101100101: data <= 7'h00; 
        10'b0101100110: data <= 7'h00; 
        10'b0101100111: data <= 7'h00; 
        10'b0101101000: data <= 7'h00; 
        10'b0101101001: data <= 7'h00; 
        10'b0101101010: data <= 7'h00; 
        10'b0101101011: data <= 7'h00; 
        10'b0101101100: data <= 7'h00; 
        10'b0101101101: data <= 7'h00; 
        10'b0101101110: data <= 7'h00; 
        10'b0101101111: data <= 7'h00; 
        10'b0101110000: data <= 7'h00; 
        10'b0101110001: data <= 7'h7f; 
        10'b0101110010: data <= 7'h7f; 
        10'b0101110011: data <= 7'h7f; 
        10'b0101110100: data <= 7'h7f; 
        10'b0101110101: data <= 7'h7f; 
        10'b0101110110: data <= 7'h7f; 
        10'b0101110111: data <= 7'h00; 
        10'b0101111000: data <= 7'h00; 
        10'b0101111001: data <= 7'h00; 
        10'b0101111010: data <= 7'h00; 
        10'b0101111011: data <= 7'h00; 
        10'b0101111100: data <= 7'h7f; 
        10'b0101111101: data <= 7'h00; 
        10'b0101111110: data <= 7'h00; 
        10'b0101111111: data <= 7'h00; 
        10'b0110000000: data <= 7'h00; 
        10'b0110000001: data <= 7'h00; 
        10'b0110000010: data <= 7'h00; 
        10'b0110000011: data <= 7'h00; 
        10'b0110000100: data <= 7'h00; 
        10'b0110000101: data <= 7'h00; 
        10'b0110000110: data <= 7'h00; 
        10'b0110000111: data <= 7'h00; 
        10'b0110001000: data <= 7'h00; 
        10'b0110001001: data <= 7'h00; 
        10'b0110001010: data <= 7'h00; 
        10'b0110001011: data <= 7'h00; 
        10'b0110001100: data <= 7'h00; 
        10'b0110001101: data <= 7'h7f; 
        10'b0110001110: data <= 7'h7f; 
        10'b0110001111: data <= 7'h7f; 
        10'b0110010000: data <= 7'h00; 
        10'b0110010001: data <= 7'h00; 
        10'b0110010010: data <= 7'h00; 
        10'b0110010011: data <= 7'h00; 
        10'b0110010100: data <= 7'h00; 
        10'b0110010101: data <= 7'h00; 
        10'b0110010110: data <= 7'h00; 
        10'b0110010111: data <= 7'h00; 
        10'b0110011000: data <= 7'h00; 
        10'b0110011001: data <= 7'h00; 
        10'b0110011010: data <= 7'h00; 
        10'b0110011011: data <= 7'h00; 
        10'b0110011100: data <= 7'h00; 
        10'b0110011101: data <= 7'h00; 
        10'b0110011110: data <= 7'h00; 
        10'b0110011111: data <= 7'h00; 
        10'b0110100000: data <= 7'h00; 
        10'b0110100001: data <= 7'h00; 
        10'b0110100010: data <= 7'h00; 
        10'b0110100011: data <= 7'h00; 
        10'b0110100100: data <= 7'h00; 
        10'b0110100101: data <= 7'h00; 
        10'b0110100110: data <= 7'h00; 
        10'b0110100111: data <= 7'h00; 
        10'b0110101000: data <= 7'h00; 
        10'b0110101001: data <= 7'h00; 
        10'b0110101010: data <= 7'h00; 
        10'b0110101011: data <= 7'h00; 
        10'b0110101100: data <= 7'h00; 
        10'b0110101101: data <= 7'h00; 
        10'b0110101110: data <= 7'h00; 
        10'b0110101111: data <= 7'h00; 
        10'b0110110000: data <= 7'h00; 
        10'b0110110001: data <= 7'h00; 
        10'b0110110010: data <= 7'h00; 
        10'b0110110011: data <= 7'h00; 
        10'b0110110100: data <= 7'h00; 
        10'b0110110101: data <= 7'h00; 
        10'b0110110110: data <= 7'h00; 
        10'b0110110111: data <= 7'h00; 
        10'b0110111000: data <= 7'h00; 
        10'b0110111001: data <= 7'h00; 
        10'b0110111010: data <= 7'h00; 
        10'b0110111011: data <= 7'h00; 
        10'b0110111100: data <= 7'h00; 
        10'b0110111101: data <= 7'h00; 
        10'b0110111110: data <= 7'h00; 
        10'b0110111111: data <= 7'h00; 
        10'b0111000000: data <= 7'h00; 
        10'b0111000001: data <= 7'h00; 
        10'b0111000010: data <= 7'h00; 
        10'b0111000011: data <= 7'h00; 
        10'b0111000100: data <= 7'h00; 
        10'b0111000101: data <= 7'h00; 
        10'b0111000110: data <= 7'h00; 
        10'b0111000111: data <= 7'h00; 
        10'b0111001000: data <= 7'h00; 
        10'b0111001001: data <= 7'h00; 
        10'b0111001010: data <= 7'h00; 
        10'b0111001011: data <= 7'h00; 
        10'b0111001100: data <= 7'h00; 
        10'b0111001101: data <= 7'h00; 
        10'b0111001110: data <= 7'h00; 
        10'b0111001111: data <= 7'h00; 
        10'b0111010000: data <= 7'h00; 
        10'b0111010001: data <= 7'h00; 
        10'b0111010010: data <= 7'h00; 
        10'b0111010011: data <= 7'h00; 
        10'b0111010100: data <= 7'h00; 
        10'b0111010101: data <= 7'h00; 
        10'b0111010110: data <= 7'h00; 
        10'b0111010111: data <= 7'h00; 
        10'b0111011000: data <= 7'h00; 
        10'b0111011001: data <= 7'h00; 
        10'b0111011010: data <= 7'h00; 
        10'b0111011011: data <= 7'h00; 
        10'b0111011100: data <= 7'h00; 
        10'b0111011101: data <= 7'h00; 
        10'b0111011110: data <= 7'h00; 
        10'b0111011111: data <= 7'h00; 
        10'b0111100000: data <= 7'h00; 
        10'b0111100001: data <= 7'h01; 
        10'b0111100010: data <= 7'h01; 
        10'b0111100011: data <= 7'h00; 
        10'b0111100100: data <= 7'h00; 
        10'b0111100101: data <= 7'h00; 
        10'b0111100110: data <= 7'h01; 
        10'b0111100111: data <= 7'h00; 
        10'b0111101000: data <= 7'h00; 
        10'b0111101001: data <= 7'h00; 
        10'b0111101010: data <= 7'h00; 
        10'b0111101011: data <= 7'h00; 
        10'b0111101100: data <= 7'h00; 
        10'b0111101101: data <= 7'h00; 
        10'b0111101110: data <= 7'h00; 
        10'b0111101111: data <= 7'h00; 
        10'b0111110000: data <= 7'h00; 
        10'b0111110001: data <= 7'h00; 
        10'b0111110010: data <= 7'h00; 
        10'b0111110011: data <= 7'h00; 
        10'b0111110100: data <= 7'h01; 
        10'b0111110101: data <= 7'h01; 
        10'b0111110110: data <= 7'h00; 
        10'b0111110111: data <= 7'h00; 
        10'b0111111000: data <= 7'h00; 
        10'b0111111001: data <= 7'h00; 
        10'b0111111010: data <= 7'h00; 
        10'b0111111011: data <= 7'h00; 
        10'b0111111100: data <= 7'h00; 
        10'b0111111101: data <= 7'h01; 
        10'b0111111110: data <= 7'h01; 
        10'b0111111111: data <= 7'h01; 
        10'b1000000000: data <= 7'h00; 
        10'b1000000001: data <= 7'h00; 
        10'b1000000010: data <= 7'h01; 
        10'b1000000011: data <= 7'h01; 
        10'b1000000100: data <= 7'h01; 
        10'b1000000101: data <= 7'h01; 
        10'b1000000110: data <= 7'h01; 
        10'b1000000111: data <= 7'h00; 
        10'b1000001000: data <= 7'h00; 
        10'b1000001001: data <= 7'h00; 
        10'b1000001010: data <= 7'h00; 
        10'b1000001011: data <= 7'h00; 
        10'b1000001100: data <= 7'h00; 
        10'b1000001101: data <= 7'h00; 
        10'b1000001110: data <= 7'h00; 
        10'b1000001111: data <= 7'h01; 
        10'b1000010000: data <= 7'h01; 
        10'b1000010001: data <= 7'h00; 
        10'b1000010010: data <= 7'h00; 
        10'b1000010011: data <= 7'h00; 
        10'b1000010100: data <= 7'h00; 
        10'b1000010101: data <= 7'h00; 
        10'b1000010110: data <= 7'h00; 
        10'b1000010111: data <= 7'h00; 
        10'b1000011000: data <= 7'h00; 
        10'b1000011001: data <= 7'h01; 
        10'b1000011010: data <= 7'h01; 
        10'b1000011011: data <= 7'h01; 
        10'b1000011100: data <= 7'h01; 
        10'b1000011101: data <= 7'h01; 
        10'b1000011110: data <= 7'h01; 
        10'b1000011111: data <= 7'h01; 
        10'b1000100000: data <= 7'h01; 
        10'b1000100001: data <= 7'h00; 
        10'b1000100010: data <= 7'h00; 
        10'b1000100011: data <= 7'h00; 
        10'b1000100100: data <= 7'h00; 
        10'b1000100101: data <= 7'h00; 
        10'b1000100110: data <= 7'h00; 
        10'b1000100111: data <= 7'h00; 
        10'b1000101000: data <= 7'h00; 
        10'b1000101001: data <= 7'h00; 
        10'b1000101010: data <= 7'h01; 
        10'b1000101011: data <= 7'h01; 
        10'b1000101100: data <= 7'h00; 
        10'b1000101101: data <= 7'h00; 
        10'b1000101110: data <= 7'h00; 
        10'b1000101111: data <= 7'h00; 
        10'b1000110000: data <= 7'h00; 
        10'b1000110001: data <= 7'h00; 
        10'b1000110010: data <= 7'h00; 
        10'b1000110011: data <= 7'h00; 
        10'b1000110100: data <= 7'h00; 
        10'b1000110101: data <= 7'h00; 
        10'b1000110110: data <= 7'h00; 
        10'b1000110111: data <= 7'h01; 
        10'b1000111000: data <= 7'h01; 
        10'b1000111001: data <= 7'h00; 
        10'b1000111010: data <= 7'h00; 
        10'b1000111011: data <= 7'h01; 
        10'b1000111100: data <= 7'h00; 
        10'b1000111101: data <= 7'h00; 
        10'b1000111110: data <= 7'h00; 
        10'b1000111111: data <= 7'h00; 
        10'b1001000000: data <= 7'h00; 
        10'b1001000001: data <= 7'h00; 
        10'b1001000010: data <= 7'h00; 
        10'b1001000011: data <= 7'h00; 
        10'b1001000100: data <= 7'h00; 
        10'b1001000101: data <= 7'h00; 
        10'b1001000110: data <= 7'h01; 
        10'b1001000111: data <= 7'h01; 
        10'b1001001000: data <= 7'h00; 
        10'b1001001001: data <= 7'h00; 
        10'b1001001010: data <= 7'h00; 
        10'b1001001011: data <= 7'h00; 
        10'b1001001100: data <= 7'h00; 
        10'b1001001101: data <= 7'h00; 
        10'b1001001110: data <= 7'h00; 
        10'b1001001111: data <= 7'h00; 
        10'b1001010000: data <= 7'h00; 
        10'b1001010001: data <= 7'h00; 
        10'b1001010010: data <= 7'h00; 
        10'b1001010011: data <= 7'h00; 
        10'b1001010100: data <= 7'h00; 
        10'b1001010101: data <= 7'h00; 
        10'b1001010110: data <= 7'h00; 
        10'b1001010111: data <= 7'h00; 
        10'b1001011000: data <= 7'h00; 
        10'b1001011001: data <= 7'h00; 
        10'b1001011010: data <= 7'h00; 
        10'b1001011011: data <= 7'h00; 
        10'b1001011100: data <= 7'h00; 
        10'b1001011101: data <= 7'h00; 
        10'b1001011110: data <= 7'h00; 
        10'b1001011111: data <= 7'h00; 
        10'b1001100000: data <= 7'h00; 
        10'b1001100001: data <= 7'h00; 
        10'b1001100010: data <= 7'h01; 
        10'b1001100011: data <= 7'h01; 
        10'b1001100100: data <= 7'h00; 
        10'b1001100101: data <= 7'h00; 
        10'b1001100110: data <= 7'h00; 
        10'b1001100111: data <= 7'h00; 
        10'b1001101000: data <= 7'h00; 
        10'b1001101001: data <= 7'h00; 
        10'b1001101010: data <= 7'h00; 
        10'b1001101011: data <= 7'h00; 
        10'b1001101100: data <= 7'h00; 
        10'b1001101101: data <= 7'h00; 
        10'b1001101110: data <= 7'h00; 
        10'b1001101111: data <= 7'h00; 
        10'b1001110000: data <= 7'h00; 
        10'b1001110001: data <= 7'h00; 
        10'b1001110010: data <= 7'h00; 
        10'b1001110011: data <= 7'h00; 
        10'b1001110100: data <= 7'h00; 
        10'b1001110101: data <= 7'h00; 
        10'b1001110110: data <= 7'h00; 
        10'b1001110111: data <= 7'h00; 
        10'b1001111000: data <= 7'h00; 
        10'b1001111001: data <= 7'h00; 
        10'b1001111010: data <= 7'h00; 
        10'b1001111011: data <= 7'h00; 
        10'b1001111100: data <= 7'h00; 
        10'b1001111101: data <= 7'h00; 
        10'b1001111110: data <= 7'h00; 
        10'b1001111111: data <= 7'h00; 
        10'b1010000000: data <= 7'h00; 
        10'b1010000001: data <= 7'h00; 
        10'b1010000010: data <= 7'h00; 
        10'b1010000011: data <= 7'h00; 
        10'b1010000100: data <= 7'h00; 
        10'b1010000101: data <= 7'h00; 
        10'b1010000110: data <= 7'h00; 
        10'b1010000111: data <= 7'h00; 
        10'b1010001000: data <= 7'h00; 
        10'b1010001001: data <= 7'h00; 
        10'b1010001010: data <= 7'h00; 
        10'b1010001011: data <= 7'h00; 
        10'b1010001100: data <= 7'h00; 
        10'b1010001101: data <= 7'h00; 
        10'b1010001110: data <= 7'h00; 
        10'b1010001111: data <= 7'h00; 
        10'b1010010000: data <= 7'h00; 
        10'b1010010001: data <= 7'h00; 
        10'b1010010010: data <= 7'h00; 
        10'b1010010011: data <= 7'h00; 
        10'b1010010100: data <= 7'h00; 
        10'b1010010101: data <= 7'h00; 
        10'b1010010110: data <= 7'h00; 
        10'b1010010111: data <= 7'h00; 
        10'b1010011000: data <= 7'h00; 
        10'b1010011001: data <= 7'h00; 
        10'b1010011010: data <= 7'h00; 
        10'b1010011011: data <= 7'h00; 
        10'b1010011100: data <= 7'h00; 
        10'b1010011101: data <= 7'h00; 
        10'b1010011110: data <= 7'h00; 
        10'b1010011111: data <= 7'h00; 
        10'b1010100000: data <= 7'h00; 
        10'b1010100001: data <= 7'h00; 
        10'b1010100010: data <= 7'h00; 
        10'b1010100011: data <= 7'h00; 
        10'b1010100100: data <= 7'h00; 
        10'b1010100101: data <= 7'h00; 
        10'b1010100110: data <= 7'h00; 
        10'b1010100111: data <= 7'h00; 
        10'b1010101000: data <= 7'h00; 
        10'b1010101001: data <= 7'h00; 
        10'b1010101010: data <= 7'h00; 
        10'b1010101011: data <= 7'h00; 
        10'b1010101100: data <= 7'h00; 
        10'b1010101101: data <= 7'h00; 
        10'b1010101110: data <= 7'h00; 
        10'b1010101111: data <= 7'h00; 
        10'b1010110000: data <= 7'h00; 
        10'b1010110001: data <= 7'h00; 
        10'b1010110010: data <= 7'h00; 
        10'b1010110011: data <= 7'h00; 
        10'b1010110100: data <= 7'h00; 
        10'b1010110101: data <= 7'h00; 
        10'b1010110110: data <= 7'h00; 
        10'b1010110111: data <= 7'h00; 
        10'b1010111000: data <= 7'h00; 
        10'b1010111001: data <= 7'h00; 
        10'b1010111010: data <= 7'h00; 
        10'b1010111011: data <= 7'h00; 
        10'b1010111100: data <= 7'h00; 
        10'b1010111101: data <= 7'h00; 
        10'b1010111110: data <= 7'h00; 
        10'b1010111111: data <= 7'h00; 
        10'b1011000000: data <= 7'h00; 
        10'b1011000001: data <= 7'h00; 
        10'b1011000010: data <= 7'h00; 
        10'b1011000011: data <= 7'h00; 
        10'b1011000100: data <= 7'h00; 
        10'b1011000101: data <= 7'h00; 
        10'b1011000110: data <= 7'h00; 
        10'b1011000111: data <= 7'h00; 
        10'b1011001000: data <= 7'h00; 
        10'b1011001001: data <= 7'h00; 
        10'b1011001010: data <= 7'h00; 
        10'b1011001011: data <= 7'h00; 
        10'b1011001100: data <= 7'h00; 
        10'b1011001101: data <= 7'h00; 
        10'b1011001110: data <= 7'h00; 
        10'b1011001111: data <= 7'h00; 
        10'b1011010000: data <= 7'h00; 
        10'b1011010001: data <= 7'h00; 
        10'b1011010010: data <= 7'h00; 
        10'b1011010011: data <= 7'h00; 
        10'b1011010100: data <= 7'h00; 
        10'b1011010101: data <= 7'h00; 
        10'b1011010110: data <= 7'h00; 
        10'b1011010111: data <= 7'h00; 
        10'b1011011000: data <= 7'h00; 
        10'b1011011001: data <= 7'h00; 
        10'b1011011010: data <= 7'h00; 
        10'b1011011011: data <= 7'h00; 
        10'b1011011100: data <= 7'h00; 
        10'b1011011101: data <= 7'h00; 
        10'b1011011110: data <= 7'h00; 
        10'b1011011111: data <= 7'h00; 
        10'b1011100000: data <= 7'h00; 
        10'b1011100001: data <= 7'h00; 
        10'b1011100010: data <= 7'h00; 
        10'b1011100011: data <= 7'h00; 
        10'b1011100100: data <= 7'h00; 
        10'b1011100101: data <= 7'h00; 
        10'b1011100110: data <= 7'h00; 
        10'b1011100111: data <= 7'h00; 
        10'b1011101000: data <= 7'h00; 
        10'b1011101001: data <= 7'h00; 
        10'b1011101010: data <= 7'h00; 
        10'b1011101011: data <= 7'h00; 
        10'b1011101100: data <= 7'h00; 
        10'b1011101101: data <= 7'h00; 
        10'b1011101110: data <= 7'h00; 
        10'b1011101111: data <= 7'h00; 
        10'b1011110000: data <= 7'h00; 
        10'b1011110001: data <= 7'h00; 
        10'b1011110010: data <= 7'h00; 
        10'b1011110011: data <= 7'h00; 
        10'b1011110100: data <= 7'h00; 
        10'b1011110101: data <= 7'h00; 
        10'b1011110110: data <= 7'h00; 
        10'b1011110111: data <= 7'h00; 
        10'b1011111000: data <= 7'h00; 
        10'b1011111001: data <= 7'h00; 
        10'b1011111010: data <= 7'h00; 
        10'b1011111011: data <= 7'h00; 
        10'b1011111100: data <= 7'h00; 
        10'b1011111101: data <= 7'h00; 
        10'b1011111110: data <= 7'h00; 
        10'b1011111111: data <= 7'h00; 
        10'b1100000000: data <= 7'h00; 
        10'b1100000001: data <= 7'h00; 
        10'b1100000010: data <= 7'h00; 
        10'b1100000011: data <= 7'h00; 
        10'b1100000100: data <= 7'h00; 
        10'b1100000101: data <= 7'h00; 
        10'b1100000110: data <= 7'h00; 
        10'b1100000111: data <= 7'h00; 
        10'b1100001000: data <= 7'h00; 
        10'b1100001001: data <= 7'h00; 
        10'b1100001010: data <= 7'h00; 
        10'b1100001011: data <= 7'h00; 
        10'b1100001100: data <= 7'h00; 
        10'b1100001101: data <= 7'h00; 
        10'b1100001110: data <= 7'h00; 
        10'b1100001111: data <= 7'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 2) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 8'h00; 
        10'b0000000001: data <= 8'h00; 
        10'b0000000010: data <= 8'h00; 
        10'b0000000011: data <= 8'h00; 
        10'b0000000100: data <= 8'h00; 
        10'b0000000101: data <= 8'h00; 
        10'b0000000110: data <= 8'h00; 
        10'b0000000111: data <= 8'h00; 
        10'b0000001000: data <= 8'h00; 
        10'b0000001001: data <= 8'h00; 
        10'b0000001010: data <= 8'h00; 
        10'b0000001011: data <= 8'h00; 
        10'b0000001100: data <= 8'h00; 
        10'b0000001101: data <= 8'h00; 
        10'b0000001110: data <= 8'h00; 
        10'b0000001111: data <= 8'h00; 
        10'b0000010000: data <= 8'h00; 
        10'b0000010001: data <= 8'h00; 
        10'b0000010010: data <= 8'h00; 
        10'b0000010011: data <= 8'h00; 
        10'b0000010100: data <= 8'h00; 
        10'b0000010101: data <= 8'h00; 
        10'b0000010110: data <= 8'h00; 
        10'b0000010111: data <= 8'h00; 
        10'b0000011000: data <= 8'h00; 
        10'b0000011001: data <= 8'h00; 
        10'b0000011010: data <= 8'h00; 
        10'b0000011011: data <= 8'h00; 
        10'b0000011100: data <= 8'h00; 
        10'b0000011101: data <= 8'h00; 
        10'b0000011110: data <= 8'h00; 
        10'b0000011111: data <= 8'h00; 
        10'b0000100000: data <= 8'h00; 
        10'b0000100001: data <= 8'h00; 
        10'b0000100010: data <= 8'h00; 
        10'b0000100011: data <= 8'h00; 
        10'b0000100100: data <= 8'h00; 
        10'b0000100101: data <= 8'h00; 
        10'b0000100110: data <= 8'h00; 
        10'b0000100111: data <= 8'h00; 
        10'b0000101000: data <= 8'h00; 
        10'b0000101001: data <= 8'h00; 
        10'b0000101010: data <= 8'h00; 
        10'b0000101011: data <= 8'h00; 
        10'b0000101100: data <= 8'h00; 
        10'b0000101101: data <= 8'h00; 
        10'b0000101110: data <= 8'h00; 
        10'b0000101111: data <= 8'h00; 
        10'b0000110000: data <= 8'h00; 
        10'b0000110001: data <= 8'h00; 
        10'b0000110010: data <= 8'h00; 
        10'b0000110011: data <= 8'h00; 
        10'b0000110100: data <= 8'h00; 
        10'b0000110101: data <= 8'h00; 
        10'b0000110110: data <= 8'h00; 
        10'b0000110111: data <= 8'h00; 
        10'b0000111000: data <= 8'h00; 
        10'b0000111001: data <= 8'h00; 
        10'b0000111010: data <= 8'h00; 
        10'b0000111011: data <= 8'h00; 
        10'b0000111100: data <= 8'h00; 
        10'b0000111101: data <= 8'h00; 
        10'b0000111110: data <= 8'h00; 
        10'b0000111111: data <= 8'h00; 
        10'b0001000000: data <= 8'h00; 
        10'b0001000001: data <= 8'h00; 
        10'b0001000010: data <= 8'h00; 
        10'b0001000011: data <= 8'h00; 
        10'b0001000100: data <= 8'h00; 
        10'b0001000101: data <= 8'h00; 
        10'b0001000110: data <= 8'h00; 
        10'b0001000111: data <= 8'h00; 
        10'b0001001000: data <= 8'h00; 
        10'b0001001001: data <= 8'h00; 
        10'b0001001010: data <= 8'h00; 
        10'b0001001011: data <= 8'h00; 
        10'b0001001100: data <= 8'h00; 
        10'b0001001101: data <= 8'h00; 
        10'b0001001110: data <= 8'h00; 
        10'b0001001111: data <= 8'h00; 
        10'b0001010000: data <= 8'h00; 
        10'b0001010001: data <= 8'h00; 
        10'b0001010010: data <= 8'h00; 
        10'b0001010011: data <= 8'h00; 
        10'b0001010100: data <= 8'h00; 
        10'b0001010101: data <= 8'h00; 
        10'b0001010110: data <= 8'h00; 
        10'b0001010111: data <= 8'h00; 
        10'b0001011000: data <= 8'h00; 
        10'b0001011001: data <= 8'h00; 
        10'b0001011010: data <= 8'h00; 
        10'b0001011011: data <= 8'h00; 
        10'b0001011100: data <= 8'h00; 
        10'b0001011101: data <= 8'h00; 
        10'b0001011110: data <= 8'h01; 
        10'b0001011111: data <= 8'h01; 
        10'b0001100000: data <= 8'h01; 
        10'b0001100001: data <= 8'h01; 
        10'b0001100010: data <= 8'h01; 
        10'b0001100011: data <= 8'h00; 
        10'b0001100100: data <= 8'h00; 
        10'b0001100101: data <= 8'h00; 
        10'b0001100110: data <= 8'h00; 
        10'b0001100111: data <= 8'h00; 
        10'b0001101000: data <= 8'h00; 
        10'b0001101001: data <= 8'h00; 
        10'b0001101010: data <= 8'h00; 
        10'b0001101011: data <= 8'h00; 
        10'b0001101100: data <= 8'h00; 
        10'b0001101101: data <= 8'h00; 
        10'b0001101110: data <= 8'h00; 
        10'b0001101111: data <= 8'h00; 
        10'b0001110000: data <= 8'h00; 
        10'b0001110001: data <= 8'h00; 
        10'b0001110010: data <= 8'h00; 
        10'b0001110011: data <= 8'h00; 
        10'b0001110100: data <= 8'h00; 
        10'b0001110101: data <= 8'h00; 
        10'b0001110110: data <= 8'h00; 
        10'b0001110111: data <= 8'h00; 
        10'b0001111000: data <= 8'h00; 
        10'b0001111001: data <= 8'h01; 
        10'b0001111010: data <= 8'h01; 
        10'b0001111011: data <= 8'h01; 
        10'b0001111100: data <= 8'h01; 
        10'b0001111101: data <= 8'h01; 
        10'b0001111110: data <= 8'h01; 
        10'b0001111111: data <= 8'h00; 
        10'b0010000000: data <= 8'h00; 
        10'b0010000001: data <= 8'h00; 
        10'b0010000010: data <= 8'h00; 
        10'b0010000011: data <= 8'h00; 
        10'b0010000100: data <= 8'h00; 
        10'b0010000101: data <= 8'h00; 
        10'b0010000110: data <= 8'hff; 
        10'b0010000111: data <= 8'hff; 
        10'b0010001000: data <= 8'h00; 
        10'b0010001001: data <= 8'h00; 
        10'b0010001010: data <= 8'h00; 
        10'b0010001011: data <= 8'h00; 
        10'b0010001100: data <= 8'h00; 
        10'b0010001101: data <= 8'h00; 
        10'b0010001110: data <= 8'h00; 
        10'b0010001111: data <= 8'h00; 
        10'b0010010000: data <= 8'h00; 
        10'b0010010001: data <= 8'h00; 
        10'b0010010010: data <= 8'h00; 
        10'b0010010011: data <= 8'h00; 
        10'b0010010100: data <= 8'h01; 
        10'b0010010101: data <= 8'h01; 
        10'b0010010110: data <= 8'h01; 
        10'b0010010111: data <= 8'h01; 
        10'b0010011000: data <= 8'h01; 
        10'b0010011001: data <= 8'h01; 
        10'b0010011010: data <= 8'h01; 
        10'b0010011011: data <= 8'h01; 
        10'b0010011100: data <= 8'h01; 
        10'b0010011101: data <= 8'h01; 
        10'b0010011110: data <= 8'h01; 
        10'b0010011111: data <= 8'h00; 
        10'b0010100000: data <= 8'h00; 
        10'b0010100001: data <= 8'h00; 
        10'b0010100010: data <= 8'h00; 
        10'b0010100011: data <= 8'hff; 
        10'b0010100100: data <= 8'h00; 
        10'b0010100101: data <= 8'h00; 
        10'b0010100110: data <= 8'h00; 
        10'b0010100111: data <= 8'h00; 
        10'b0010101000: data <= 8'h00; 
        10'b0010101001: data <= 8'h00; 
        10'b0010101010: data <= 8'h00; 
        10'b0010101011: data <= 8'h00; 
        10'b0010101100: data <= 8'h00; 
        10'b0010101101: data <= 8'h00; 
        10'b0010101110: data <= 8'h00; 
        10'b0010101111: data <= 8'h01; 
        10'b0010110000: data <= 8'h01; 
        10'b0010110001: data <= 8'h01; 
        10'b0010110010: data <= 8'h01; 
        10'b0010110011: data <= 8'h01; 
        10'b0010110100: data <= 8'h01; 
        10'b0010110101: data <= 8'h01; 
        10'b0010110110: data <= 8'h01; 
        10'b0010110111: data <= 8'h00; 
        10'b0010111000: data <= 8'h00; 
        10'b0010111001: data <= 8'h00; 
        10'b0010111010: data <= 8'h00; 
        10'b0010111011: data <= 8'h00; 
        10'b0010111100: data <= 8'h00; 
        10'b0010111101: data <= 8'hff; 
        10'b0010111110: data <= 8'hff; 
        10'b0010111111: data <= 8'hff; 
        10'b0011000000: data <= 8'h00; 
        10'b0011000001: data <= 8'h00; 
        10'b0011000010: data <= 8'h00; 
        10'b0011000011: data <= 8'h00; 
        10'b0011000100: data <= 8'h00; 
        10'b0011000101: data <= 8'h00; 
        10'b0011000110: data <= 8'h00; 
        10'b0011000111: data <= 8'h00; 
        10'b0011001000: data <= 8'h00; 
        10'b0011001001: data <= 8'h00; 
        10'b0011001010: data <= 8'h01; 
        10'b0011001011: data <= 8'h01; 
        10'b0011001100: data <= 8'h01; 
        10'b0011001101: data <= 8'h01; 
        10'b0011001110: data <= 8'h00; 
        10'b0011001111: data <= 8'h00; 
        10'b0011010000: data <= 8'h00; 
        10'b0011010001: data <= 8'h00; 
        10'b0011010010: data <= 8'h01; 
        10'b0011010011: data <= 8'h00; 
        10'b0011010100: data <= 8'h00; 
        10'b0011010101: data <= 8'hff; 
        10'b0011010110: data <= 8'h00; 
        10'b0011010111: data <= 8'h00; 
        10'b0011011000: data <= 8'h00; 
        10'b0011011001: data <= 8'h00; 
        10'b0011011010: data <= 8'h00; 
        10'b0011011011: data <= 8'hff; 
        10'b0011011100: data <= 8'h00; 
        10'b0011011101: data <= 8'h00; 
        10'b0011011110: data <= 8'h00; 
        10'b0011011111: data <= 8'h00; 
        10'b0011100000: data <= 8'h00; 
        10'b0011100001: data <= 8'h00; 
        10'b0011100010: data <= 8'h00; 
        10'b0011100011: data <= 8'h00; 
        10'b0011100100: data <= 8'h00; 
        10'b0011100101: data <= 8'h00; 
        10'b0011100110: data <= 8'h00; 
        10'b0011100111: data <= 8'h00; 
        10'b0011101000: data <= 8'h00; 
        10'b0011101001: data <= 8'h00; 
        10'b0011101010: data <= 8'h00; 
        10'b0011101011: data <= 8'h00; 
        10'b0011101100: data <= 8'h00; 
        10'b0011101101: data <= 8'h00; 
        10'b0011101110: data <= 8'h01; 
        10'b0011101111: data <= 8'h01; 
        10'b0011110000: data <= 8'h00; 
        10'b0011110001: data <= 8'h00; 
        10'b0011110010: data <= 8'h00; 
        10'b0011110011: data <= 8'h00; 
        10'b0011110100: data <= 8'h00; 
        10'b0011110101: data <= 8'h00; 
        10'b0011110110: data <= 8'h00; 
        10'b0011110111: data <= 8'hff; 
        10'b0011111000: data <= 8'hff; 
        10'b0011111001: data <= 8'h00; 
        10'b0011111010: data <= 8'h00; 
        10'b0011111011: data <= 8'h00; 
        10'b0011111100: data <= 8'h00; 
        10'b0011111101: data <= 8'h00; 
        10'b0011111110: data <= 8'h00; 
        10'b0011111111: data <= 8'h00; 
        10'b0100000000: data <= 8'h00; 
        10'b0100000001: data <= 8'h00; 
        10'b0100000010: data <= 8'h00; 
        10'b0100000011: data <= 8'h00; 
        10'b0100000100: data <= 8'h00; 
        10'b0100000101: data <= 8'h00; 
        10'b0100000110: data <= 8'h00; 
        10'b0100000111: data <= 8'h00; 
        10'b0100001000: data <= 8'h00; 
        10'b0100001001: data <= 8'h00; 
        10'b0100001010: data <= 8'h01; 
        10'b0100001011: data <= 8'h01; 
        10'b0100001100: data <= 8'h00; 
        10'b0100001101: data <= 8'h00; 
        10'b0100001110: data <= 8'h00; 
        10'b0100001111: data <= 8'h00; 
        10'b0100010000: data <= 8'h00; 
        10'b0100010001: data <= 8'h00; 
        10'b0100010010: data <= 8'h00; 
        10'b0100010011: data <= 8'hff; 
        10'b0100010100: data <= 8'hff; 
        10'b0100010101: data <= 8'h00; 
        10'b0100010110: data <= 8'h00; 
        10'b0100010111: data <= 8'h00; 
        10'b0100011000: data <= 8'h00; 
        10'b0100011001: data <= 8'h00; 
        10'b0100011010: data <= 8'h00; 
        10'b0100011011: data <= 8'h00; 
        10'b0100011100: data <= 8'h00; 
        10'b0100011101: data <= 8'h00; 
        10'b0100011110: data <= 8'h00; 
        10'b0100011111: data <= 8'hff; 
        10'b0100100000: data <= 8'hff; 
        10'b0100100001: data <= 8'hff; 
        10'b0100100010: data <= 8'hff; 
        10'b0100100011: data <= 8'hff; 
        10'b0100100100: data <= 8'hff; 
        10'b0100100101: data <= 8'hff; 
        10'b0100100110: data <= 8'hff; 
        10'b0100100111: data <= 8'h00; 
        10'b0100101000: data <= 8'h00; 
        10'b0100101001: data <= 8'h00; 
        10'b0100101010: data <= 8'h00; 
        10'b0100101011: data <= 8'h00; 
        10'b0100101100: data <= 8'h00; 
        10'b0100101101: data <= 8'h00; 
        10'b0100101110: data <= 8'h00; 
        10'b0100101111: data <= 8'hff; 
        10'b0100110000: data <= 8'h00; 
        10'b0100110001: data <= 8'h00; 
        10'b0100110010: data <= 8'h00; 
        10'b0100110011: data <= 8'h00; 
        10'b0100110100: data <= 8'h00; 
        10'b0100110101: data <= 8'h00; 
        10'b0100110110: data <= 8'h00; 
        10'b0100110111: data <= 8'h00; 
        10'b0100111000: data <= 8'h00; 
        10'b0100111001: data <= 8'hff; 
        10'b0100111010: data <= 8'hff; 
        10'b0100111011: data <= 8'hfe; 
        10'b0100111100: data <= 8'hfe; 
        10'b0100111101: data <= 8'hfe; 
        10'b0100111110: data <= 8'hfe; 
        10'b0100111111: data <= 8'hfe; 
        10'b0101000000: data <= 8'hfe; 
        10'b0101000001: data <= 8'hfd; 
        10'b0101000010: data <= 8'hfe; 
        10'b0101000011: data <= 8'hff; 
        10'b0101000100: data <= 8'h00; 
        10'b0101000101: data <= 8'h00; 
        10'b0101000110: data <= 8'h00; 
        10'b0101000111: data <= 8'h00; 
        10'b0101001000: data <= 8'h00; 
        10'b0101001001: data <= 8'h00; 
        10'b0101001010: data <= 8'h00; 
        10'b0101001011: data <= 8'h00; 
        10'b0101001100: data <= 8'h00; 
        10'b0101001101: data <= 8'h00; 
        10'b0101001110: data <= 8'h00; 
        10'b0101001111: data <= 8'h00; 
        10'b0101010000: data <= 8'h00; 
        10'b0101010001: data <= 8'h00; 
        10'b0101010010: data <= 8'h00; 
        10'b0101010011: data <= 8'h00; 
        10'b0101010100: data <= 8'h00; 
        10'b0101010101: data <= 8'hff; 
        10'b0101010110: data <= 8'hfe; 
        10'b0101010111: data <= 8'hfd; 
        10'b0101011000: data <= 8'hfd; 
        10'b0101011001: data <= 8'hfd; 
        10'b0101011010: data <= 8'hfe; 
        10'b0101011011: data <= 8'hfe; 
        10'b0101011100: data <= 8'hfe; 
        10'b0101011101: data <= 8'hfe; 
        10'b0101011110: data <= 8'hfe; 
        10'b0101011111: data <= 8'hff; 
        10'b0101100000: data <= 8'hff; 
        10'b0101100001: data <= 8'hff; 
        10'b0101100010: data <= 8'h00; 
        10'b0101100011: data <= 8'h00; 
        10'b0101100100: data <= 8'h00; 
        10'b0101100101: data <= 8'h00; 
        10'b0101100110: data <= 8'h00; 
        10'b0101100111: data <= 8'hff; 
        10'b0101101000: data <= 8'h00; 
        10'b0101101001: data <= 8'h00; 
        10'b0101101010: data <= 8'h00; 
        10'b0101101011: data <= 8'h00; 
        10'b0101101100: data <= 8'h00; 
        10'b0101101101: data <= 8'h00; 
        10'b0101101110: data <= 8'h00; 
        10'b0101101111: data <= 8'h00; 
        10'b0101110000: data <= 8'hff; 
        10'b0101110001: data <= 8'hfe; 
        10'b0101110010: data <= 8'hfe; 
        10'b0101110011: data <= 8'hfe; 
        10'b0101110100: data <= 8'hfe; 
        10'b0101110101: data <= 8'hff; 
        10'b0101110110: data <= 8'hff; 
        10'b0101110111: data <= 8'h00; 
        10'b0101111000: data <= 8'hff; 
        10'b0101111001: data <= 8'h00; 
        10'b0101111010: data <= 8'hff; 
        10'b0101111011: data <= 8'hff; 
        10'b0101111100: data <= 8'hff; 
        10'b0101111101: data <= 8'hff; 
        10'b0101111110: data <= 8'h00; 
        10'b0101111111: data <= 8'h00; 
        10'b0110000000: data <= 8'h00; 
        10'b0110000001: data <= 8'h00; 
        10'b0110000010: data <= 8'hff; 
        10'b0110000011: data <= 8'hff; 
        10'b0110000100: data <= 8'h00; 
        10'b0110000101: data <= 8'h00; 
        10'b0110000110: data <= 8'h00; 
        10'b0110000111: data <= 8'h00; 
        10'b0110001000: data <= 8'h00; 
        10'b0110001001: data <= 8'h00; 
        10'b0110001010: data <= 8'h00; 
        10'b0110001011: data <= 8'h00; 
        10'b0110001100: data <= 8'h00; 
        10'b0110001101: data <= 8'hff; 
        10'b0110001110: data <= 8'hff; 
        10'b0110001111: data <= 8'hff; 
        10'b0110010000: data <= 8'h00; 
        10'b0110010001: data <= 8'h00; 
        10'b0110010010: data <= 8'h00; 
        10'b0110010011: data <= 8'h00; 
        10'b0110010100: data <= 8'h00; 
        10'b0110010101: data <= 8'h01; 
        10'b0110010110: data <= 8'h00; 
        10'b0110010111: data <= 8'h00; 
        10'b0110011000: data <= 8'h00; 
        10'b0110011001: data <= 8'hff; 
        10'b0110011010: data <= 8'h00; 
        10'b0110011011: data <= 8'h00; 
        10'b0110011100: data <= 8'h00; 
        10'b0110011101: data <= 8'h00; 
        10'b0110011110: data <= 8'hff; 
        10'b0110011111: data <= 8'hff; 
        10'b0110100000: data <= 8'h00; 
        10'b0110100001: data <= 8'h00; 
        10'b0110100010: data <= 8'h00; 
        10'b0110100011: data <= 8'h00; 
        10'b0110100100: data <= 8'h00; 
        10'b0110100101: data <= 8'h00; 
        10'b0110100110: data <= 8'h00; 
        10'b0110100111: data <= 8'h00; 
        10'b0110101000: data <= 8'h00; 
        10'b0110101001: data <= 8'h00; 
        10'b0110101010: data <= 8'h00; 
        10'b0110101011: data <= 8'h00; 
        10'b0110101100: data <= 8'h01; 
        10'b0110101101: data <= 8'h00; 
        10'b0110101110: data <= 8'h01; 
        10'b0110101111: data <= 8'h00; 
        10'b0110110000: data <= 8'h00; 
        10'b0110110001: data <= 8'h01; 
        10'b0110110010: data <= 8'h00; 
        10'b0110110011: data <= 8'h00; 
        10'b0110110100: data <= 8'h00; 
        10'b0110110101: data <= 8'hff; 
        10'b0110110110: data <= 8'h00; 
        10'b0110110111: data <= 8'h00; 
        10'b0110111000: data <= 8'h00; 
        10'b0110111001: data <= 8'h00; 
        10'b0110111010: data <= 8'hff; 
        10'b0110111011: data <= 8'h00; 
        10'b0110111100: data <= 8'h00; 
        10'b0110111101: data <= 8'h00; 
        10'b0110111110: data <= 8'h00; 
        10'b0110111111: data <= 8'h00; 
        10'b0111000000: data <= 8'h00; 
        10'b0111000001: data <= 8'h00; 
        10'b0111000010: data <= 8'h00; 
        10'b0111000011: data <= 8'h00; 
        10'b0111000100: data <= 8'h01; 
        10'b0111000101: data <= 8'h01; 
        10'b0111000110: data <= 8'h01; 
        10'b0111000111: data <= 8'h01; 
        10'b0111001000: data <= 8'h00; 
        10'b0111001001: data <= 8'h00; 
        10'b0111001010: data <= 8'h00; 
        10'b0111001011: data <= 8'h00; 
        10'b0111001100: data <= 8'h01; 
        10'b0111001101: data <= 8'h01; 
        10'b0111001110: data <= 8'h00; 
        10'b0111001111: data <= 8'h00; 
        10'b0111010000: data <= 8'h00; 
        10'b0111010001: data <= 8'h00; 
        10'b0111010010: data <= 8'h00; 
        10'b0111010011: data <= 8'h00; 
        10'b0111010100: data <= 8'h00; 
        10'b0111010101: data <= 8'h00; 
        10'b0111010110: data <= 8'h00; 
        10'b0111010111: data <= 8'h00; 
        10'b0111011000: data <= 8'h01; 
        10'b0111011001: data <= 8'h01; 
        10'b0111011010: data <= 8'h00; 
        10'b0111011011: data <= 8'h00; 
        10'b0111011100: data <= 8'h00; 
        10'b0111011101: data <= 8'h00; 
        10'b0111011110: data <= 8'h00; 
        10'b0111011111: data <= 8'h00; 
        10'b0111100000: data <= 8'h01; 
        10'b0111100001: data <= 8'h01; 
        10'b0111100010: data <= 8'h01; 
        10'b0111100011: data <= 8'h01; 
        10'b0111100100: data <= 8'h01; 
        10'b0111100101: data <= 8'h01; 
        10'b0111100110: data <= 8'h01; 
        10'b0111100111: data <= 8'h01; 
        10'b0111101000: data <= 8'h01; 
        10'b0111101001: data <= 8'h00; 
        10'b0111101010: data <= 8'h00; 
        10'b0111101011: data <= 8'h00; 
        10'b0111101100: data <= 8'h00; 
        10'b0111101101: data <= 8'h00; 
        10'b0111101110: data <= 8'h00; 
        10'b0111101111: data <= 8'h00; 
        10'b0111110000: data <= 8'h00; 
        10'b0111110001: data <= 8'h00; 
        10'b0111110010: data <= 8'h00; 
        10'b0111110011: data <= 8'h00; 
        10'b0111110100: data <= 8'h01; 
        10'b0111110101: data <= 8'h01; 
        10'b0111110110: data <= 8'h00; 
        10'b0111110111: data <= 8'h00; 
        10'b0111111000: data <= 8'h00; 
        10'b0111111001: data <= 8'h00; 
        10'b0111111010: data <= 8'h00; 
        10'b0111111011: data <= 8'h00; 
        10'b0111111100: data <= 8'h01; 
        10'b0111111101: data <= 8'h02; 
        10'b0111111110: data <= 8'h02; 
        10'b0111111111: data <= 8'h01; 
        10'b1000000000: data <= 8'h01; 
        10'b1000000001: data <= 8'h01; 
        10'b1000000010: data <= 8'h01; 
        10'b1000000011: data <= 8'h01; 
        10'b1000000100: data <= 8'h02; 
        10'b1000000101: data <= 8'h01; 
        10'b1000000110: data <= 8'h01; 
        10'b1000000111: data <= 8'h01; 
        10'b1000001000: data <= 8'h00; 
        10'b1000001001: data <= 8'h01; 
        10'b1000001010: data <= 8'h00; 
        10'b1000001011: data <= 8'h00; 
        10'b1000001100: data <= 8'h01; 
        10'b1000001101: data <= 8'h01; 
        10'b1000001110: data <= 8'h01; 
        10'b1000001111: data <= 8'h01; 
        10'b1000010000: data <= 8'h02; 
        10'b1000010001: data <= 8'h01; 
        10'b1000010010: data <= 8'h00; 
        10'b1000010011: data <= 8'h00; 
        10'b1000010100: data <= 8'h00; 
        10'b1000010101: data <= 8'h00; 
        10'b1000010110: data <= 8'h00; 
        10'b1000010111: data <= 8'h00; 
        10'b1000011000: data <= 8'h01; 
        10'b1000011001: data <= 8'h01; 
        10'b1000011010: data <= 8'h01; 
        10'b1000011011: data <= 8'h01; 
        10'b1000011100: data <= 8'h01; 
        10'b1000011101: data <= 8'h01; 
        10'b1000011110: data <= 8'h01; 
        10'b1000011111: data <= 8'h01; 
        10'b1000100000: data <= 8'h01; 
        10'b1000100001: data <= 8'h01; 
        10'b1000100010: data <= 8'h01; 
        10'b1000100011: data <= 8'h00; 
        10'b1000100100: data <= 8'h00; 
        10'b1000100101: data <= 8'h01; 
        10'b1000100110: data <= 8'h00; 
        10'b1000100111: data <= 8'h00; 
        10'b1000101000: data <= 8'h01; 
        10'b1000101001: data <= 8'h01; 
        10'b1000101010: data <= 8'h01; 
        10'b1000101011: data <= 8'h01; 
        10'b1000101100: data <= 8'h01; 
        10'b1000101101: data <= 8'h00; 
        10'b1000101110: data <= 8'h00; 
        10'b1000101111: data <= 8'h00; 
        10'b1000110000: data <= 8'h00; 
        10'b1000110001: data <= 8'h00; 
        10'b1000110010: data <= 8'h00; 
        10'b1000110011: data <= 8'h00; 
        10'b1000110100: data <= 8'h00; 
        10'b1000110101: data <= 8'h01; 
        10'b1000110110: data <= 8'h01; 
        10'b1000110111: data <= 8'h01; 
        10'b1000111000: data <= 8'h01; 
        10'b1000111001: data <= 8'h01; 
        10'b1000111010: data <= 8'h01; 
        10'b1000111011: data <= 8'h01; 
        10'b1000111100: data <= 8'h01; 
        10'b1000111101: data <= 8'h00; 
        10'b1000111110: data <= 8'h00; 
        10'b1000111111: data <= 8'h00; 
        10'b1001000000: data <= 8'h00; 
        10'b1001000001: data <= 8'h00; 
        10'b1001000010: data <= 8'h01; 
        10'b1001000011: data <= 8'h01; 
        10'b1001000100: data <= 8'h01; 
        10'b1001000101: data <= 8'h01; 
        10'b1001000110: data <= 8'h01; 
        10'b1001000111: data <= 8'h01; 
        10'b1001001000: data <= 8'h01; 
        10'b1001001001: data <= 8'h00; 
        10'b1001001010: data <= 8'h00; 
        10'b1001001011: data <= 8'h00; 
        10'b1001001100: data <= 8'h00; 
        10'b1001001101: data <= 8'h00; 
        10'b1001001110: data <= 8'h00; 
        10'b1001001111: data <= 8'h00; 
        10'b1001010000: data <= 8'h00; 
        10'b1001010001: data <= 8'h00; 
        10'b1001010010: data <= 8'h01; 
        10'b1001010011: data <= 8'h01; 
        10'b1001010100: data <= 8'h01; 
        10'b1001010101: data <= 8'h01; 
        10'b1001010110: data <= 8'h01; 
        10'b1001010111: data <= 8'h01; 
        10'b1001011000: data <= 8'h00; 
        10'b1001011001: data <= 8'h00; 
        10'b1001011010: data <= 8'h00; 
        10'b1001011011: data <= 8'h00; 
        10'b1001011100: data <= 8'h00; 
        10'b1001011101: data <= 8'h00; 
        10'b1001011110: data <= 8'h01; 
        10'b1001011111: data <= 8'h01; 
        10'b1001100000: data <= 8'h00; 
        10'b1001100001: data <= 8'h01; 
        10'b1001100010: data <= 8'h01; 
        10'b1001100011: data <= 8'h01; 
        10'b1001100100: data <= 8'h01; 
        10'b1001100101: data <= 8'h00; 
        10'b1001100110: data <= 8'h00; 
        10'b1001100111: data <= 8'h00; 
        10'b1001101000: data <= 8'h00; 
        10'b1001101001: data <= 8'h00; 
        10'b1001101010: data <= 8'h00; 
        10'b1001101011: data <= 8'h00; 
        10'b1001101100: data <= 8'h00; 
        10'b1001101101: data <= 8'h00; 
        10'b1001101110: data <= 8'h00; 
        10'b1001101111: data <= 8'h00; 
        10'b1001110000: data <= 8'h00; 
        10'b1001110001: data <= 8'h00; 
        10'b1001110010: data <= 8'h00; 
        10'b1001110011: data <= 8'h01; 
        10'b1001110100: data <= 8'h00; 
        10'b1001110101: data <= 8'h00; 
        10'b1001110110: data <= 8'hff; 
        10'b1001110111: data <= 8'h00; 
        10'b1001111000: data <= 8'h00; 
        10'b1001111001: data <= 8'h00; 
        10'b1001111010: data <= 8'h01; 
        10'b1001111011: data <= 8'h01; 
        10'b1001111100: data <= 8'h01; 
        10'b1001111101: data <= 8'h01; 
        10'b1001111110: data <= 8'h01; 
        10'b1001111111: data <= 8'h01; 
        10'b1010000000: data <= 8'h00; 
        10'b1010000001: data <= 8'h00; 
        10'b1010000010: data <= 8'h00; 
        10'b1010000011: data <= 8'h00; 
        10'b1010000100: data <= 8'h00; 
        10'b1010000101: data <= 8'h00; 
        10'b1010000110: data <= 8'h00; 
        10'b1010000111: data <= 8'h00; 
        10'b1010001000: data <= 8'h00; 
        10'b1010001001: data <= 8'h00; 
        10'b1010001010: data <= 8'h00; 
        10'b1010001011: data <= 8'h00; 
        10'b1010001100: data <= 8'h00; 
        10'b1010001101: data <= 8'h00; 
        10'b1010001110: data <= 8'h00; 
        10'b1010001111: data <= 8'h00; 
        10'b1010010000: data <= 8'h00; 
        10'b1010010001: data <= 8'h00; 
        10'b1010010010: data <= 8'h00; 
        10'b1010010011: data <= 8'hff; 
        10'b1010010100: data <= 8'hff; 
        10'b1010010101: data <= 8'h00; 
        10'b1010010110: data <= 8'h00; 
        10'b1010010111: data <= 8'h01; 
        10'b1010011000: data <= 8'h01; 
        10'b1010011001: data <= 8'h01; 
        10'b1010011010: data <= 8'h01; 
        10'b1010011011: data <= 8'h00; 
        10'b1010011100: data <= 8'h00; 
        10'b1010011101: data <= 8'h00; 
        10'b1010011110: data <= 8'h00; 
        10'b1010011111: data <= 8'h00; 
        10'b1010100000: data <= 8'h00; 
        10'b1010100001: data <= 8'h00; 
        10'b1010100010: data <= 8'h00; 
        10'b1010100011: data <= 8'h00; 
        10'b1010100100: data <= 8'h00; 
        10'b1010100101: data <= 8'h00; 
        10'b1010100110: data <= 8'hff; 
        10'b1010100111: data <= 8'hff; 
        10'b1010101000: data <= 8'hff; 
        10'b1010101001: data <= 8'hff; 
        10'b1010101010: data <= 8'hff; 
        10'b1010101011: data <= 8'hff; 
        10'b1010101100: data <= 8'hff; 
        10'b1010101101: data <= 8'h00; 
        10'b1010101110: data <= 8'h00; 
        10'b1010101111: data <= 8'hff; 
        10'b1010110000: data <= 8'h00; 
        10'b1010110001: data <= 8'h00; 
        10'b1010110010: data <= 8'h00; 
        10'b1010110011: data <= 8'h00; 
        10'b1010110100: data <= 8'h00; 
        10'b1010110101: data <= 8'h00; 
        10'b1010110110: data <= 8'h00; 
        10'b1010110111: data <= 8'h00; 
        10'b1010111000: data <= 8'h00; 
        10'b1010111001: data <= 8'h00; 
        10'b1010111010: data <= 8'h00; 
        10'b1010111011: data <= 8'h00; 
        10'b1010111100: data <= 8'h00; 
        10'b1010111101: data <= 8'h00; 
        10'b1010111110: data <= 8'h00; 
        10'b1010111111: data <= 8'h00; 
        10'b1011000000: data <= 8'h00; 
        10'b1011000001: data <= 8'h00; 
        10'b1011000010: data <= 8'h00; 
        10'b1011000011: data <= 8'hff; 
        10'b1011000100: data <= 8'hff; 
        10'b1011000101: data <= 8'hff; 
        10'b1011000110: data <= 8'hff; 
        10'b1011000111: data <= 8'hff; 
        10'b1011001000: data <= 8'h00; 
        10'b1011001001: data <= 8'h00; 
        10'b1011001010: data <= 8'hff; 
        10'b1011001011: data <= 8'h00; 
        10'b1011001100: data <= 8'h00; 
        10'b1011001101: data <= 8'h00; 
        10'b1011001110: data <= 8'h00; 
        10'b1011001111: data <= 8'h00; 
        10'b1011010000: data <= 8'h00; 
        10'b1011010001: data <= 8'h00; 
        10'b1011010010: data <= 8'h00; 
        10'b1011010011: data <= 8'h00; 
        10'b1011010100: data <= 8'h00; 
        10'b1011010101: data <= 8'h00; 
        10'b1011010110: data <= 8'h00; 
        10'b1011010111: data <= 8'h00; 
        10'b1011011000: data <= 8'h00; 
        10'b1011011001: data <= 8'h00; 
        10'b1011011010: data <= 8'h00; 
        10'b1011011011: data <= 8'h00; 
        10'b1011011100: data <= 8'h00; 
        10'b1011011101: data <= 8'h00; 
        10'b1011011110: data <= 8'h00; 
        10'b1011011111: data <= 8'h00; 
        10'b1011100000: data <= 8'h00; 
        10'b1011100001: data <= 8'h00; 
        10'b1011100010: data <= 8'h00; 
        10'b1011100011: data <= 8'h00; 
        10'b1011100100: data <= 8'h00; 
        10'b1011100101: data <= 8'h00; 
        10'b1011100110: data <= 8'h00; 
        10'b1011100111: data <= 8'h00; 
        10'b1011101000: data <= 8'h00; 
        10'b1011101001: data <= 8'h00; 
        10'b1011101010: data <= 8'h00; 
        10'b1011101011: data <= 8'h00; 
        10'b1011101100: data <= 8'h00; 
        10'b1011101101: data <= 8'h00; 
        10'b1011101110: data <= 8'h00; 
        10'b1011101111: data <= 8'h00; 
        10'b1011110000: data <= 8'h00; 
        10'b1011110001: data <= 8'h00; 
        10'b1011110010: data <= 8'h00; 
        10'b1011110011: data <= 8'h00; 
        10'b1011110100: data <= 8'h00; 
        10'b1011110101: data <= 8'h00; 
        10'b1011110110: data <= 8'h00; 
        10'b1011110111: data <= 8'h00; 
        10'b1011111000: data <= 8'h00; 
        10'b1011111001: data <= 8'h00; 
        10'b1011111010: data <= 8'h00; 
        10'b1011111011: data <= 8'h00; 
        10'b1011111100: data <= 8'h00; 
        10'b1011111101: data <= 8'h00; 
        10'b1011111110: data <= 8'h00; 
        10'b1011111111: data <= 8'h00; 
        10'b1100000000: data <= 8'h00; 
        10'b1100000001: data <= 8'h00; 
        10'b1100000010: data <= 8'h00; 
        10'b1100000011: data <= 8'h00; 
        10'b1100000100: data <= 8'h00; 
        10'b1100000101: data <= 8'h00; 
        10'b1100000110: data <= 8'h00; 
        10'b1100000111: data <= 8'h00; 
        10'b1100001000: data <= 8'h00; 
        10'b1100001001: data <= 8'h00; 
        10'b1100001010: data <= 8'h00; 
        10'b1100001011: data <= 8'h00; 
        10'b1100001100: data <= 8'h00; 
        10'b1100001101: data <= 8'h00; 
        10'b1100001110: data <= 8'h00; 
        10'b1100001111: data <= 8'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 3) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 9'h000; 
        10'b0000000001: data <= 9'h000; 
        10'b0000000010: data <= 9'h000; 
        10'b0000000011: data <= 9'h000; 
        10'b0000000100: data <= 9'h000; 
        10'b0000000101: data <= 9'h000; 
        10'b0000000110: data <= 9'h000; 
        10'b0000000111: data <= 9'h000; 
        10'b0000001000: data <= 9'h000; 
        10'b0000001001: data <= 9'h000; 
        10'b0000001010: data <= 9'h000; 
        10'b0000001011: data <= 9'h000; 
        10'b0000001100: data <= 9'h000; 
        10'b0000001101: data <= 9'h000; 
        10'b0000001110: data <= 9'h000; 
        10'b0000001111: data <= 9'h000; 
        10'b0000010000: data <= 9'h000; 
        10'b0000010001: data <= 9'h000; 
        10'b0000010010: data <= 9'h000; 
        10'b0000010011: data <= 9'h000; 
        10'b0000010100: data <= 9'h000; 
        10'b0000010101: data <= 9'h000; 
        10'b0000010110: data <= 9'h000; 
        10'b0000010111: data <= 9'h000; 
        10'b0000011000: data <= 9'h000; 
        10'b0000011001: data <= 9'h000; 
        10'b0000011010: data <= 9'h000; 
        10'b0000011011: data <= 9'h000; 
        10'b0000011100: data <= 9'h000; 
        10'b0000011101: data <= 9'h000; 
        10'b0000011110: data <= 9'h000; 
        10'b0000011111: data <= 9'h000; 
        10'b0000100000: data <= 9'h000; 
        10'b0000100001: data <= 9'h000; 
        10'b0000100010: data <= 9'h000; 
        10'b0000100011: data <= 9'h000; 
        10'b0000100100: data <= 9'h000; 
        10'b0000100101: data <= 9'h000; 
        10'b0000100110: data <= 9'h000; 
        10'b0000100111: data <= 9'h000; 
        10'b0000101000: data <= 9'h000; 
        10'b0000101001: data <= 9'h000; 
        10'b0000101010: data <= 9'h000; 
        10'b0000101011: data <= 9'h000; 
        10'b0000101100: data <= 9'h000; 
        10'b0000101101: data <= 9'h000; 
        10'b0000101110: data <= 9'h000; 
        10'b0000101111: data <= 9'h000; 
        10'b0000110000: data <= 9'h000; 
        10'b0000110001: data <= 9'h000; 
        10'b0000110010: data <= 9'h000; 
        10'b0000110011: data <= 9'h000; 
        10'b0000110100: data <= 9'h000; 
        10'b0000110101: data <= 9'h000; 
        10'b0000110110: data <= 9'h000; 
        10'b0000110111: data <= 9'h000; 
        10'b0000111000: data <= 9'h000; 
        10'b0000111001: data <= 9'h000; 
        10'b0000111010: data <= 9'h000; 
        10'b0000111011: data <= 9'h000; 
        10'b0000111100: data <= 9'h000; 
        10'b0000111101: data <= 9'h000; 
        10'b0000111110: data <= 9'h000; 
        10'b0000111111: data <= 9'h000; 
        10'b0001000000: data <= 9'h000; 
        10'b0001000001: data <= 9'h000; 
        10'b0001000010: data <= 9'h000; 
        10'b0001000011: data <= 9'h000; 
        10'b0001000100: data <= 9'h001; 
        10'b0001000101: data <= 9'h000; 
        10'b0001000110: data <= 9'h000; 
        10'b0001000111: data <= 9'h000; 
        10'b0001001000: data <= 9'h001; 
        10'b0001001001: data <= 9'h000; 
        10'b0001001010: data <= 9'h000; 
        10'b0001001011: data <= 9'h000; 
        10'b0001001100: data <= 9'h000; 
        10'b0001001101: data <= 9'h000; 
        10'b0001001110: data <= 9'h1ff; 
        10'b0001001111: data <= 9'h000; 
        10'b0001010000: data <= 9'h000; 
        10'b0001010001: data <= 9'h000; 
        10'b0001010010: data <= 9'h000; 
        10'b0001010011: data <= 9'h000; 
        10'b0001010100: data <= 9'h000; 
        10'b0001010101: data <= 9'h000; 
        10'b0001010110: data <= 9'h000; 
        10'b0001010111: data <= 9'h000; 
        10'b0001011000: data <= 9'h000; 
        10'b0001011001: data <= 9'h000; 
        10'b0001011010: data <= 9'h000; 
        10'b0001011011: data <= 9'h000; 
        10'b0001011100: data <= 9'h000; 
        10'b0001011101: data <= 9'h001; 
        10'b0001011110: data <= 9'h001; 
        10'b0001011111: data <= 9'h001; 
        10'b0001100000: data <= 9'h001; 
        10'b0001100001: data <= 9'h002; 
        10'b0001100010: data <= 9'h001; 
        10'b0001100011: data <= 9'h000; 
        10'b0001100100: data <= 9'h001; 
        10'b0001100101: data <= 9'h000; 
        10'b0001100110: data <= 9'h000; 
        10'b0001100111: data <= 9'h000; 
        10'b0001101000: data <= 9'h000; 
        10'b0001101001: data <= 9'h1ff; 
        10'b0001101010: data <= 9'h1ff; 
        10'b0001101011: data <= 9'h000; 
        10'b0001101100: data <= 9'h000; 
        10'b0001101101: data <= 9'h000; 
        10'b0001101110: data <= 9'h000; 
        10'b0001101111: data <= 9'h000; 
        10'b0001110000: data <= 9'h000; 
        10'b0001110001: data <= 9'h000; 
        10'b0001110010: data <= 9'h000; 
        10'b0001110011: data <= 9'h000; 
        10'b0001110100: data <= 9'h000; 
        10'b0001110101: data <= 9'h000; 
        10'b0001110110: data <= 9'h000; 
        10'b0001110111: data <= 9'h000; 
        10'b0001111000: data <= 9'h001; 
        10'b0001111001: data <= 9'h002; 
        10'b0001111010: data <= 9'h002; 
        10'b0001111011: data <= 9'h002; 
        10'b0001111100: data <= 9'h002; 
        10'b0001111101: data <= 9'h001; 
        10'b0001111110: data <= 9'h001; 
        10'b0001111111: data <= 9'h001; 
        10'b0010000000: data <= 9'h001; 
        10'b0010000001: data <= 9'h001; 
        10'b0010000010: data <= 9'h000; 
        10'b0010000011: data <= 9'h000; 
        10'b0010000100: data <= 9'h000; 
        10'b0010000101: data <= 9'h1ff; 
        10'b0010000110: data <= 9'h1ff; 
        10'b0010000111: data <= 9'h1ff; 
        10'b0010001000: data <= 9'h000; 
        10'b0010001001: data <= 9'h000; 
        10'b0010001010: data <= 9'h000; 
        10'b0010001011: data <= 9'h000; 
        10'b0010001100: data <= 9'h000; 
        10'b0010001101: data <= 9'h000; 
        10'b0010001110: data <= 9'h000; 
        10'b0010001111: data <= 9'h000; 
        10'b0010010000: data <= 9'h000; 
        10'b0010010001: data <= 9'h000; 
        10'b0010010010: data <= 9'h000; 
        10'b0010010011: data <= 9'h001; 
        10'b0010010100: data <= 9'h001; 
        10'b0010010101: data <= 9'h002; 
        10'b0010010110: data <= 9'h002; 
        10'b0010010111: data <= 9'h002; 
        10'b0010011000: data <= 9'h002; 
        10'b0010011001: data <= 9'h002; 
        10'b0010011010: data <= 9'h002; 
        10'b0010011011: data <= 9'h002; 
        10'b0010011100: data <= 9'h002; 
        10'b0010011101: data <= 9'h002; 
        10'b0010011110: data <= 9'h001; 
        10'b0010011111: data <= 9'h1ff; 
        10'b0010100000: data <= 9'h1ff; 
        10'b0010100001: data <= 9'h1ff; 
        10'b0010100010: data <= 9'h1ff; 
        10'b0010100011: data <= 9'h1ff; 
        10'b0010100100: data <= 9'h1ff; 
        10'b0010100101: data <= 9'h000; 
        10'b0010100110: data <= 9'h000; 
        10'b0010100111: data <= 9'h000; 
        10'b0010101000: data <= 9'h000; 
        10'b0010101001: data <= 9'h000; 
        10'b0010101010: data <= 9'h000; 
        10'b0010101011: data <= 9'h000; 
        10'b0010101100: data <= 9'h000; 
        10'b0010101101: data <= 9'h000; 
        10'b0010101110: data <= 9'h001; 
        10'b0010101111: data <= 9'h002; 
        10'b0010110000: data <= 9'h001; 
        10'b0010110001: data <= 9'h001; 
        10'b0010110010: data <= 9'h002; 
        10'b0010110011: data <= 9'h001; 
        10'b0010110100: data <= 9'h001; 
        10'b0010110101: data <= 9'h002; 
        10'b0010110110: data <= 9'h001; 
        10'b0010110111: data <= 9'h001; 
        10'b0010111000: data <= 9'h001; 
        10'b0010111001: data <= 9'h000; 
        10'b0010111010: data <= 9'h000; 
        10'b0010111011: data <= 9'h1ff; 
        10'b0010111100: data <= 9'h000; 
        10'b0010111101: data <= 9'h1ff; 
        10'b0010111110: data <= 9'h1ff; 
        10'b0010111111: data <= 9'h1fe; 
        10'b0011000000: data <= 9'h1ff; 
        10'b0011000001: data <= 9'h1ff; 
        10'b0011000010: data <= 9'h000; 
        10'b0011000011: data <= 9'h000; 
        10'b0011000100: data <= 9'h000; 
        10'b0011000101: data <= 9'h000; 
        10'b0011000110: data <= 9'h000; 
        10'b0011000111: data <= 9'h000; 
        10'b0011001000: data <= 9'h000; 
        10'b0011001001: data <= 9'h000; 
        10'b0011001010: data <= 9'h001; 
        10'b0011001011: data <= 9'h002; 
        10'b0011001100: data <= 9'h001; 
        10'b0011001101: data <= 9'h001; 
        10'b0011001110: data <= 9'h000; 
        10'b0011001111: data <= 9'h001; 
        10'b0011010000: data <= 9'h000; 
        10'b0011010001: data <= 9'h001; 
        10'b0011010010: data <= 9'h001; 
        10'b0011010011: data <= 9'h000; 
        10'b0011010100: data <= 9'h000; 
        10'b0011010101: data <= 9'h1ff; 
        10'b0011010110: data <= 9'h000; 
        10'b0011010111: data <= 9'h000; 
        10'b0011011000: data <= 9'h000; 
        10'b0011011001: data <= 9'h000; 
        10'b0011011010: data <= 9'h000; 
        10'b0011011011: data <= 9'h1ff; 
        10'b0011011100: data <= 9'h1ff; 
        10'b0011011101: data <= 9'h000; 
        10'b0011011110: data <= 9'h000; 
        10'b0011011111: data <= 9'h000; 
        10'b0011100000: data <= 9'h000; 
        10'b0011100001: data <= 9'h000; 
        10'b0011100010: data <= 9'h000; 
        10'b0011100011: data <= 9'h000; 
        10'b0011100100: data <= 9'h000; 
        10'b0011100101: data <= 9'h001; 
        10'b0011100110: data <= 9'h001; 
        10'b0011100111: data <= 9'h001; 
        10'b0011101000: data <= 9'h001; 
        10'b0011101001: data <= 9'h001; 
        10'b0011101010: data <= 9'h001; 
        10'b0011101011: data <= 9'h001; 
        10'b0011101100: data <= 9'h001; 
        10'b0011101101: data <= 9'h001; 
        10'b0011101110: data <= 9'h002; 
        10'b0011101111: data <= 9'h001; 
        10'b0011110000: data <= 9'h000; 
        10'b0011110001: data <= 9'h000; 
        10'b0011110010: data <= 9'h000; 
        10'b0011110011: data <= 9'h000; 
        10'b0011110100: data <= 9'h000; 
        10'b0011110101: data <= 9'h000; 
        10'b0011110110: data <= 9'h1ff; 
        10'b0011110111: data <= 9'h1ff; 
        10'b0011111000: data <= 9'h1ff; 
        10'b0011111001: data <= 9'h000; 
        10'b0011111010: data <= 9'h000; 
        10'b0011111011: data <= 9'h000; 
        10'b0011111100: data <= 9'h000; 
        10'b0011111101: data <= 9'h000; 
        10'b0011111110: data <= 9'h000; 
        10'b0011111111: data <= 9'h000; 
        10'b0100000000: data <= 9'h000; 
        10'b0100000001: data <= 9'h001; 
        10'b0100000010: data <= 9'h000; 
        10'b0100000011: data <= 9'h000; 
        10'b0100000100: data <= 9'h000; 
        10'b0100000101: data <= 9'h000; 
        10'b0100000110: data <= 9'h000; 
        10'b0100000111: data <= 9'h000; 
        10'b0100001000: data <= 9'h000; 
        10'b0100001001: data <= 9'h000; 
        10'b0100001010: data <= 9'h001; 
        10'b0100001011: data <= 9'h001; 
        10'b0100001100: data <= 9'h000; 
        10'b0100001101: data <= 9'h000; 
        10'b0100001110: data <= 9'h000; 
        10'b0100001111: data <= 9'h000; 
        10'b0100010000: data <= 9'h000; 
        10'b0100010001: data <= 9'h000; 
        10'b0100010010: data <= 9'h000; 
        10'b0100010011: data <= 9'h1ff; 
        10'b0100010100: data <= 9'h1ff; 
        10'b0100010101: data <= 9'h000; 
        10'b0100010110: data <= 9'h000; 
        10'b0100010111: data <= 9'h000; 
        10'b0100011000: data <= 9'h000; 
        10'b0100011001: data <= 9'h000; 
        10'b0100011010: data <= 9'h000; 
        10'b0100011011: data <= 9'h000; 
        10'b0100011100: data <= 9'h000; 
        10'b0100011101: data <= 9'h000; 
        10'b0100011110: data <= 9'h000; 
        10'b0100011111: data <= 9'h1fe; 
        10'b0100100000: data <= 9'h1fe; 
        10'b0100100001: data <= 9'h1ff; 
        10'b0100100010: data <= 9'h1fe; 
        10'b0100100011: data <= 9'h1fe; 
        10'b0100100100: data <= 9'h1fd; 
        10'b0100100101: data <= 9'h1fd; 
        10'b0100100110: data <= 9'h1ff; 
        10'b0100100111: data <= 9'h000; 
        10'b0100101000: data <= 9'h000; 
        10'b0100101001: data <= 9'h000; 
        10'b0100101010: data <= 9'h000; 
        10'b0100101011: data <= 9'h000; 
        10'b0100101100: data <= 9'h000; 
        10'b0100101101: data <= 9'h000; 
        10'b0100101110: data <= 9'h1ff; 
        10'b0100101111: data <= 9'h1ff; 
        10'b0100110000: data <= 9'h1ff; 
        10'b0100110001: data <= 9'h000; 
        10'b0100110010: data <= 9'h000; 
        10'b0100110011: data <= 9'h000; 
        10'b0100110100: data <= 9'h000; 
        10'b0100110101: data <= 9'h000; 
        10'b0100110110: data <= 9'h000; 
        10'b0100110111: data <= 9'h000; 
        10'b0100111000: data <= 9'h1ff; 
        10'b0100111001: data <= 9'h1fe; 
        10'b0100111010: data <= 9'h1fd; 
        10'b0100111011: data <= 9'h1fc; 
        10'b0100111100: data <= 9'h1fc; 
        10'b0100111101: data <= 9'h1fc; 
        10'b0100111110: data <= 9'h1fc; 
        10'b0100111111: data <= 9'h1fc; 
        10'b0101000000: data <= 9'h1fc; 
        10'b0101000001: data <= 9'h1fb; 
        10'b0101000010: data <= 9'h1fc; 
        10'b0101000011: data <= 9'h1fe; 
        10'b0101000100: data <= 9'h1ff; 
        10'b0101000101: data <= 9'h1ff; 
        10'b0101000110: data <= 9'h1ff; 
        10'b0101000111: data <= 9'h000; 
        10'b0101001000: data <= 9'h000; 
        10'b0101001001: data <= 9'h000; 
        10'b0101001010: data <= 9'h1ff; 
        10'b0101001011: data <= 9'h1ff; 
        10'b0101001100: data <= 9'h000; 
        10'b0101001101: data <= 9'h000; 
        10'b0101001110: data <= 9'h000; 
        10'b0101001111: data <= 9'h000; 
        10'b0101010000: data <= 9'h000; 
        10'b0101010001: data <= 9'h000; 
        10'b0101010010: data <= 9'h000; 
        10'b0101010011: data <= 9'h000; 
        10'b0101010100: data <= 9'h1ff; 
        10'b0101010101: data <= 9'h1fe; 
        10'b0101010110: data <= 9'h1fb; 
        10'b0101010111: data <= 9'h1fa; 
        10'b0101011000: data <= 9'h1fb; 
        10'b0101011001: data <= 9'h1fb; 
        10'b0101011010: data <= 9'h1fb; 
        10'b0101011011: data <= 9'h1fc; 
        10'b0101011100: data <= 9'h1fc; 
        10'b0101011101: data <= 9'h1fb; 
        10'b0101011110: data <= 9'h1fc; 
        10'b0101011111: data <= 9'h1fe; 
        10'b0101100000: data <= 9'h1fe; 
        10'b0101100001: data <= 9'h1fe; 
        10'b0101100010: data <= 9'h1ff; 
        10'b0101100011: data <= 9'h000; 
        10'b0101100100: data <= 9'h000; 
        10'b0101100101: data <= 9'h000; 
        10'b0101100110: data <= 9'h1ff; 
        10'b0101100111: data <= 9'h1fe; 
        10'b0101101000: data <= 9'h000; 
        10'b0101101001: data <= 9'h000; 
        10'b0101101010: data <= 9'h000; 
        10'b0101101011: data <= 9'h000; 
        10'b0101101100: data <= 9'h000; 
        10'b0101101101: data <= 9'h000; 
        10'b0101101110: data <= 9'h000; 
        10'b0101101111: data <= 9'h000; 
        10'b0101110000: data <= 9'h1ff; 
        10'b0101110001: data <= 9'h1fd; 
        10'b0101110010: data <= 9'h1fb; 
        10'b0101110011: data <= 9'h1fc; 
        10'b0101110100: data <= 9'h1fc; 
        10'b0101110101: data <= 9'h1fd; 
        10'b0101110110: data <= 9'h1fe; 
        10'b0101110111: data <= 9'h1ff; 
        10'b0101111000: data <= 9'h1fe; 
        10'b0101111001: data <= 9'h1ff; 
        10'b0101111010: data <= 9'h1fe; 
        10'b0101111011: data <= 9'h1fe; 
        10'b0101111100: data <= 9'h1fe; 
        10'b0101111101: data <= 9'h1fe; 
        10'b0101111110: data <= 9'h1ff; 
        10'b0101111111: data <= 9'h000; 
        10'b0110000000: data <= 9'h000; 
        10'b0110000001: data <= 9'h1ff; 
        10'b0110000010: data <= 9'h1ff; 
        10'b0110000011: data <= 9'h1ff; 
        10'b0110000100: data <= 9'h1ff; 
        10'b0110000101: data <= 9'h000; 
        10'b0110000110: data <= 9'h000; 
        10'b0110000111: data <= 9'h000; 
        10'b0110001000: data <= 9'h000; 
        10'b0110001001: data <= 9'h000; 
        10'b0110001010: data <= 9'h000; 
        10'b0110001011: data <= 9'h000; 
        10'b0110001100: data <= 9'h000; 
        10'b0110001101: data <= 9'h1fe; 
        10'b0110001110: data <= 9'h1fd; 
        10'b0110001111: data <= 9'h1fe; 
        10'b0110010000: data <= 9'h1ff; 
        10'b0110010001: data <= 9'h000; 
        10'b0110010010: data <= 9'h001; 
        10'b0110010011: data <= 9'h001; 
        10'b0110010100: data <= 9'h001; 
        10'b0110010101: data <= 9'h001; 
        10'b0110010110: data <= 9'h000; 
        10'b0110010111: data <= 9'h1ff; 
        10'b0110011000: data <= 9'h1ff; 
        10'b0110011001: data <= 9'h1ff; 
        10'b0110011010: data <= 9'h000; 
        10'b0110011011: data <= 9'h1ff; 
        10'b0110011100: data <= 9'h000; 
        10'b0110011101: data <= 9'h1ff; 
        10'b0110011110: data <= 9'h1ff; 
        10'b0110011111: data <= 9'h1ff; 
        10'b0110100000: data <= 9'h000; 
        10'b0110100001: data <= 9'h001; 
        10'b0110100010: data <= 9'h001; 
        10'b0110100011: data <= 9'h000; 
        10'b0110100100: data <= 9'h000; 
        10'b0110100101: data <= 9'h000; 
        10'b0110100110: data <= 9'h000; 
        10'b0110100111: data <= 9'h000; 
        10'b0110101000: data <= 9'h000; 
        10'b0110101001: data <= 9'h000; 
        10'b0110101010: data <= 9'h001; 
        10'b0110101011: data <= 9'h001; 
        10'b0110101100: data <= 9'h001; 
        10'b0110101101: data <= 9'h001; 
        10'b0110101110: data <= 9'h001; 
        10'b0110101111: data <= 9'h001; 
        10'b0110110000: data <= 9'h001; 
        10'b0110110001: data <= 9'h001; 
        10'b0110110010: data <= 9'h000; 
        10'b0110110011: data <= 9'h000; 
        10'b0110110100: data <= 9'h000; 
        10'b0110110101: data <= 9'h1ff; 
        10'b0110110110: data <= 9'h1ff; 
        10'b0110110111: data <= 9'h1ff; 
        10'b0110111000: data <= 9'h000; 
        10'b0110111001: data <= 9'h1ff; 
        10'b0110111010: data <= 9'h1ff; 
        10'b0110111011: data <= 9'h1ff; 
        10'b0110111100: data <= 9'h000; 
        10'b0110111101: data <= 9'h001; 
        10'b0110111110: data <= 9'h000; 
        10'b0110111111: data <= 9'h000; 
        10'b0111000000: data <= 9'h000; 
        10'b0111000001: data <= 9'h000; 
        10'b0111000010: data <= 9'h000; 
        10'b0111000011: data <= 9'h001; 
        10'b0111000100: data <= 9'h001; 
        10'b0111000101: data <= 9'h002; 
        10'b0111000110: data <= 9'h002; 
        10'b0111000111: data <= 9'h001; 
        10'b0111001000: data <= 9'h000; 
        10'b0111001001: data <= 9'h001; 
        10'b0111001010: data <= 9'h001; 
        10'b0111001011: data <= 9'h001; 
        10'b0111001100: data <= 9'h002; 
        10'b0111001101: data <= 9'h001; 
        10'b0111001110: data <= 9'h000; 
        10'b0111001111: data <= 9'h000; 
        10'b0111010000: data <= 9'h000; 
        10'b0111010001: data <= 9'h1ff; 
        10'b0111010010: data <= 9'h1ff; 
        10'b0111010011: data <= 9'h1ff; 
        10'b0111010100: data <= 9'h000; 
        10'b0111010101: data <= 9'h000; 
        10'b0111010110: data <= 9'h000; 
        10'b0111010111: data <= 9'h000; 
        10'b0111011000: data <= 9'h001; 
        10'b0111011001: data <= 9'h002; 
        10'b0111011010: data <= 9'h000; 
        10'b0111011011: data <= 9'h000; 
        10'b0111011100: data <= 9'h000; 
        10'b0111011101: data <= 9'h000; 
        10'b0111011110: data <= 9'h000; 
        10'b0111011111: data <= 9'h001; 
        10'b0111100000: data <= 9'h002; 
        10'b0111100001: data <= 9'h003; 
        10'b0111100010: data <= 9'h002; 
        10'b0111100011: data <= 9'h002; 
        10'b0111100100: data <= 9'h001; 
        10'b0111100101: data <= 9'h001; 
        10'b0111100110: data <= 9'h002; 
        10'b0111100111: data <= 9'h002; 
        10'b0111101000: data <= 9'h002; 
        10'b0111101001: data <= 9'h001; 
        10'b0111101010: data <= 9'h000; 
        10'b0111101011: data <= 9'h001; 
        10'b0111101100: data <= 9'h001; 
        10'b0111101101: data <= 9'h000; 
        10'b0111101110: data <= 9'h000; 
        10'b0111101111: data <= 9'h000; 
        10'b0111110000: data <= 9'h001; 
        10'b0111110001: data <= 9'h001; 
        10'b0111110010: data <= 9'h001; 
        10'b0111110011: data <= 9'h001; 
        10'b0111110100: data <= 9'h002; 
        10'b0111110101: data <= 9'h002; 
        10'b0111110110: data <= 9'h000; 
        10'b0111110111: data <= 9'h000; 
        10'b0111111000: data <= 9'h000; 
        10'b0111111001: data <= 9'h000; 
        10'b0111111010: data <= 9'h1ff; 
        10'b0111111011: data <= 9'h000; 
        10'b0111111100: data <= 9'h002; 
        10'b0111111101: data <= 9'h003; 
        10'b0111111110: data <= 9'h003; 
        10'b0111111111: data <= 9'h002; 
        10'b1000000000: data <= 9'h001; 
        10'b1000000001: data <= 9'h002; 
        10'b1000000010: data <= 9'h003; 
        10'b1000000011: data <= 9'h002; 
        10'b1000000100: data <= 9'h004; 
        10'b1000000101: data <= 9'h003; 
        10'b1000000110: data <= 9'h002; 
        10'b1000000111: data <= 9'h001; 
        10'b1000001000: data <= 9'h001; 
        10'b1000001001: data <= 9'h001; 
        10'b1000001010: data <= 9'h001; 
        10'b1000001011: data <= 9'h001; 
        10'b1000001100: data <= 9'h002; 
        10'b1000001101: data <= 9'h002; 
        10'b1000001110: data <= 9'h002; 
        10'b1000001111: data <= 9'h003; 
        10'b1000010000: data <= 9'h003; 
        10'b1000010001: data <= 9'h002; 
        10'b1000010010: data <= 9'h000; 
        10'b1000010011: data <= 9'h000; 
        10'b1000010100: data <= 9'h000; 
        10'b1000010101: data <= 9'h000; 
        10'b1000010110: data <= 9'h000; 
        10'b1000010111: data <= 9'h000; 
        10'b1000011000: data <= 9'h001; 
        10'b1000011001: data <= 9'h002; 
        10'b1000011010: data <= 9'h003; 
        10'b1000011011: data <= 9'h002; 
        10'b1000011100: data <= 9'h002; 
        10'b1000011101: data <= 9'h002; 
        10'b1000011110: data <= 9'h002; 
        10'b1000011111: data <= 9'h002; 
        10'b1000100000: data <= 9'h002; 
        10'b1000100001: data <= 9'h002; 
        10'b1000100010: data <= 9'h001; 
        10'b1000100011: data <= 9'h001; 
        10'b1000100100: data <= 9'h001; 
        10'b1000100101: data <= 9'h002; 
        10'b1000100110: data <= 9'h001; 
        10'b1000100111: data <= 9'h001; 
        10'b1000101000: data <= 9'h001; 
        10'b1000101001: data <= 9'h002; 
        10'b1000101010: data <= 9'h002; 
        10'b1000101011: data <= 9'h002; 
        10'b1000101100: data <= 9'h002; 
        10'b1000101101: data <= 9'h001; 
        10'b1000101110: data <= 9'h000; 
        10'b1000101111: data <= 9'h000; 
        10'b1000110000: data <= 9'h000; 
        10'b1000110001: data <= 9'h000; 
        10'b1000110010: data <= 9'h000; 
        10'b1000110011: data <= 9'h1ff; 
        10'b1000110100: data <= 9'h001; 
        10'b1000110101: data <= 9'h001; 
        10'b1000110110: data <= 9'h002; 
        10'b1000110111: data <= 9'h003; 
        10'b1000111000: data <= 9'h002; 
        10'b1000111001: data <= 9'h002; 
        10'b1000111010: data <= 9'h002; 
        10'b1000111011: data <= 9'h003; 
        10'b1000111100: data <= 9'h001; 
        10'b1000111101: data <= 9'h000; 
        10'b1000111110: data <= 9'h000; 
        10'b1000111111: data <= 9'h000; 
        10'b1001000000: data <= 9'h001; 
        10'b1001000001: data <= 9'h000; 
        10'b1001000010: data <= 9'h001; 
        10'b1001000011: data <= 9'h002; 
        10'b1001000100: data <= 9'h001; 
        10'b1001000101: data <= 9'h002; 
        10'b1001000110: data <= 9'h002; 
        10'b1001000111: data <= 9'h002; 
        10'b1001001000: data <= 9'h001; 
        10'b1001001001: data <= 9'h001; 
        10'b1001001010: data <= 9'h000; 
        10'b1001001011: data <= 9'h000; 
        10'b1001001100: data <= 9'h000; 
        10'b1001001101: data <= 9'h000; 
        10'b1001001110: data <= 9'h000; 
        10'b1001001111: data <= 9'h000; 
        10'b1001010000: data <= 9'h000; 
        10'b1001010001: data <= 9'h001; 
        10'b1001010010: data <= 9'h001; 
        10'b1001010011: data <= 9'h001; 
        10'b1001010100: data <= 9'h001; 
        10'b1001010101: data <= 9'h002; 
        10'b1001010110: data <= 9'h001; 
        10'b1001010111: data <= 9'h001; 
        10'b1001011000: data <= 9'h001; 
        10'b1001011001: data <= 9'h000; 
        10'b1001011010: data <= 9'h000; 
        10'b1001011011: data <= 9'h000; 
        10'b1001011100: data <= 9'h001; 
        10'b1001011101: data <= 9'h001; 
        10'b1001011110: data <= 9'h002; 
        10'b1001011111: data <= 9'h002; 
        10'b1001100000: data <= 9'h001; 
        10'b1001100001: data <= 9'h002; 
        10'b1001100010: data <= 9'h002; 
        10'b1001100011: data <= 9'h002; 
        10'b1001100100: data <= 9'h001; 
        10'b1001100101: data <= 9'h000; 
        10'b1001100110: data <= 9'h000; 
        10'b1001100111: data <= 9'h000; 
        10'b1001101000: data <= 9'h000; 
        10'b1001101001: data <= 9'h000; 
        10'b1001101010: data <= 9'h000; 
        10'b1001101011: data <= 9'h000; 
        10'b1001101100: data <= 9'h000; 
        10'b1001101101: data <= 9'h000; 
        10'b1001101110: data <= 9'h001; 
        10'b1001101111: data <= 9'h001; 
        10'b1001110000: data <= 9'h001; 
        10'b1001110001: data <= 9'h001; 
        10'b1001110010: data <= 9'h001; 
        10'b1001110011: data <= 9'h001; 
        10'b1001110100: data <= 9'h000; 
        10'b1001110101: data <= 9'h1ff; 
        10'b1001110110: data <= 9'h1ff; 
        10'b1001110111: data <= 9'h1ff; 
        10'b1001111000: data <= 9'h1ff; 
        10'b1001111001: data <= 9'h000; 
        10'b1001111010: data <= 9'h002; 
        10'b1001111011: data <= 9'h002; 
        10'b1001111100: data <= 9'h002; 
        10'b1001111101: data <= 9'h002; 
        10'b1001111110: data <= 9'h001; 
        10'b1001111111: data <= 9'h002; 
        10'b1010000000: data <= 9'h001; 
        10'b1010000001: data <= 9'h000; 
        10'b1010000010: data <= 9'h000; 
        10'b1010000011: data <= 9'h000; 
        10'b1010000100: data <= 9'h000; 
        10'b1010000101: data <= 9'h000; 
        10'b1010000110: data <= 9'h000; 
        10'b1010000111: data <= 9'h000; 
        10'b1010001000: data <= 9'h000; 
        10'b1010001001: data <= 9'h000; 
        10'b1010001010: data <= 9'h1ff; 
        10'b1010001011: data <= 9'h000; 
        10'b1010001100: data <= 9'h1ff; 
        10'b1010001101: data <= 9'h000; 
        10'b1010001110: data <= 9'h000; 
        10'b1010001111: data <= 9'h000; 
        10'b1010010000: data <= 9'h000; 
        10'b1010010001: data <= 9'h1ff; 
        10'b1010010010: data <= 9'h1ff; 
        10'b1010010011: data <= 9'h1ff; 
        10'b1010010100: data <= 9'h1ff; 
        10'b1010010101: data <= 9'h1ff; 
        10'b1010010110: data <= 9'h000; 
        10'b1010010111: data <= 9'h002; 
        10'b1010011000: data <= 9'h001; 
        10'b1010011001: data <= 9'h002; 
        10'b1010011010: data <= 9'h001; 
        10'b1010011011: data <= 9'h000; 
        10'b1010011100: data <= 9'h000; 
        10'b1010011101: data <= 9'h000; 
        10'b1010011110: data <= 9'h000; 
        10'b1010011111: data <= 9'h000; 
        10'b1010100000: data <= 9'h000; 
        10'b1010100001: data <= 9'h000; 
        10'b1010100010: data <= 9'h000; 
        10'b1010100011: data <= 9'h000; 
        10'b1010100100: data <= 9'h000; 
        10'b1010100101: data <= 9'h1ff; 
        10'b1010100110: data <= 9'h1fe; 
        10'b1010100111: data <= 9'h1ff; 
        10'b1010101000: data <= 9'h1ff; 
        10'b1010101001: data <= 9'h1ff; 
        10'b1010101010: data <= 9'h1ff; 
        10'b1010101011: data <= 9'h1ff; 
        10'b1010101100: data <= 9'h1ff; 
        10'b1010101101: data <= 9'h1ff; 
        10'b1010101110: data <= 9'h1ff; 
        10'b1010101111: data <= 9'h1ff; 
        10'b1010110000: data <= 9'h1ff; 
        10'b1010110001: data <= 9'h1ff; 
        10'b1010110010: data <= 9'h1ff; 
        10'b1010110011: data <= 9'h1ff; 
        10'b1010110100: data <= 9'h000; 
        10'b1010110101: data <= 9'h000; 
        10'b1010110110: data <= 9'h000; 
        10'b1010110111: data <= 9'h000; 
        10'b1010111000: data <= 9'h000; 
        10'b1010111001: data <= 9'h000; 
        10'b1010111010: data <= 9'h000; 
        10'b1010111011: data <= 9'h000; 
        10'b1010111100: data <= 9'h000; 
        10'b1010111101: data <= 9'h000; 
        10'b1010111110: data <= 9'h000; 
        10'b1010111111: data <= 9'h000; 
        10'b1011000000: data <= 9'h000; 
        10'b1011000001: data <= 9'h1ff; 
        10'b1011000010: data <= 9'h1ff; 
        10'b1011000011: data <= 9'h1ff; 
        10'b1011000100: data <= 9'h1ff; 
        10'b1011000101: data <= 9'h1ff; 
        10'b1011000110: data <= 9'h1ff; 
        10'b1011000111: data <= 9'h1ff; 
        10'b1011001000: data <= 9'h1ff; 
        10'b1011001001: data <= 9'h1ff; 
        10'b1011001010: data <= 9'h1ff; 
        10'b1011001011: data <= 9'h1ff; 
        10'b1011001100: data <= 9'h1ff; 
        10'b1011001101: data <= 9'h1ff; 
        10'b1011001110: data <= 9'h000; 
        10'b1011001111: data <= 9'h1ff; 
        10'b1011010000: data <= 9'h000; 
        10'b1011010001: data <= 9'h000; 
        10'b1011010010: data <= 9'h000; 
        10'b1011010011: data <= 9'h000; 
        10'b1011010100: data <= 9'h000; 
        10'b1011010101: data <= 9'h000; 
        10'b1011010110: data <= 9'h000; 
        10'b1011010111: data <= 9'h000; 
        10'b1011011000: data <= 9'h000; 
        10'b1011011001: data <= 9'h000; 
        10'b1011011010: data <= 9'h000; 
        10'b1011011011: data <= 9'h000; 
        10'b1011011100: data <= 9'h000; 
        10'b1011011101: data <= 9'h000; 
        10'b1011011110: data <= 9'h000; 
        10'b1011011111: data <= 9'h000; 
        10'b1011100000: data <= 9'h000; 
        10'b1011100001: data <= 9'h000; 
        10'b1011100010: data <= 9'h000; 
        10'b1011100011: data <= 9'h000; 
        10'b1011100100: data <= 9'h000; 
        10'b1011100101: data <= 9'h000; 
        10'b1011100110: data <= 9'h000; 
        10'b1011100111: data <= 9'h000; 
        10'b1011101000: data <= 9'h000; 
        10'b1011101001: data <= 9'h000; 
        10'b1011101010: data <= 9'h000; 
        10'b1011101011: data <= 9'h000; 
        10'b1011101100: data <= 9'h000; 
        10'b1011101101: data <= 9'h000; 
        10'b1011101110: data <= 9'h000; 
        10'b1011101111: data <= 9'h000; 
        10'b1011110000: data <= 9'h000; 
        10'b1011110001: data <= 9'h000; 
        10'b1011110010: data <= 9'h000; 
        10'b1011110011: data <= 9'h000; 
        10'b1011110100: data <= 9'h000; 
        10'b1011110101: data <= 9'h000; 
        10'b1011110110: data <= 9'h000; 
        10'b1011110111: data <= 9'h000; 
        10'b1011111000: data <= 9'h000; 
        10'b1011111001: data <= 9'h000; 
        10'b1011111010: data <= 9'h000; 
        10'b1011111011: data <= 9'h000; 
        10'b1011111100: data <= 9'h000; 
        10'b1011111101: data <= 9'h000; 
        10'b1011111110: data <= 9'h000; 
        10'b1011111111: data <= 9'h000; 
        10'b1100000000: data <= 9'h000; 
        10'b1100000001: data <= 9'h000; 
        10'b1100000010: data <= 9'h000; 
        10'b1100000011: data <= 9'h000; 
        10'b1100000100: data <= 9'h000; 
        10'b1100000101: data <= 9'h000; 
        10'b1100000110: data <= 9'h000; 
        10'b1100000111: data <= 9'h000; 
        10'b1100001000: data <= 9'h000; 
        10'b1100001001: data <= 9'h000; 
        10'b1100001010: data <= 9'h000; 
        10'b1100001011: data <= 9'h000; 
        10'b1100001100: data <= 9'h000; 
        10'b1100001101: data <= 9'h000; 
        10'b1100001110: data <= 9'h000; 
        10'b1100001111: data <= 9'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 4) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 10'h3ff; 
        10'b0000000001: data <= 10'h000; 
        10'b0000000010: data <= 10'h000; 
        10'b0000000011: data <= 10'h3ff; 
        10'b0000000100: data <= 10'h000; 
        10'b0000000101: data <= 10'h3ff; 
        10'b0000000110: data <= 10'h000; 
        10'b0000000111: data <= 10'h000; 
        10'b0000001000: data <= 10'h3ff; 
        10'b0000001001: data <= 10'h000; 
        10'b0000001010: data <= 10'h3ff; 
        10'b0000001011: data <= 10'h3ff; 
        10'b0000001100: data <= 10'h000; 
        10'b0000001101: data <= 10'h000; 
        10'b0000001110: data <= 10'h3ff; 
        10'b0000001111: data <= 10'h000; 
        10'b0000010000: data <= 10'h3ff; 
        10'b0000010001: data <= 10'h3ff; 
        10'b0000010010: data <= 10'h000; 
        10'b0000010011: data <= 10'h000; 
        10'b0000010100: data <= 10'h3ff; 
        10'b0000010101: data <= 10'h000; 
        10'b0000010110: data <= 10'h3ff; 
        10'b0000010111: data <= 10'h3ff; 
        10'b0000011000: data <= 10'h3ff; 
        10'b0000011001: data <= 10'h000; 
        10'b0000011010: data <= 10'h000; 
        10'b0000011011: data <= 10'h000; 
        10'b0000011100: data <= 10'h000; 
        10'b0000011101: data <= 10'h000; 
        10'b0000011110: data <= 10'h000; 
        10'b0000011111: data <= 10'h000; 
        10'b0000100000: data <= 10'h3ff; 
        10'b0000100001: data <= 10'h3ff; 
        10'b0000100010: data <= 10'h3ff; 
        10'b0000100011: data <= 10'h3ff; 
        10'b0000100100: data <= 10'h3ff; 
        10'b0000100101: data <= 10'h000; 
        10'b0000100110: data <= 10'h000; 
        10'b0000100111: data <= 10'h3ff; 
        10'b0000101000: data <= 10'h000; 
        10'b0000101001: data <= 10'h3ff; 
        10'b0000101010: data <= 10'h000; 
        10'b0000101011: data <= 10'h3ff; 
        10'b0000101100: data <= 10'h000; 
        10'b0000101101: data <= 10'h3ff; 
        10'b0000101110: data <= 10'h000; 
        10'b0000101111: data <= 10'h3ff; 
        10'b0000110000: data <= 10'h000; 
        10'b0000110001: data <= 10'h3ff; 
        10'b0000110010: data <= 10'h3ff; 
        10'b0000110011: data <= 10'h3ff; 
        10'b0000110100: data <= 10'h000; 
        10'b0000110101: data <= 10'h000; 
        10'b0000110110: data <= 10'h000; 
        10'b0000110111: data <= 10'h3ff; 
        10'b0000111000: data <= 10'h000; 
        10'b0000111001: data <= 10'h3ff; 
        10'b0000111010: data <= 10'h3ff; 
        10'b0000111011: data <= 10'h000; 
        10'b0000111100: data <= 10'h3ff; 
        10'b0000111101: data <= 10'h3ff; 
        10'b0000111110: data <= 10'h000; 
        10'b0000111111: data <= 10'h000; 
        10'b0001000000: data <= 10'h000; 
        10'b0001000001: data <= 10'h000; 
        10'b0001000010: data <= 10'h000; 
        10'b0001000011: data <= 10'h000; 
        10'b0001000100: data <= 10'h001; 
        10'b0001000101: data <= 10'h001; 
        10'b0001000110: data <= 10'h001; 
        10'b0001000111: data <= 10'h000; 
        10'b0001001000: data <= 10'h001; 
        10'b0001001001: data <= 10'h000; 
        10'b0001001010: data <= 10'h000; 
        10'b0001001011: data <= 10'h3ff; 
        10'b0001001100: data <= 10'h000; 
        10'b0001001101: data <= 10'h000; 
        10'b0001001110: data <= 10'h3ff; 
        10'b0001001111: data <= 10'h000; 
        10'b0001010000: data <= 10'h000; 
        10'b0001010001: data <= 10'h000; 
        10'b0001010010: data <= 10'h000; 
        10'b0001010011: data <= 10'h000; 
        10'b0001010100: data <= 10'h3ff; 
        10'b0001010101: data <= 10'h3ff; 
        10'b0001010110: data <= 10'h000; 
        10'b0001010111: data <= 10'h3ff; 
        10'b0001011000: data <= 10'h000; 
        10'b0001011001: data <= 10'h3ff; 
        10'b0001011010: data <= 10'h000; 
        10'b0001011011: data <= 10'h000; 
        10'b0001011100: data <= 10'h000; 
        10'b0001011101: data <= 10'h002; 
        10'b0001011110: data <= 10'h003; 
        10'b0001011111: data <= 10'h003; 
        10'b0001100000: data <= 10'h003; 
        10'b0001100001: data <= 10'h004; 
        10'b0001100010: data <= 10'h002; 
        10'b0001100011: data <= 10'h001; 
        10'b0001100100: data <= 10'h002; 
        10'b0001100101: data <= 10'h001; 
        10'b0001100110: data <= 10'h3ff; 
        10'b0001100111: data <= 10'h000; 
        10'b0001101000: data <= 10'h3ff; 
        10'b0001101001: data <= 10'h3ff; 
        10'b0001101010: data <= 10'h3ff; 
        10'b0001101011: data <= 10'h3ff; 
        10'b0001101100: data <= 10'h000; 
        10'b0001101101: data <= 10'h000; 
        10'b0001101110: data <= 10'h3ff; 
        10'b0001101111: data <= 10'h000; 
        10'b0001110000: data <= 10'h3ff; 
        10'b0001110001: data <= 10'h000; 
        10'b0001110010: data <= 10'h000; 
        10'b0001110011: data <= 10'h3ff; 
        10'b0001110100: data <= 10'h3ff; 
        10'b0001110101: data <= 10'h000; 
        10'b0001110110: data <= 10'h000; 
        10'b0001110111: data <= 10'h000; 
        10'b0001111000: data <= 10'h001; 
        10'b0001111001: data <= 10'h004; 
        10'b0001111010: data <= 10'h004; 
        10'b0001111011: data <= 10'h004; 
        10'b0001111100: data <= 10'h004; 
        10'b0001111101: data <= 10'h003; 
        10'b0001111110: data <= 10'h003; 
        10'b0001111111: data <= 10'h001; 
        10'b0010000000: data <= 10'h002; 
        10'b0010000001: data <= 10'h001; 
        10'b0010000010: data <= 10'h000; 
        10'b0010000011: data <= 10'h3ff; 
        10'b0010000100: data <= 10'h3ff; 
        10'b0010000101: data <= 10'h3fe; 
        10'b0010000110: data <= 10'h3fe; 
        10'b0010000111: data <= 10'h3fe; 
        10'b0010001000: data <= 10'h000; 
        10'b0010001001: data <= 10'h000; 
        10'b0010001010: data <= 10'h3ff; 
        10'b0010001011: data <= 10'h000; 
        10'b0010001100: data <= 10'h000; 
        10'b0010001101: data <= 10'h000; 
        10'b0010001110: data <= 10'h3ff; 
        10'b0010001111: data <= 10'h3ff; 
        10'b0010010000: data <= 10'h3ff; 
        10'b0010010001: data <= 10'h3ff; 
        10'b0010010010: data <= 10'h000; 
        10'b0010010011: data <= 10'h002; 
        10'b0010010100: data <= 10'h002; 
        10'b0010010101: data <= 10'h004; 
        10'b0010010110: data <= 10'h005; 
        10'b0010010111: data <= 10'h005; 
        10'b0010011000: data <= 10'h004; 
        10'b0010011001: data <= 10'h005; 
        10'b0010011010: data <= 10'h004; 
        10'b0010011011: data <= 10'h004; 
        10'b0010011100: data <= 10'h005; 
        10'b0010011101: data <= 10'h004; 
        10'b0010011110: data <= 10'h003; 
        10'b0010011111: data <= 10'h3ff; 
        10'b0010100000: data <= 10'h3ff; 
        10'b0010100001: data <= 10'h3fe; 
        10'b0010100010: data <= 10'h3fe; 
        10'b0010100011: data <= 10'h3fd; 
        10'b0010100100: data <= 10'h3ff; 
        10'b0010100101: data <= 10'h3ff; 
        10'b0010100110: data <= 10'h000; 
        10'b0010100111: data <= 10'h3ff; 
        10'b0010101000: data <= 10'h000; 
        10'b0010101001: data <= 10'h3ff; 
        10'b0010101010: data <= 10'h000; 
        10'b0010101011: data <= 10'h000; 
        10'b0010101100: data <= 10'h000; 
        10'b0010101101: data <= 10'h000; 
        10'b0010101110: data <= 10'h002; 
        10'b0010101111: data <= 10'h003; 
        10'b0010110000: data <= 10'h002; 
        10'b0010110001: data <= 10'h003; 
        10'b0010110010: data <= 10'h004; 
        10'b0010110011: data <= 10'h002; 
        10'b0010110100: data <= 10'h003; 
        10'b0010110101: data <= 10'h003; 
        10'b0010110110: data <= 10'h003; 
        10'b0010110111: data <= 10'h002; 
        10'b0010111000: data <= 10'h002; 
        10'b0010111001: data <= 10'h000; 
        10'b0010111010: data <= 10'h000; 
        10'b0010111011: data <= 10'h3ff; 
        10'b0010111100: data <= 10'h3ff; 
        10'b0010111101: data <= 10'h3fe; 
        10'b0010111110: data <= 10'h3fe; 
        10'b0010111111: data <= 10'h3fd; 
        10'b0011000000: data <= 10'h3fe; 
        10'b0011000001: data <= 10'h3ff; 
        10'b0011000010: data <= 10'h000; 
        10'b0011000011: data <= 10'h000; 
        10'b0011000100: data <= 10'h000; 
        10'b0011000101: data <= 10'h000; 
        10'b0011000110: data <= 10'h000; 
        10'b0011000111: data <= 10'h000; 
        10'b0011001000: data <= 10'h000; 
        10'b0011001001: data <= 10'h001; 
        10'b0011001010: data <= 10'h002; 
        10'b0011001011: data <= 10'h003; 
        10'b0011001100: data <= 10'h003; 
        10'b0011001101: data <= 10'h002; 
        10'b0011001110: data <= 10'h001; 
        10'b0011001111: data <= 10'h001; 
        10'b0011010000: data <= 10'h000; 
        10'b0011010001: data <= 10'h002; 
        10'b0011010010: data <= 10'h002; 
        10'b0011010011: data <= 10'h000; 
        10'b0011010100: data <= 10'h000; 
        10'b0011010101: data <= 10'h3fd; 
        10'b0011010110: data <= 10'h3ff; 
        10'b0011010111: data <= 10'h3ff; 
        10'b0011011000: data <= 10'h3ff; 
        10'b0011011001: data <= 10'h3ff; 
        10'b0011011010: data <= 10'h3ff; 
        10'b0011011011: data <= 10'h3fd; 
        10'b0011011100: data <= 10'h3fe; 
        10'b0011011101: data <= 10'h3ff; 
        10'b0011011110: data <= 10'h3ff; 
        10'b0011011111: data <= 10'h3ff; 
        10'b0011100000: data <= 10'h000; 
        10'b0011100001: data <= 10'h000; 
        10'b0011100010: data <= 10'h000; 
        10'b0011100011: data <= 10'h000; 
        10'b0011100100: data <= 10'h000; 
        10'b0011100101: data <= 10'h001; 
        10'b0011100110: data <= 10'h001; 
        10'b0011100111: data <= 10'h002; 
        10'b0011101000: data <= 10'h002; 
        10'b0011101001: data <= 10'h002; 
        10'b0011101010: data <= 10'h002; 
        10'b0011101011: data <= 10'h002; 
        10'b0011101100: data <= 10'h001; 
        10'b0011101101: data <= 10'h001; 
        10'b0011101110: data <= 10'h004; 
        10'b0011101111: data <= 10'h002; 
        10'b0011110000: data <= 10'h000; 
        10'b0011110001: data <= 10'h3ff; 
        10'b0011110010: data <= 10'h000; 
        10'b0011110011: data <= 10'h001; 
        10'b0011110100: data <= 10'h000; 
        10'b0011110101: data <= 10'h3ff; 
        10'b0011110110: data <= 10'h3ff; 
        10'b0011110111: data <= 10'h3fd; 
        10'b0011111000: data <= 10'h3fe; 
        10'b0011111001: data <= 10'h3ff; 
        10'b0011111010: data <= 10'h000; 
        10'b0011111011: data <= 10'h3ff; 
        10'b0011111100: data <= 10'h3ff; 
        10'b0011111101: data <= 10'h000; 
        10'b0011111110: data <= 10'h000; 
        10'b0011111111: data <= 10'h000; 
        10'b0100000000: data <= 10'h001; 
        10'b0100000001: data <= 10'h002; 
        10'b0100000010: data <= 10'h001; 
        10'b0100000011: data <= 10'h000; 
        10'b0100000100: data <= 10'h3ff; 
        10'b0100000101: data <= 10'h001; 
        10'b0100000110: data <= 10'h001; 
        10'b0100000111: data <= 10'h001; 
        10'b0100001000: data <= 10'h000; 
        10'b0100001001: data <= 10'h000; 
        10'b0100001010: data <= 10'h002; 
        10'b0100001011: data <= 10'h003; 
        10'b0100001100: data <= 10'h001; 
        10'b0100001101: data <= 10'h000; 
        10'b0100001110: data <= 10'h000; 
        10'b0100001111: data <= 10'h000; 
        10'b0100010000: data <= 10'h000; 
        10'b0100010001: data <= 10'h000; 
        10'b0100010010: data <= 10'h3ff; 
        10'b0100010011: data <= 10'h3fd; 
        10'b0100010100: data <= 10'h3fe; 
        10'b0100010101: data <= 10'h3ff; 
        10'b0100010110: data <= 10'h000; 
        10'b0100010111: data <= 10'h3ff; 
        10'b0100011000: data <= 10'h000; 
        10'b0100011001: data <= 10'h000; 
        10'b0100011010: data <= 10'h000; 
        10'b0100011011: data <= 10'h3ff; 
        10'b0100011100: data <= 10'h000; 
        10'b0100011101: data <= 10'h000; 
        10'b0100011110: data <= 10'h3ff; 
        10'b0100011111: data <= 10'h3fc; 
        10'b0100100000: data <= 10'h3fc; 
        10'b0100100001: data <= 10'h3fd; 
        10'b0100100010: data <= 10'h3fc; 
        10'b0100100011: data <= 10'h3fb; 
        10'b0100100100: data <= 10'h3fb; 
        10'b0100100101: data <= 10'h3fa; 
        10'b0100100110: data <= 10'h3fd; 
        10'b0100100111: data <= 10'h000; 
        10'b0100101000: data <= 10'h001; 
        10'b0100101001: data <= 10'h000; 
        10'b0100101010: data <= 10'h000; 
        10'b0100101011: data <= 10'h000; 
        10'b0100101100: data <= 10'h000; 
        10'b0100101101: data <= 10'h000; 
        10'b0100101110: data <= 10'h3ff; 
        10'b0100101111: data <= 10'h3fd; 
        10'b0100110000: data <= 10'h3fe; 
        10'b0100110001: data <= 10'h000; 
        10'b0100110010: data <= 10'h000; 
        10'b0100110011: data <= 10'h3ff; 
        10'b0100110100: data <= 10'h3ff; 
        10'b0100110101: data <= 10'h000; 
        10'b0100110110: data <= 10'h000; 
        10'b0100110111: data <= 10'h3ff; 
        10'b0100111000: data <= 10'h3ff; 
        10'b0100111001: data <= 10'h3fd; 
        10'b0100111010: data <= 10'h3fa; 
        10'b0100111011: data <= 10'h3f8; 
        10'b0100111100: data <= 10'h3f8; 
        10'b0100111101: data <= 10'h3f7; 
        10'b0100111110: data <= 10'h3f7; 
        10'b0100111111: data <= 10'h3f8; 
        10'b0101000000: data <= 10'h3f7; 
        10'b0101000001: data <= 10'h3f5; 
        10'b0101000010: data <= 10'h3f8; 
        10'b0101000011: data <= 10'h3fc; 
        10'b0101000100: data <= 10'h3ff; 
        10'b0101000101: data <= 10'h3ff; 
        10'b0101000110: data <= 10'h3ff; 
        10'b0101000111: data <= 10'h000; 
        10'b0101001000: data <= 10'h3ff; 
        10'b0101001001: data <= 10'h3ff; 
        10'b0101001010: data <= 10'h3fe; 
        10'b0101001011: data <= 10'h3ff; 
        10'b0101001100: data <= 10'h000; 
        10'b0101001101: data <= 10'h000; 
        10'b0101001110: data <= 10'h3ff; 
        10'b0101001111: data <= 10'h000; 
        10'b0101010000: data <= 10'h000; 
        10'b0101010001: data <= 10'h000; 
        10'b0101010010: data <= 10'h000; 
        10'b0101010011: data <= 10'h000; 
        10'b0101010100: data <= 10'h3fe; 
        10'b0101010101: data <= 10'h3fb; 
        10'b0101010110: data <= 10'h3f7; 
        10'b0101010111: data <= 10'h3f4; 
        10'b0101011000: data <= 10'h3f5; 
        10'b0101011001: data <= 10'h3f6; 
        10'b0101011010: data <= 10'h3f7; 
        10'b0101011011: data <= 10'h3f7; 
        10'b0101011100: data <= 10'h3f7; 
        10'b0101011101: data <= 10'h3f7; 
        10'b0101011110: data <= 10'h3f9; 
        10'b0101011111: data <= 10'h3fb; 
        10'b0101100000: data <= 10'h3fd; 
        10'b0101100001: data <= 10'h3fd; 
        10'b0101100010: data <= 10'h3fe; 
        10'b0101100011: data <= 10'h000; 
        10'b0101100100: data <= 10'h000; 
        10'b0101100101: data <= 10'h3ff; 
        10'b0101100110: data <= 10'h3fe; 
        10'b0101100111: data <= 10'h3fd; 
        10'b0101101000: data <= 10'h000; 
        10'b0101101001: data <= 10'h000; 
        10'b0101101010: data <= 10'h000; 
        10'b0101101011: data <= 10'h000; 
        10'b0101101100: data <= 10'h3ff; 
        10'b0101101101: data <= 10'h000; 
        10'b0101101110: data <= 10'h000; 
        10'b0101101111: data <= 10'h3ff; 
        10'b0101110000: data <= 10'h3fd; 
        10'b0101110001: data <= 10'h3fa; 
        10'b0101110010: data <= 10'h3f6; 
        10'b0101110011: data <= 10'h3f7; 
        10'b0101110100: data <= 10'h3f8; 
        10'b0101110101: data <= 10'h3fa; 
        10'b0101110110: data <= 10'h3fc; 
        10'b0101110111: data <= 10'h3fe; 
        10'b0101111000: data <= 10'h3fd; 
        10'b0101111001: data <= 10'h3ff; 
        10'b0101111010: data <= 10'h3fd; 
        10'b0101111011: data <= 10'h3fc; 
        10'b0101111100: data <= 10'h3fc; 
        10'b0101111101: data <= 10'h3fd; 
        10'b0101111110: data <= 10'h3fe; 
        10'b0101111111: data <= 10'h000; 
        10'b0110000000: data <= 10'h000; 
        10'b0110000001: data <= 10'h3ff; 
        10'b0110000010: data <= 10'h3fe; 
        10'b0110000011: data <= 10'h3fe; 
        10'b0110000100: data <= 10'h3ff; 
        10'b0110000101: data <= 10'h000; 
        10'b0110000110: data <= 10'h000; 
        10'b0110000111: data <= 10'h000; 
        10'b0110001000: data <= 10'h000; 
        10'b0110001001: data <= 10'h000; 
        10'b0110001010: data <= 10'h000; 
        10'b0110001011: data <= 10'h3ff; 
        10'b0110001100: data <= 10'h3ff; 
        10'b0110001101: data <= 10'h3fc; 
        10'b0110001110: data <= 10'h3fb; 
        10'b0110001111: data <= 10'h3fc; 
        10'b0110010000: data <= 10'h3fe; 
        10'b0110010001: data <= 10'h000; 
        10'b0110010010: data <= 10'h001; 
        10'b0110010011: data <= 10'h001; 
        10'b0110010100: data <= 10'h002; 
        10'b0110010101: data <= 10'h003; 
        10'b0110010110: data <= 10'h000; 
        10'b0110010111: data <= 10'h3fe; 
        10'b0110011000: data <= 10'h3ff; 
        10'b0110011001: data <= 10'h3fe; 
        10'b0110011010: data <= 10'h000; 
        10'b0110011011: data <= 10'h3ff; 
        10'b0110011100: data <= 10'h000; 
        10'b0110011101: data <= 10'h3fe; 
        10'b0110011110: data <= 10'h3fd; 
        10'b0110011111: data <= 10'h3fe; 
        10'b0110100000: data <= 10'h000; 
        10'b0110100001: data <= 10'h001; 
        10'b0110100010: data <= 10'h001; 
        10'b0110100011: data <= 10'h3ff; 
        10'b0110100100: data <= 10'h000; 
        10'b0110100101: data <= 10'h000; 
        10'b0110100110: data <= 10'h000; 
        10'b0110100111: data <= 10'h001; 
        10'b0110101000: data <= 10'h000; 
        10'b0110101001: data <= 10'h000; 
        10'b0110101010: data <= 10'h001; 
        10'b0110101011: data <= 10'h001; 
        10'b0110101100: data <= 10'h002; 
        10'b0110101101: data <= 10'h002; 
        10'b0110101110: data <= 10'h002; 
        10'b0110101111: data <= 10'h001; 
        10'b0110110000: data <= 10'h001; 
        10'b0110110001: data <= 10'h003; 
        10'b0110110010: data <= 10'h000; 
        10'b0110110011: data <= 10'h001; 
        10'b0110110100: data <= 10'h000; 
        10'b0110110101: data <= 10'h3fe; 
        10'b0110110110: data <= 10'h3fe; 
        10'b0110110111: data <= 10'h3ff; 
        10'b0110111000: data <= 10'h3ff; 
        10'b0110111001: data <= 10'h3ff; 
        10'b0110111010: data <= 10'h3fd; 
        10'b0110111011: data <= 10'h3ff; 
        10'b0110111100: data <= 10'h001; 
        10'b0110111101: data <= 10'h001; 
        10'b0110111110: data <= 10'h001; 
        10'b0110111111: data <= 10'h3ff; 
        10'b0111000000: data <= 10'h3ff; 
        10'b0111000001: data <= 10'h3ff; 
        10'b0111000010: data <= 10'h3ff; 
        10'b0111000011: data <= 10'h001; 
        10'b0111000100: data <= 10'h002; 
        10'b0111000101: data <= 10'h003; 
        10'b0111000110: data <= 10'h004; 
        10'b0111000111: data <= 10'h002; 
        10'b0111001000: data <= 10'h001; 
        10'b0111001001: data <= 10'h002; 
        10'b0111001010: data <= 10'h002; 
        10'b0111001011: data <= 10'h002; 
        10'b0111001100: data <= 10'h003; 
        10'b0111001101: data <= 10'h003; 
        10'b0111001110: data <= 10'h001; 
        10'b0111001111: data <= 10'h000; 
        10'b0111010000: data <= 10'h000; 
        10'b0111010001: data <= 10'h3ff; 
        10'b0111010010: data <= 10'h3ff; 
        10'b0111010011: data <= 10'h3fe; 
        10'b0111010100: data <= 10'h3ff; 
        10'b0111010101: data <= 10'h000; 
        10'b0111010110: data <= 10'h000; 
        10'b0111010111: data <= 10'h001; 
        10'b0111011000: data <= 10'h003; 
        10'b0111011001: data <= 10'h004; 
        10'b0111011010: data <= 10'h001; 
        10'b0111011011: data <= 10'h3ff; 
        10'b0111011100: data <= 10'h000; 
        10'b0111011101: data <= 10'h000; 
        10'b0111011110: data <= 10'h000; 
        10'b0111011111: data <= 10'h001; 
        10'b0111100000: data <= 10'h004; 
        10'b0111100001: data <= 10'h005; 
        10'b0111100010: data <= 10'h005; 
        10'b0111100011: data <= 10'h003; 
        10'b0111100100: data <= 10'h002; 
        10'b0111100101: data <= 10'h003; 
        10'b0111100110: data <= 10'h004; 
        10'b0111100111: data <= 10'h003; 
        10'b0111101000: data <= 10'h004; 
        10'b0111101001: data <= 10'h002; 
        10'b0111101010: data <= 10'h001; 
        10'b0111101011: data <= 10'h001; 
        10'b0111101100: data <= 10'h001; 
        10'b0111101101: data <= 10'h000; 
        10'b0111101110: data <= 10'h001; 
        10'b0111101111: data <= 10'h3ff; 
        10'b0111110000: data <= 10'h002; 
        10'b0111110001: data <= 10'h002; 
        10'b0111110010: data <= 10'h001; 
        10'b0111110011: data <= 10'h002; 
        10'b0111110100: data <= 10'h005; 
        10'b0111110101: data <= 10'h004; 
        10'b0111110110: data <= 10'h001; 
        10'b0111110111: data <= 10'h000; 
        10'b0111111000: data <= 10'h000; 
        10'b0111111001: data <= 10'h000; 
        10'b0111111010: data <= 10'h3ff; 
        10'b0111111011: data <= 10'h000; 
        10'b0111111100: data <= 10'h004; 
        10'b0111111101: data <= 10'h007; 
        10'b0111111110: data <= 10'h006; 
        10'b0111111111: data <= 10'h004; 
        10'b1000000000: data <= 10'h003; 
        10'b1000000001: data <= 10'h003; 
        10'b1000000010: data <= 10'h005; 
        10'b1000000011: data <= 10'h005; 
        10'b1000000100: data <= 10'h007; 
        10'b1000000101: data <= 10'h005; 
        10'b1000000110: data <= 10'h005; 
        10'b1000000111: data <= 10'h002; 
        10'b1000001000: data <= 10'h002; 
        10'b1000001001: data <= 10'h003; 
        10'b1000001010: data <= 10'h002; 
        10'b1000001011: data <= 10'h001; 
        10'b1000001100: data <= 10'h003; 
        10'b1000001101: data <= 10'h003; 
        10'b1000001110: data <= 10'h004; 
        10'b1000001111: data <= 10'h005; 
        10'b1000010000: data <= 10'h006; 
        10'b1000010001: data <= 10'h004; 
        10'b1000010010: data <= 10'h000; 
        10'b1000010011: data <= 10'h3ff; 
        10'b1000010100: data <= 10'h3ff; 
        10'b1000010101: data <= 10'h3ff; 
        10'b1000010110: data <= 10'h3ff; 
        10'b1000010111: data <= 10'h000; 
        10'b1000011000: data <= 10'h002; 
        10'b1000011001: data <= 10'h004; 
        10'b1000011010: data <= 10'h005; 
        10'b1000011011: data <= 10'h004; 
        10'b1000011100: data <= 10'h004; 
        10'b1000011101: data <= 10'h004; 
        10'b1000011110: data <= 10'h004; 
        10'b1000011111: data <= 10'h004; 
        10'b1000100000: data <= 10'h005; 
        10'b1000100001: data <= 10'h004; 
        10'b1000100010: data <= 10'h002; 
        10'b1000100011: data <= 10'h001; 
        10'b1000100100: data <= 10'h002; 
        10'b1000100101: data <= 10'h003; 
        10'b1000100110: data <= 10'h002; 
        10'b1000100111: data <= 10'h001; 
        10'b1000101000: data <= 10'h003; 
        10'b1000101001: data <= 10'h003; 
        10'b1000101010: data <= 10'h004; 
        10'b1000101011: data <= 10'h004; 
        10'b1000101100: data <= 10'h004; 
        10'b1000101101: data <= 10'h002; 
        10'b1000101110: data <= 10'h000; 
        10'b1000101111: data <= 10'h000; 
        10'b1000110000: data <= 10'h3ff; 
        10'b1000110001: data <= 10'h000; 
        10'b1000110010: data <= 10'h000; 
        10'b1000110011: data <= 10'h3ff; 
        10'b1000110100: data <= 10'h002; 
        10'b1000110101: data <= 10'h002; 
        10'b1000110110: data <= 10'h004; 
        10'b1000110111: data <= 10'h005; 
        10'b1000111000: data <= 10'h005; 
        10'b1000111001: data <= 10'h003; 
        10'b1000111010: data <= 10'h003; 
        10'b1000111011: data <= 10'h005; 
        10'b1000111100: data <= 10'h003; 
        10'b1000111101: data <= 10'h001; 
        10'b1000111110: data <= 10'h001; 
        10'b1000111111: data <= 10'h001; 
        10'b1001000000: data <= 10'h001; 
        10'b1001000001: data <= 10'h000; 
        10'b1001000010: data <= 10'h002; 
        10'b1001000011: data <= 10'h003; 
        10'b1001000100: data <= 10'h002; 
        10'b1001000101: data <= 10'h003; 
        10'b1001000110: data <= 10'h005; 
        10'b1001000111: data <= 10'h004; 
        10'b1001001000: data <= 10'h003; 
        10'b1001001001: data <= 10'h001; 
        10'b1001001010: data <= 10'h000; 
        10'b1001001011: data <= 10'h000; 
        10'b1001001100: data <= 10'h000; 
        10'b1001001101: data <= 10'h3ff; 
        10'b1001001110: data <= 10'h000; 
        10'b1001001111: data <= 10'h000; 
        10'b1001010000: data <= 10'h000; 
        10'b1001010001: data <= 10'h001; 
        10'b1001010010: data <= 10'h003; 
        10'b1001010011: data <= 10'h003; 
        10'b1001010100: data <= 10'h003; 
        10'b1001010101: data <= 10'h003; 
        10'b1001010110: data <= 10'h003; 
        10'b1001010111: data <= 10'h003; 
        10'b1001011000: data <= 10'h001; 
        10'b1001011001: data <= 10'h001; 
        10'b1001011010: data <= 10'h000; 
        10'b1001011011: data <= 10'h000; 
        10'b1001011100: data <= 10'h001; 
        10'b1001011101: data <= 10'h001; 
        10'b1001011110: data <= 10'h003; 
        10'b1001011111: data <= 10'h003; 
        10'b1001100000: data <= 10'h002; 
        10'b1001100001: data <= 10'h003; 
        10'b1001100010: data <= 10'h004; 
        10'b1001100011: data <= 10'h005; 
        10'b1001100100: data <= 10'h002; 
        10'b1001100101: data <= 10'h001; 
        10'b1001100110: data <= 10'h000; 
        10'b1001100111: data <= 10'h000; 
        10'b1001101000: data <= 10'h3ff; 
        10'b1001101001: data <= 10'h000; 
        10'b1001101010: data <= 10'h3ff; 
        10'b1001101011: data <= 10'h000; 
        10'b1001101100: data <= 10'h001; 
        10'b1001101101: data <= 10'h000; 
        10'b1001101110: data <= 10'h002; 
        10'b1001101111: data <= 10'h002; 
        10'b1001110000: data <= 10'h001; 
        10'b1001110001: data <= 10'h002; 
        10'b1001110010: data <= 10'h002; 
        10'b1001110011: data <= 10'h002; 
        10'b1001110100: data <= 10'h000; 
        10'b1001110101: data <= 10'h3fe; 
        10'b1001110110: data <= 10'h3fe; 
        10'b1001110111: data <= 10'h3ff; 
        10'b1001111000: data <= 10'h3ff; 
        10'b1001111001: data <= 10'h001; 
        10'b1001111010: data <= 10'h003; 
        10'b1001111011: data <= 10'h004; 
        10'b1001111100: data <= 10'h004; 
        10'b1001111101: data <= 10'h003; 
        10'b1001111110: data <= 10'h003; 
        10'b1001111111: data <= 10'h003; 
        10'b1010000000: data <= 10'h001; 
        10'b1010000001: data <= 10'h000; 
        10'b1010000010: data <= 10'h000; 
        10'b1010000011: data <= 10'h3ff; 
        10'b1010000100: data <= 10'h000; 
        10'b1010000101: data <= 10'h000; 
        10'b1010000110: data <= 10'h000; 
        10'b1010000111: data <= 10'h000; 
        10'b1010001000: data <= 10'h000; 
        10'b1010001001: data <= 10'h3ff; 
        10'b1010001010: data <= 10'h3ff; 
        10'b1010001011: data <= 10'h3ff; 
        10'b1010001100: data <= 10'h3fe; 
        10'b1010001101: data <= 10'h3ff; 
        10'b1010001110: data <= 10'h3ff; 
        10'b1010001111: data <= 10'h001; 
        10'b1010010000: data <= 10'h000; 
        10'b1010010001: data <= 10'h3ff; 
        10'b1010010010: data <= 10'h3fe; 
        10'b1010010011: data <= 10'h3fe; 
        10'b1010010100: data <= 10'h3fe; 
        10'b1010010101: data <= 10'h3ff; 
        10'b1010010110: data <= 10'h000; 
        10'b1010010111: data <= 10'h003; 
        10'b1010011000: data <= 10'h003; 
        10'b1010011001: data <= 10'h003; 
        10'b1010011010: data <= 10'h002; 
        10'b1010011011: data <= 10'h001; 
        10'b1010011100: data <= 10'h001; 
        10'b1010011101: data <= 10'h000; 
        10'b1010011110: data <= 10'h000; 
        10'b1010011111: data <= 10'h000; 
        10'b1010100000: data <= 10'h000; 
        10'b1010100001: data <= 10'h3ff; 
        10'b1010100010: data <= 10'h000; 
        10'b1010100011: data <= 10'h000; 
        10'b1010100100: data <= 10'h3ff; 
        10'b1010100101: data <= 10'h3fe; 
        10'b1010100110: data <= 10'h3fd; 
        10'b1010100111: data <= 10'h3fe; 
        10'b1010101000: data <= 10'h3fd; 
        10'b1010101001: data <= 10'h3fd; 
        10'b1010101010: data <= 10'h3fd; 
        10'b1010101011: data <= 10'h3fe; 
        10'b1010101100: data <= 10'h3fe; 
        10'b1010101101: data <= 10'h3ff; 
        10'b1010101110: data <= 10'h3ff; 
        10'b1010101111: data <= 10'h3fe; 
        10'b1010110000: data <= 10'h3fe; 
        10'b1010110001: data <= 10'h3fe; 
        10'b1010110010: data <= 10'h3fe; 
        10'b1010110011: data <= 10'h3ff; 
        10'b1010110100: data <= 10'h3ff; 
        10'b1010110101: data <= 10'h3ff; 
        10'b1010110110: data <= 10'h3ff; 
        10'b1010110111: data <= 10'h000; 
        10'b1010111000: data <= 10'h000; 
        10'b1010111001: data <= 10'h000; 
        10'b1010111010: data <= 10'h3ff; 
        10'b1010111011: data <= 10'h3ff; 
        10'b1010111100: data <= 10'h000; 
        10'b1010111101: data <= 10'h3ff; 
        10'b1010111110: data <= 10'h000; 
        10'b1010111111: data <= 10'h3ff; 
        10'b1011000000: data <= 10'h3ff; 
        10'b1011000001: data <= 10'h3ff; 
        10'b1011000010: data <= 10'h3fe; 
        10'b1011000011: data <= 10'h3fe; 
        10'b1011000100: data <= 10'h3fd; 
        10'b1011000101: data <= 10'h3fe; 
        10'b1011000110: data <= 10'h3fe; 
        10'b1011000111: data <= 10'h3fd; 
        10'b1011001000: data <= 10'h3fe; 
        10'b1011001001: data <= 10'h3fe; 
        10'b1011001010: data <= 10'h3fe; 
        10'b1011001011: data <= 10'h3fe; 
        10'b1011001100: data <= 10'h3ff; 
        10'b1011001101: data <= 10'h3ff; 
        10'b1011001110: data <= 10'h3ff; 
        10'b1011001111: data <= 10'h3ff; 
        10'b1011010000: data <= 10'h000; 
        10'b1011010001: data <= 10'h000; 
        10'b1011010010: data <= 10'h000; 
        10'b1011010011: data <= 10'h3ff; 
        10'b1011010100: data <= 10'h000; 
        10'b1011010101: data <= 10'h3ff; 
        10'b1011010110: data <= 10'h3ff; 
        10'b1011010111: data <= 10'h3ff; 
        10'b1011011000: data <= 10'h3ff; 
        10'b1011011001: data <= 10'h3ff; 
        10'b1011011010: data <= 10'h000; 
        10'b1011011011: data <= 10'h000; 
        10'b1011011100: data <= 10'h000; 
        10'b1011011101: data <= 10'h000; 
        10'b1011011110: data <= 10'h000; 
        10'b1011011111: data <= 10'h000; 
        10'b1011100000: data <= 10'h000; 
        10'b1011100001: data <= 10'h000; 
        10'b1011100010: data <= 10'h000; 
        10'b1011100011: data <= 10'h000; 
        10'b1011100100: data <= 10'h000; 
        10'b1011100101: data <= 10'h000; 
        10'b1011100110: data <= 10'h3ff; 
        10'b1011100111: data <= 10'h3ff; 
        10'b1011101000: data <= 10'h000; 
        10'b1011101001: data <= 10'h000; 
        10'b1011101010: data <= 10'h000; 
        10'b1011101011: data <= 10'h3ff; 
        10'b1011101100: data <= 10'h000; 
        10'b1011101101: data <= 10'h000; 
        10'b1011101110: data <= 10'h3ff; 
        10'b1011101111: data <= 10'h3ff; 
        10'b1011110000: data <= 10'h3ff; 
        10'b1011110001: data <= 10'h000; 
        10'b1011110010: data <= 10'h000; 
        10'b1011110011: data <= 10'h000; 
        10'b1011110100: data <= 10'h000; 
        10'b1011110101: data <= 10'h3ff; 
        10'b1011110110: data <= 10'h3ff; 
        10'b1011110111: data <= 10'h000; 
        10'b1011111000: data <= 10'h3ff; 
        10'b1011111001: data <= 10'h000; 
        10'b1011111010: data <= 10'h000; 
        10'b1011111011: data <= 10'h000; 
        10'b1011111100: data <= 10'h000; 
        10'b1011111101: data <= 10'h3ff; 
        10'b1011111110: data <= 10'h000; 
        10'b1011111111: data <= 10'h3ff; 
        10'b1100000000: data <= 10'h000; 
        10'b1100000001: data <= 10'h000; 
        10'b1100000010: data <= 10'h000; 
        10'b1100000011: data <= 10'h3ff; 
        10'b1100000100: data <= 10'h000; 
        10'b1100000101: data <= 10'h000; 
        10'b1100000110: data <= 10'h000; 
        10'b1100000111: data <= 10'h000; 
        10'b1100001000: data <= 10'h000; 
        10'b1100001001: data <= 10'h3ff; 
        10'b1100001010: data <= 10'h000; 
        10'b1100001011: data <= 10'h000; 
        10'b1100001100: data <= 10'h3ff; 
        10'b1100001101: data <= 10'h000; 
        10'b1100001110: data <= 10'h000; 
        10'b1100001111: data <= 10'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 5) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 11'h7fe; 
        10'b0000000001: data <= 11'h000; 
        10'b0000000010: data <= 11'h7ff; 
        10'b0000000011: data <= 11'h7ff; 
        10'b0000000100: data <= 11'h7ff; 
        10'b0000000101: data <= 11'h7ff; 
        10'b0000000110: data <= 11'h7ff; 
        10'b0000000111: data <= 11'h000; 
        10'b0000001000: data <= 11'h7fe; 
        10'b0000001001: data <= 11'h7ff; 
        10'b0000001010: data <= 11'h7fe; 
        10'b0000001011: data <= 11'h7ff; 
        10'b0000001100: data <= 11'h000; 
        10'b0000001101: data <= 11'h000; 
        10'b0000001110: data <= 11'h7fe; 
        10'b0000001111: data <= 11'h7ff; 
        10'b0000010000: data <= 11'h7ff; 
        10'b0000010001: data <= 11'h7ff; 
        10'b0000010010: data <= 11'h000; 
        10'b0000010011: data <= 11'h000; 
        10'b0000010100: data <= 11'h7ff; 
        10'b0000010101: data <= 11'h7ff; 
        10'b0000010110: data <= 11'h7ff; 
        10'b0000010111: data <= 11'h7fe; 
        10'b0000011000: data <= 11'h7fe; 
        10'b0000011001: data <= 11'h7ff; 
        10'b0000011010: data <= 11'h000; 
        10'b0000011011: data <= 11'h000; 
        10'b0000011100: data <= 11'h7ff; 
        10'b0000011101: data <= 11'h7ff; 
        10'b0000011110: data <= 11'h000; 
        10'b0000011111: data <= 11'h000; 
        10'b0000100000: data <= 11'h7fe; 
        10'b0000100001: data <= 11'h7fe; 
        10'b0000100010: data <= 11'h7fe; 
        10'b0000100011: data <= 11'h7ff; 
        10'b0000100100: data <= 11'h7ff; 
        10'b0000100101: data <= 11'h7ff; 
        10'b0000100110: data <= 11'h000; 
        10'b0000100111: data <= 11'h7ff; 
        10'b0000101000: data <= 11'h7ff; 
        10'b0000101001: data <= 11'h7fe; 
        10'b0000101010: data <= 11'h7ff; 
        10'b0000101011: data <= 11'h7fe; 
        10'b0000101100: data <= 11'h000; 
        10'b0000101101: data <= 11'h7ff; 
        10'b0000101110: data <= 11'h7ff; 
        10'b0000101111: data <= 11'h7ff; 
        10'b0000110000: data <= 11'h7ff; 
        10'b0000110001: data <= 11'h7ff; 
        10'b0000110010: data <= 11'h7fe; 
        10'b0000110011: data <= 11'h7fe; 
        10'b0000110100: data <= 11'h000; 
        10'b0000110101: data <= 11'h000; 
        10'b0000110110: data <= 11'h000; 
        10'b0000110111: data <= 11'h7ff; 
        10'b0000111000: data <= 11'h7ff; 
        10'b0000111001: data <= 11'h7fe; 
        10'b0000111010: data <= 11'h7fe; 
        10'b0000111011: data <= 11'h000; 
        10'b0000111100: data <= 11'h7fe; 
        10'b0000111101: data <= 11'h7fe; 
        10'b0000111110: data <= 11'h7ff; 
        10'b0000111111: data <= 11'h7ff; 
        10'b0001000000: data <= 11'h000; 
        10'b0001000001: data <= 11'h7ff; 
        10'b0001000010: data <= 11'h001; 
        10'b0001000011: data <= 11'h001; 
        10'b0001000100: data <= 11'h002; 
        10'b0001000101: data <= 11'h002; 
        10'b0001000110: data <= 11'h002; 
        10'b0001000111: data <= 11'h001; 
        10'b0001001000: data <= 11'h002; 
        10'b0001001001: data <= 11'h001; 
        10'b0001001010: data <= 11'h001; 
        10'b0001001011: data <= 11'h7ff; 
        10'b0001001100: data <= 11'h000; 
        10'b0001001101: data <= 11'h7ff; 
        10'b0001001110: data <= 11'h7fe; 
        10'b0001001111: data <= 11'h7ff; 
        10'b0001010000: data <= 11'h000; 
        10'b0001010001: data <= 11'h001; 
        10'b0001010010: data <= 11'h7ff; 
        10'b0001010011: data <= 11'h7ff; 
        10'b0001010100: data <= 11'h7ff; 
        10'b0001010101: data <= 11'h7ff; 
        10'b0001010110: data <= 11'h000; 
        10'b0001010111: data <= 11'h7ff; 
        10'b0001011000: data <= 11'h000; 
        10'b0001011001: data <= 11'h7ff; 
        10'b0001011010: data <= 11'h7ff; 
        10'b0001011011: data <= 11'h000; 
        10'b0001011100: data <= 11'h000; 
        10'b0001011101: data <= 11'h004; 
        10'b0001011110: data <= 11'h006; 
        10'b0001011111: data <= 11'h006; 
        10'b0001100000: data <= 11'h005; 
        10'b0001100001: data <= 11'h008; 
        10'b0001100010: data <= 11'h004; 
        10'b0001100011: data <= 11'h002; 
        10'b0001100100: data <= 11'h004; 
        10'b0001100101: data <= 11'h002; 
        10'b0001100110: data <= 11'h7fe; 
        10'b0001100111: data <= 11'h000; 
        10'b0001101000: data <= 11'h7fe; 
        10'b0001101001: data <= 11'h7fe; 
        10'b0001101010: data <= 11'h7fd; 
        10'b0001101011: data <= 11'h7ff; 
        10'b0001101100: data <= 11'h000; 
        10'b0001101101: data <= 11'h001; 
        10'b0001101110: data <= 11'h7ff; 
        10'b0001101111: data <= 11'h000; 
        10'b0001110000: data <= 11'h7ff; 
        10'b0001110001: data <= 11'h7ff; 
        10'b0001110010: data <= 11'h000; 
        10'b0001110011: data <= 11'h7fe; 
        10'b0001110100: data <= 11'h7fe; 
        10'b0001110101: data <= 11'h7ff; 
        10'b0001110110: data <= 11'h001; 
        10'b0001110111: data <= 11'h001; 
        10'b0001111000: data <= 11'h002; 
        10'b0001111001: data <= 11'h007; 
        10'b0001111010: data <= 11'h007; 
        10'b0001111011: data <= 11'h009; 
        10'b0001111100: data <= 11'h008; 
        10'b0001111101: data <= 11'h006; 
        10'b0001111110: data <= 11'h005; 
        10'b0001111111: data <= 11'h002; 
        10'b0010000000: data <= 11'h003; 
        10'b0010000001: data <= 11'h003; 
        10'b0010000010: data <= 11'h7ff; 
        10'b0010000011: data <= 11'h7fe; 
        10'b0010000100: data <= 11'h7ff; 
        10'b0010000101: data <= 11'h7fc; 
        10'b0010000110: data <= 11'h7fc; 
        10'b0010000111: data <= 11'h7fc; 
        10'b0010001000: data <= 11'h7ff; 
        10'b0010001001: data <= 11'h7ff; 
        10'b0010001010: data <= 11'h7fe; 
        10'b0010001011: data <= 11'h000; 
        10'b0010001100: data <= 11'h000; 
        10'b0010001101: data <= 11'h7ff; 
        10'b0010001110: data <= 11'h7ff; 
        10'b0010001111: data <= 11'h7fe; 
        10'b0010010000: data <= 11'h7ff; 
        10'b0010010001: data <= 11'h7ff; 
        10'b0010010010: data <= 11'h001; 
        10'b0010010011: data <= 11'h003; 
        10'b0010010100: data <= 11'h005; 
        10'b0010010101: data <= 11'h008; 
        10'b0010010110: data <= 11'h009; 
        10'b0010010111: data <= 11'h009; 
        10'b0010011000: data <= 11'h009; 
        10'b0010011001: data <= 11'h00a; 
        10'b0010011010: data <= 11'h009; 
        10'b0010011011: data <= 11'h008; 
        10'b0010011100: data <= 11'h009; 
        10'b0010011101: data <= 11'h007; 
        10'b0010011110: data <= 11'h005; 
        10'b0010011111: data <= 11'h7fe; 
        10'b0010100000: data <= 11'h7fe; 
        10'b0010100001: data <= 11'h7fc; 
        10'b0010100010: data <= 11'h7fc; 
        10'b0010100011: data <= 11'h7fa; 
        10'b0010100100: data <= 11'h7fe; 
        10'b0010100101: data <= 11'h7ff; 
        10'b0010100110: data <= 11'h000; 
        10'b0010100111: data <= 11'h7ff; 
        10'b0010101000: data <= 11'h7ff; 
        10'b0010101001: data <= 11'h7ff; 
        10'b0010101010: data <= 11'h000; 
        10'b0010101011: data <= 11'h7ff; 
        10'b0010101100: data <= 11'h7ff; 
        10'b0010101101: data <= 11'h001; 
        10'b0010101110: data <= 11'h003; 
        10'b0010101111: data <= 11'h007; 
        10'b0010110000: data <= 11'h005; 
        10'b0010110001: data <= 11'h006; 
        10'b0010110010: data <= 11'h008; 
        10'b0010110011: data <= 11'h005; 
        10'b0010110100: data <= 11'h005; 
        10'b0010110101: data <= 11'h007; 
        10'b0010110110: data <= 11'h006; 
        10'b0010110111: data <= 11'h003; 
        10'b0010111000: data <= 11'h003; 
        10'b0010111001: data <= 11'h001; 
        10'b0010111010: data <= 11'h001; 
        10'b0010111011: data <= 11'h7fe; 
        10'b0010111100: data <= 11'h7ff; 
        10'b0010111101: data <= 11'h7fc; 
        10'b0010111110: data <= 11'h7fc; 
        10'b0010111111: data <= 11'h7fa; 
        10'b0011000000: data <= 11'h7fc; 
        10'b0011000001: data <= 11'h7fe; 
        10'b0011000010: data <= 11'h000; 
        10'b0011000011: data <= 11'h000; 
        10'b0011000100: data <= 11'h7ff; 
        10'b0011000101: data <= 11'h000; 
        10'b0011000110: data <= 11'h000; 
        10'b0011000111: data <= 11'h7ff; 
        10'b0011001000: data <= 11'h000; 
        10'b0011001001: data <= 11'h002; 
        10'b0011001010: data <= 11'h004; 
        10'b0011001011: data <= 11'h006; 
        10'b0011001100: data <= 11'h005; 
        10'b0011001101: data <= 11'h005; 
        10'b0011001110: data <= 11'h002; 
        10'b0011001111: data <= 11'h002; 
        10'b0011010000: data <= 11'h000; 
        10'b0011010001: data <= 11'h003; 
        10'b0011010010: data <= 11'h004; 
        10'b0011010011: data <= 11'h001; 
        10'b0011010100: data <= 11'h001; 
        10'b0011010101: data <= 11'h7fb; 
        10'b0011010110: data <= 11'h7fe; 
        10'b0011010111: data <= 11'h7ff; 
        10'b0011011000: data <= 11'h7fe; 
        10'b0011011001: data <= 11'h7fe; 
        10'b0011011010: data <= 11'h7ff; 
        10'b0011011011: data <= 11'h7fb; 
        10'b0011011100: data <= 11'h7fc; 
        10'b0011011101: data <= 11'h7ff; 
        10'b0011011110: data <= 11'h7ff; 
        10'b0011011111: data <= 11'h7fe; 
        10'b0011100000: data <= 11'h000; 
        10'b0011100001: data <= 11'h000; 
        10'b0011100010: data <= 11'h7ff; 
        10'b0011100011: data <= 11'h000; 
        10'b0011100100: data <= 11'h001; 
        10'b0011100101: data <= 11'h003; 
        10'b0011100110: data <= 11'h002; 
        10'b0011100111: data <= 11'h003; 
        10'b0011101000: data <= 11'h003; 
        10'b0011101001: data <= 11'h003; 
        10'b0011101010: data <= 11'h003; 
        10'b0011101011: data <= 11'h004; 
        10'b0011101100: data <= 11'h002; 
        10'b0011101101: data <= 11'h003; 
        10'b0011101110: data <= 11'h007; 
        10'b0011101111: data <= 11'h004; 
        10'b0011110000: data <= 11'h7ff; 
        10'b0011110001: data <= 11'h7fe; 
        10'b0011110010: data <= 11'h000; 
        10'b0011110011: data <= 11'h002; 
        10'b0011110100: data <= 11'h000; 
        10'b0011110101: data <= 11'h7ff; 
        10'b0011110110: data <= 11'h7fd; 
        10'b0011110111: data <= 11'h7fa; 
        10'b0011111000: data <= 11'h7fb; 
        10'b0011111001: data <= 11'h7fe; 
        10'b0011111010: data <= 11'h7ff; 
        10'b0011111011: data <= 11'h7ff; 
        10'b0011111100: data <= 11'h7ff; 
        10'b0011111101: data <= 11'h000; 
        10'b0011111110: data <= 11'h000; 
        10'b0011111111: data <= 11'h001; 
        10'b0100000000: data <= 11'h001; 
        10'b0100000001: data <= 11'h003; 
        10'b0100000010: data <= 11'h001; 
        10'b0100000011: data <= 11'h000; 
        10'b0100000100: data <= 11'h7ff; 
        10'b0100000101: data <= 11'h002; 
        10'b0100000110: data <= 11'h001; 
        10'b0100000111: data <= 11'h002; 
        10'b0100001000: data <= 11'h000; 
        10'b0100001001: data <= 11'h000; 
        10'b0100001010: data <= 11'h005; 
        10'b0100001011: data <= 11'h005; 
        10'b0100001100: data <= 11'h002; 
        10'b0100001101: data <= 11'h000; 
        10'b0100001110: data <= 11'h000; 
        10'b0100001111: data <= 11'h000; 
        10'b0100010000: data <= 11'h000; 
        10'b0100010001: data <= 11'h000; 
        10'b0100010010: data <= 11'h7fe; 
        10'b0100010011: data <= 11'h7fb; 
        10'b0100010100: data <= 11'h7fc; 
        10'b0100010101: data <= 11'h7ff; 
        10'b0100010110: data <= 11'h000; 
        10'b0100010111: data <= 11'h7fe; 
        10'b0100011000: data <= 11'h000; 
        10'b0100011001: data <= 11'h000; 
        10'b0100011010: data <= 11'h7ff; 
        10'b0100011011: data <= 11'h7ff; 
        10'b0100011100: data <= 11'h000; 
        10'b0100011101: data <= 11'h7ff; 
        10'b0100011110: data <= 11'h7fe; 
        10'b0100011111: data <= 11'h7f8; 
        10'b0100100000: data <= 11'h7f9; 
        10'b0100100001: data <= 11'h7fb; 
        10'b0100100010: data <= 11'h7f8; 
        10'b0100100011: data <= 11'h7f7; 
        10'b0100100100: data <= 11'h7f5; 
        10'b0100100101: data <= 11'h7f4; 
        10'b0100100110: data <= 11'h7fb; 
        10'b0100100111: data <= 11'h001; 
        10'b0100101000: data <= 11'h001; 
        10'b0100101001: data <= 11'h000; 
        10'b0100101010: data <= 11'h001; 
        10'b0100101011: data <= 11'h7ff; 
        10'b0100101100: data <= 11'h7ff; 
        10'b0100101101: data <= 11'h7ff; 
        10'b0100101110: data <= 11'h7fd; 
        10'b0100101111: data <= 11'h7fa; 
        10'b0100110000: data <= 11'h7fd; 
        10'b0100110001: data <= 11'h000; 
        10'b0100110010: data <= 11'h000; 
        10'b0100110011: data <= 11'h7ff; 
        10'b0100110100: data <= 11'h7fe; 
        10'b0100110101: data <= 11'h000; 
        10'b0100110110: data <= 11'h000; 
        10'b0100110111: data <= 11'h7fe; 
        10'b0100111000: data <= 11'h7fd; 
        10'b0100111001: data <= 11'h7f9; 
        10'b0100111010: data <= 11'h7f5; 
        10'b0100111011: data <= 11'h7f0; 
        10'b0100111100: data <= 11'h7f1; 
        10'b0100111101: data <= 11'h7ee; 
        10'b0100111110: data <= 11'h7ee; 
        10'b0100111111: data <= 11'h7f0; 
        10'b0101000000: data <= 11'h7ef; 
        10'b0101000001: data <= 11'h7eb; 
        10'b0101000010: data <= 11'h7f0; 
        10'b0101000011: data <= 11'h7f8; 
        10'b0101000100: data <= 11'h7fd; 
        10'b0101000101: data <= 11'h7fe; 
        10'b0101000110: data <= 11'h7fe; 
        10'b0101000111: data <= 11'h000; 
        10'b0101001000: data <= 11'h7ff; 
        10'b0101001001: data <= 11'h7ff; 
        10'b0101001010: data <= 11'h7fc; 
        10'b0101001011: data <= 11'h7fd; 
        10'b0101001100: data <= 11'h000; 
        10'b0101001101: data <= 11'h7ff; 
        10'b0101001110: data <= 11'h7ff; 
        10'b0101001111: data <= 11'h000; 
        10'b0101010000: data <= 11'h7ff; 
        10'b0101010001: data <= 11'h000; 
        10'b0101010010: data <= 11'h000; 
        10'b0101010011: data <= 11'h7ff; 
        10'b0101010100: data <= 11'h7fd; 
        10'b0101010101: data <= 11'h7f6; 
        10'b0101010110: data <= 11'h7ed; 
        10'b0101010111: data <= 11'h7e9; 
        10'b0101011000: data <= 11'h7ea; 
        10'b0101011001: data <= 11'h7eb; 
        10'b0101011010: data <= 11'h7ed; 
        10'b0101011011: data <= 11'h7ee; 
        10'b0101011100: data <= 11'h7ef; 
        10'b0101011101: data <= 11'h7ee; 
        10'b0101011110: data <= 11'h7f1; 
        10'b0101011111: data <= 11'h7f6; 
        10'b0101100000: data <= 11'h7f9; 
        10'b0101100001: data <= 11'h7fa; 
        10'b0101100010: data <= 11'h7fd; 
        10'b0101100011: data <= 11'h000; 
        10'b0101100100: data <= 11'h000; 
        10'b0101100101: data <= 11'h7fe; 
        10'b0101100110: data <= 11'h7fc; 
        10'b0101100111: data <= 11'h7fa; 
        10'b0101101000: data <= 11'h7ff; 
        10'b0101101001: data <= 11'h7ff; 
        10'b0101101010: data <= 11'h000; 
        10'b0101101011: data <= 11'h000; 
        10'b0101101100: data <= 11'h7ff; 
        10'b0101101101: data <= 11'h7ff; 
        10'b0101101110: data <= 11'h000; 
        10'b0101101111: data <= 11'h7ff; 
        10'b0101110000: data <= 11'h7fb; 
        10'b0101110001: data <= 11'h7f4; 
        10'b0101110010: data <= 11'h7ec; 
        10'b0101110011: data <= 11'h7ee; 
        10'b0101110100: data <= 11'h7ef; 
        10'b0101110101: data <= 11'h7f5; 
        10'b0101110110: data <= 11'h7f8; 
        10'b0101110111: data <= 11'h7fc; 
        10'b0101111000: data <= 11'h7fa; 
        10'b0101111001: data <= 11'h7fd; 
        10'b0101111010: data <= 11'h7f9; 
        10'b0101111011: data <= 11'h7f9; 
        10'b0101111100: data <= 11'h7f8; 
        10'b0101111101: data <= 11'h7fa; 
        10'b0101111110: data <= 11'h7fd; 
        10'b0101111111: data <= 11'h7ff; 
        10'b0110000000: data <= 11'h7ff; 
        10'b0110000001: data <= 11'h7fe; 
        10'b0110000010: data <= 11'h7fb; 
        10'b0110000011: data <= 11'h7fb; 
        10'b0110000100: data <= 11'h7fe; 
        10'b0110000101: data <= 11'h001; 
        10'b0110000110: data <= 11'h7ff; 
        10'b0110000111: data <= 11'h000; 
        10'b0110001000: data <= 11'h000; 
        10'b0110001001: data <= 11'h000; 
        10'b0110001010: data <= 11'h000; 
        10'b0110001011: data <= 11'h7ff; 
        10'b0110001100: data <= 11'h7fe; 
        10'b0110001101: data <= 11'h7f8; 
        10'b0110001110: data <= 11'h7f5; 
        10'b0110001111: data <= 11'h7f7; 
        10'b0110010000: data <= 11'h7fd; 
        10'b0110010001: data <= 11'h7ff; 
        10'b0110010010: data <= 11'h002; 
        10'b0110010011: data <= 11'h003; 
        10'b0110010100: data <= 11'h003; 
        10'b0110010101: data <= 11'h005; 
        10'b0110010110: data <= 11'h000; 
        10'b0110010111: data <= 11'h7fd; 
        10'b0110011000: data <= 11'h7fe; 
        10'b0110011001: data <= 11'h7fc; 
        10'b0110011010: data <= 11'h7ff; 
        10'b0110011011: data <= 11'h7fd; 
        10'b0110011100: data <= 11'h7ff; 
        10'b0110011101: data <= 11'h7fd; 
        10'b0110011110: data <= 11'h7fa; 
        10'b0110011111: data <= 11'h7fc; 
        10'b0110100000: data <= 11'h7ff; 
        10'b0110100001: data <= 11'h002; 
        10'b0110100010: data <= 11'h002; 
        10'b0110100011: data <= 11'h7ff; 
        10'b0110100100: data <= 11'h7ff; 
        10'b0110100101: data <= 11'h7ff; 
        10'b0110100110: data <= 11'h7ff; 
        10'b0110100111: data <= 11'h002; 
        10'b0110101000: data <= 11'h001; 
        10'b0110101001: data <= 11'h000; 
        10'b0110101010: data <= 11'h002; 
        10'b0110101011: data <= 11'h003; 
        10'b0110101100: data <= 11'h005; 
        10'b0110101101: data <= 11'h003; 
        10'b0110101110: data <= 11'h004; 
        10'b0110101111: data <= 11'h002; 
        10'b0110110000: data <= 11'h002; 
        10'b0110110001: data <= 11'h005; 
        10'b0110110010: data <= 11'h000; 
        10'b0110110011: data <= 11'h002; 
        10'b0110110100: data <= 11'h000; 
        10'b0110110101: data <= 11'h7fc; 
        10'b0110110110: data <= 11'h7fc; 
        10'b0110110111: data <= 11'h7fe; 
        10'b0110111000: data <= 11'h7fe; 
        10'b0110111001: data <= 11'h7fd; 
        10'b0110111010: data <= 11'h7fb; 
        10'b0110111011: data <= 11'h7fd; 
        10'b0110111100: data <= 11'h002; 
        10'b0110111101: data <= 11'h003; 
        10'b0110111110: data <= 11'h001; 
        10'b0110111111: data <= 11'h7ff; 
        10'b0111000000: data <= 11'h7ff; 
        10'b0111000001: data <= 11'h7fe; 
        10'b0111000010: data <= 11'h7fe; 
        10'b0111000011: data <= 11'h002; 
        10'b0111000100: data <= 11'h004; 
        10'b0111000101: data <= 11'h007; 
        10'b0111000110: data <= 11'h007; 
        10'b0111000111: data <= 11'h004; 
        10'b0111001000: data <= 11'h002; 
        10'b0111001001: data <= 11'h004; 
        10'b0111001010: data <= 11'h003; 
        10'b0111001011: data <= 11'h003; 
        10'b0111001100: data <= 11'h006; 
        10'b0111001101: data <= 11'h006; 
        10'b0111001110: data <= 11'h001; 
        10'b0111001111: data <= 11'h7ff; 
        10'b0111010000: data <= 11'h000; 
        10'b0111010001: data <= 11'h7fd; 
        10'b0111010010: data <= 11'h7fe; 
        10'b0111010011: data <= 11'h7fc; 
        10'b0111010100: data <= 11'h7ff; 
        10'b0111010101: data <= 11'h000; 
        10'b0111010110: data <= 11'h001; 
        10'b0111010111: data <= 11'h002; 
        10'b0111011000: data <= 11'h006; 
        10'b0111011001: data <= 11'h007; 
        10'b0111011010: data <= 11'h001; 
        10'b0111011011: data <= 11'h7ff; 
        10'b0111011100: data <= 11'h7ff; 
        10'b0111011101: data <= 11'h000; 
        10'b0111011110: data <= 11'h7ff; 
        10'b0111011111: data <= 11'h002; 
        10'b0111100000: data <= 11'h007; 
        10'b0111100001: data <= 11'h00a; 
        10'b0111100010: data <= 11'h009; 
        10'b0111100011: data <= 11'h006; 
        10'b0111100100: data <= 11'h004; 
        10'b0111100101: data <= 11'h005; 
        10'b0111100110: data <= 11'h008; 
        10'b0111100111: data <= 11'h007; 
        10'b0111101000: data <= 11'h008; 
        10'b0111101001: data <= 11'h004; 
        10'b0111101010: data <= 11'h002; 
        10'b0111101011: data <= 11'h003; 
        10'b0111101100: data <= 11'h003; 
        10'b0111101101: data <= 11'h000; 
        10'b0111101110: data <= 11'h002; 
        10'b0111101111: data <= 11'h7ff; 
        10'b0111110000: data <= 11'h003; 
        10'b0111110001: data <= 11'h003; 
        10'b0111110010: data <= 11'h002; 
        10'b0111110011: data <= 11'h003; 
        10'b0111110100: data <= 11'h009; 
        10'b0111110101: data <= 11'h008; 
        10'b0111110110: data <= 11'h002; 
        10'b0111110111: data <= 11'h000; 
        10'b0111111000: data <= 11'h000; 
        10'b0111111001: data <= 11'h000; 
        10'b0111111010: data <= 11'h7fe; 
        10'b0111111011: data <= 11'h001; 
        10'b0111111100: data <= 11'h008; 
        10'b0111111101: data <= 11'h00d; 
        10'b0111111110: data <= 11'h00c; 
        10'b0111111111: data <= 11'h009; 
        10'b1000000000: data <= 11'h006; 
        10'b1000000001: data <= 11'h007; 
        10'b1000000010: data <= 11'h00a; 
        10'b1000000011: data <= 11'h009; 
        10'b1000000100: data <= 11'h00f; 
        10'b1000000101: data <= 11'h00b; 
        10'b1000000110: data <= 11'h009; 
        10'b1000000111: data <= 11'h005; 
        10'b1000001000: data <= 11'h003; 
        10'b1000001001: data <= 11'h006; 
        10'b1000001010: data <= 11'h004; 
        10'b1000001011: data <= 11'h003; 
        10'b1000001100: data <= 11'h007; 
        10'b1000001101: data <= 11'h007; 
        10'b1000001110: data <= 11'h008; 
        10'b1000001111: data <= 11'h00a; 
        10'b1000010000: data <= 11'h00c; 
        10'b1000010001: data <= 11'h007; 
        10'b1000010010: data <= 11'h7ff; 
        10'b1000010011: data <= 11'h7ff; 
        10'b1000010100: data <= 11'h7ff; 
        10'b1000010101: data <= 11'h7ff; 
        10'b1000010110: data <= 11'h7fe; 
        10'b1000010111: data <= 11'h000; 
        10'b1000011000: data <= 11'h004; 
        10'b1000011001: data <= 11'h008; 
        10'b1000011010: data <= 11'h00a; 
        10'b1000011011: data <= 11'h009; 
        10'b1000011100: data <= 11'h008; 
        10'b1000011101: data <= 11'h009; 
        10'b1000011110: data <= 11'h008; 
        10'b1000011111: data <= 11'h009; 
        10'b1000100000: data <= 11'h00a; 
        10'b1000100001: data <= 11'h008; 
        10'b1000100010: data <= 11'h005; 
        10'b1000100011: data <= 11'h002; 
        10'b1000100100: data <= 11'h004; 
        10'b1000100101: data <= 11'h006; 
        10'b1000100110: data <= 11'h003; 
        10'b1000100111: data <= 11'h003; 
        10'b1000101000: data <= 11'h005; 
        10'b1000101001: data <= 11'h006; 
        10'b1000101010: data <= 11'h008; 
        10'b1000101011: data <= 11'h009; 
        10'b1000101100: data <= 11'h008; 
        10'b1000101101: data <= 11'h004; 
        10'b1000101110: data <= 11'h000; 
        10'b1000101111: data <= 11'h000; 
        10'b1000110000: data <= 11'h7fe; 
        10'b1000110001: data <= 11'h000; 
        10'b1000110010: data <= 11'h000; 
        10'b1000110011: data <= 11'h7fe; 
        10'b1000110100: data <= 11'h004; 
        10'b1000110101: data <= 11'h005; 
        10'b1000110110: data <= 11'h007; 
        10'b1000110111: data <= 11'h00a; 
        10'b1000111000: data <= 11'h00a; 
        10'b1000111001: data <= 11'h006; 
        10'b1000111010: data <= 11'h006; 
        10'b1000111011: data <= 11'h00a; 
        10'b1000111100: data <= 11'h006; 
        10'b1000111101: data <= 11'h002; 
        10'b1000111110: data <= 11'h001; 
        10'b1000111111: data <= 11'h002; 
        10'b1001000000: data <= 11'h002; 
        10'b1001000001: data <= 11'h000; 
        10'b1001000010: data <= 11'h004; 
        10'b1001000011: data <= 11'h007; 
        10'b1001000100: data <= 11'h005; 
        10'b1001000101: data <= 11'h007; 
        10'b1001000110: data <= 11'h009; 
        10'b1001000111: data <= 11'h008; 
        10'b1001001000: data <= 11'h006; 
        10'b1001001001: data <= 11'h003; 
        10'b1001001010: data <= 11'h000; 
        10'b1001001011: data <= 11'h000; 
        10'b1001001100: data <= 11'h7ff; 
        10'b1001001101: data <= 11'h7ff; 
        10'b1001001110: data <= 11'h000; 
        10'b1001001111: data <= 11'h7ff; 
        10'b1001010000: data <= 11'h001; 
        10'b1001010001: data <= 11'h002; 
        10'b1001010010: data <= 11'h005; 
        10'b1001010011: data <= 11'h006; 
        10'b1001010100: data <= 11'h005; 
        10'b1001010101: data <= 11'h006; 
        10'b1001010110: data <= 11'h006; 
        10'b1001010111: data <= 11'h005; 
        10'b1001011000: data <= 11'h002; 
        10'b1001011001: data <= 11'h001; 
        10'b1001011010: data <= 11'h7ff; 
        10'b1001011011: data <= 11'h000; 
        10'b1001011100: data <= 11'h003; 
        10'b1001011101: data <= 11'h003; 
        10'b1001011110: data <= 11'h007; 
        10'b1001011111: data <= 11'h007; 
        10'b1001100000: data <= 11'h003; 
        10'b1001100001: data <= 11'h007; 
        10'b1001100010: data <= 11'h008; 
        10'b1001100011: data <= 11'h009; 
        10'b1001100100: data <= 11'h005; 
        10'b1001100101: data <= 11'h002; 
        10'b1001100110: data <= 11'h000; 
        10'b1001100111: data <= 11'h000; 
        10'b1001101000: data <= 11'h7fe; 
        10'b1001101001: data <= 11'h000; 
        10'b1001101010: data <= 11'h7ff; 
        10'b1001101011: data <= 11'h000; 
        10'b1001101100: data <= 11'h002; 
        10'b1001101101: data <= 11'h001; 
        10'b1001101110: data <= 11'h003; 
        10'b1001101111: data <= 11'h003; 
        10'b1001110000: data <= 11'h003; 
        10'b1001110001: data <= 11'h004; 
        10'b1001110010: data <= 11'h004; 
        10'b1001110011: data <= 11'h005; 
        10'b1001110100: data <= 11'h001; 
        10'b1001110101: data <= 11'h7fc; 
        10'b1001110110: data <= 11'h7fb; 
        10'b1001110111: data <= 11'h7fd; 
        10'b1001111000: data <= 11'h7fe; 
        10'b1001111001: data <= 11'h002; 
        10'b1001111010: data <= 11'h006; 
        10'b1001111011: data <= 11'h008; 
        10'b1001111100: data <= 11'h007; 
        10'b1001111101: data <= 11'h007; 
        10'b1001111110: data <= 11'h006; 
        10'b1001111111: data <= 11'h006; 
        10'b1010000000: data <= 11'h002; 
        10'b1010000001: data <= 11'h000; 
        10'b1010000010: data <= 11'h000; 
        10'b1010000011: data <= 11'h7ff; 
        10'b1010000100: data <= 11'h000; 
        10'b1010000101: data <= 11'h000; 
        10'b1010000110: data <= 11'h7ff; 
        10'b1010000111: data <= 11'h7ff; 
        10'b1010001000: data <= 11'h7ff; 
        10'b1010001001: data <= 11'h7fe; 
        10'b1010001010: data <= 11'h7fe; 
        10'b1010001011: data <= 11'h7fe; 
        10'b1010001100: data <= 11'h7fd; 
        10'b1010001101: data <= 11'h7fe; 
        10'b1010001110: data <= 11'h7ff; 
        10'b1010001111: data <= 11'h002; 
        10'b1010010000: data <= 11'h000; 
        10'b1010010001: data <= 11'h7fe; 
        10'b1010010010: data <= 11'h7fd; 
        10'b1010010011: data <= 11'h7fc; 
        10'b1010010100: data <= 11'h7fb; 
        10'b1010010101: data <= 11'h7fe; 
        10'b1010010110: data <= 11'h001; 
        10'b1010010111: data <= 11'h006; 
        10'b1010011000: data <= 11'h005; 
        10'b1010011001: data <= 11'h006; 
        10'b1010011010: data <= 11'h005; 
        10'b1010011011: data <= 11'h002; 
        10'b1010011100: data <= 11'h001; 
        10'b1010011101: data <= 11'h001; 
        10'b1010011110: data <= 11'h000; 
        10'b1010011111: data <= 11'h7ff; 
        10'b1010100000: data <= 11'h7ff; 
        10'b1010100001: data <= 11'h7ff; 
        10'b1010100010: data <= 11'h000; 
        10'b1010100011: data <= 11'h000; 
        10'b1010100100: data <= 11'h7ff; 
        10'b1010100101: data <= 11'h7fd; 
        10'b1010100110: data <= 11'h7f9; 
        10'b1010100111: data <= 11'h7fb; 
        10'b1010101000: data <= 11'h7fb; 
        10'b1010101001: data <= 11'h7fb; 
        10'b1010101010: data <= 11'h7fb; 
        10'b1010101011: data <= 11'h7fc; 
        10'b1010101100: data <= 11'h7fc; 
        10'b1010101101: data <= 11'h7fe; 
        10'b1010101110: data <= 11'h7fd; 
        10'b1010101111: data <= 11'h7fc; 
        10'b1010110000: data <= 11'h7fc; 
        10'b1010110001: data <= 11'h7fd; 
        10'b1010110010: data <= 11'h7fc; 
        10'b1010110011: data <= 11'h7fe; 
        10'b1010110100: data <= 11'h7fe; 
        10'b1010110101: data <= 11'h7fe; 
        10'b1010110110: data <= 11'h7ff; 
        10'b1010110111: data <= 11'h7ff; 
        10'b1010111000: data <= 11'h000; 
        10'b1010111001: data <= 11'h001; 
        10'b1010111010: data <= 11'h7ff; 
        10'b1010111011: data <= 11'h7ff; 
        10'b1010111100: data <= 11'h000; 
        10'b1010111101: data <= 11'h7fe; 
        10'b1010111110: data <= 11'h7ff; 
        10'b1010111111: data <= 11'h7ff; 
        10'b1011000000: data <= 11'h7ff; 
        10'b1011000001: data <= 11'h7fe; 
        10'b1011000010: data <= 11'h7fd; 
        10'b1011000011: data <= 11'h7fb; 
        10'b1011000100: data <= 11'h7fb; 
        10'b1011000101: data <= 11'h7fb; 
        10'b1011000110: data <= 11'h7fb; 
        10'b1011000111: data <= 11'h7fa; 
        10'b1011001000: data <= 11'h7fc; 
        10'b1011001001: data <= 11'h7fc; 
        10'b1011001010: data <= 11'h7fb; 
        10'b1011001011: data <= 11'h7fc; 
        10'b1011001100: data <= 11'h7fd; 
        10'b1011001101: data <= 11'h7fd; 
        10'b1011001110: data <= 11'h7ff; 
        10'b1011001111: data <= 11'h7fd; 
        10'b1011010000: data <= 11'h7ff; 
        10'b1011010001: data <= 11'h7ff; 
        10'b1011010010: data <= 11'h000; 
        10'b1011010011: data <= 11'h7ff; 
        10'b1011010100: data <= 11'h7ff; 
        10'b1011010101: data <= 11'h7ff; 
        10'b1011010110: data <= 11'h7fe; 
        10'b1011010111: data <= 11'h7ff; 
        10'b1011011000: data <= 11'h7fe; 
        10'b1011011001: data <= 11'h7ff; 
        10'b1011011010: data <= 11'h7ff; 
        10'b1011011011: data <= 11'h000; 
        10'b1011011100: data <= 11'h000; 
        10'b1011011101: data <= 11'h7ff; 
        10'b1011011110: data <= 11'h000; 
        10'b1011011111: data <= 11'h000; 
        10'b1011100000: data <= 11'h7ff; 
        10'b1011100001: data <= 11'h000; 
        10'b1011100010: data <= 11'h000; 
        10'b1011100011: data <= 11'h000; 
        10'b1011100100: data <= 11'h000; 
        10'b1011100101: data <= 11'h7ff; 
        10'b1011100110: data <= 11'h7ff; 
        10'b1011100111: data <= 11'h7fe; 
        10'b1011101000: data <= 11'h7ff; 
        10'b1011101001: data <= 11'h7ff; 
        10'b1011101010: data <= 11'h7ff; 
        10'b1011101011: data <= 11'h7ff; 
        10'b1011101100: data <= 11'h000; 
        10'b1011101101: data <= 11'h000; 
        10'b1011101110: data <= 11'h7ff; 
        10'b1011101111: data <= 11'h7ff; 
        10'b1011110000: data <= 11'h7fe; 
        10'b1011110001: data <= 11'h000; 
        10'b1011110010: data <= 11'h000; 
        10'b1011110011: data <= 11'h000; 
        10'b1011110100: data <= 11'h000; 
        10'b1011110101: data <= 11'h7ff; 
        10'b1011110110: data <= 11'h7fe; 
        10'b1011110111: data <= 11'h7ff; 
        10'b1011111000: data <= 11'h7fe; 
        10'b1011111001: data <= 11'h000; 
        10'b1011111010: data <= 11'h000; 
        10'b1011111011: data <= 11'h7ff; 
        10'b1011111100: data <= 11'h000; 
        10'b1011111101: data <= 11'h7ff; 
        10'b1011111110: data <= 11'h000; 
        10'b1011111111: data <= 11'h7fe; 
        10'b1100000000: data <= 11'h000; 
        10'b1100000001: data <= 11'h7ff; 
        10'b1100000010: data <= 11'h000; 
        10'b1100000011: data <= 11'h7ff; 
        10'b1100000100: data <= 11'h7ff; 
        10'b1100000101: data <= 11'h7ff; 
        10'b1100000110: data <= 11'h7ff; 
        10'b1100000111: data <= 11'h7ff; 
        10'b1100001000: data <= 11'h000; 
        10'b1100001001: data <= 11'h7fe; 
        10'b1100001010: data <= 11'h7ff; 
        10'b1100001011: data <= 11'h000; 
        10'b1100001100: data <= 11'h7fe; 
        10'b1100001101: data <= 11'h7ff; 
        10'b1100001110: data <= 11'h000; 
        10'b1100001111: data <= 11'h7ff; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 6) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 12'hffd; 
        10'b0000000001: data <= 12'h000; 
        10'b0000000010: data <= 12'hffe; 
        10'b0000000011: data <= 12'hffd; 
        10'b0000000100: data <= 12'hffe; 
        10'b0000000101: data <= 12'hffe; 
        10'b0000000110: data <= 12'hfff; 
        10'b0000000111: data <= 12'hfff; 
        10'b0000001000: data <= 12'hffd; 
        10'b0000001001: data <= 12'hfff; 
        10'b0000001010: data <= 12'hffd; 
        10'b0000001011: data <= 12'hffe; 
        10'b0000001100: data <= 12'h001; 
        10'b0000001101: data <= 12'h001; 
        10'b0000001110: data <= 12'hffd; 
        10'b0000001111: data <= 12'hfff; 
        10'b0000010000: data <= 12'hffd; 
        10'b0000010001: data <= 12'hffd; 
        10'b0000010010: data <= 12'h001; 
        10'b0000010011: data <= 12'h000; 
        10'b0000010100: data <= 12'hffe; 
        10'b0000010101: data <= 12'hfff; 
        10'b0000010110: data <= 12'hffe; 
        10'b0000010111: data <= 12'hffc; 
        10'b0000011000: data <= 12'hffd; 
        10'b0000011001: data <= 12'hfff; 
        10'b0000011010: data <= 12'h000; 
        10'b0000011011: data <= 12'hfff; 
        10'b0000011100: data <= 12'hfff; 
        10'b0000011101: data <= 12'hffe; 
        10'b0000011110: data <= 12'h001; 
        10'b0000011111: data <= 12'hfff; 
        10'b0000100000: data <= 12'hffd; 
        10'b0000100001: data <= 12'hffd; 
        10'b0000100010: data <= 12'hffd; 
        10'b0000100011: data <= 12'hffe; 
        10'b0000100100: data <= 12'hffe; 
        10'b0000100101: data <= 12'hfff; 
        10'b0000100110: data <= 12'h000; 
        10'b0000100111: data <= 12'hffd; 
        10'b0000101000: data <= 12'hffe; 
        10'b0000101001: data <= 12'hffd; 
        10'b0000101010: data <= 12'hfff; 
        10'b0000101011: data <= 12'hffd; 
        10'b0000101100: data <= 12'hfff; 
        10'b0000101101: data <= 12'hffd; 
        10'b0000101110: data <= 12'hffe; 
        10'b0000101111: data <= 12'hffd; 
        10'b0000110000: data <= 12'hfff; 
        10'b0000110001: data <= 12'hffd; 
        10'b0000110010: data <= 12'hffd; 
        10'b0000110011: data <= 12'hffc; 
        10'b0000110100: data <= 12'h000; 
        10'b0000110101: data <= 12'hfff; 
        10'b0000110110: data <= 12'h000; 
        10'b0000110111: data <= 12'hffe; 
        10'b0000111000: data <= 12'hffe; 
        10'b0000111001: data <= 12'hffd; 
        10'b0000111010: data <= 12'hffd; 
        10'b0000111011: data <= 12'h000; 
        10'b0000111100: data <= 12'hffd; 
        10'b0000111101: data <= 12'hffd; 
        10'b0000111110: data <= 12'hffe; 
        10'b0000111111: data <= 12'hfff; 
        10'b0001000000: data <= 12'h000; 
        10'b0001000001: data <= 12'hffe; 
        10'b0001000010: data <= 12'h002; 
        10'b0001000011: data <= 12'h001; 
        10'b0001000100: data <= 12'h005; 
        10'b0001000101: data <= 12'h004; 
        10'b0001000110: data <= 12'h003; 
        10'b0001000111: data <= 12'h001; 
        10'b0001001000: data <= 12'h005; 
        10'b0001001001: data <= 12'h002; 
        10'b0001001010: data <= 12'h001; 
        10'b0001001011: data <= 12'hffe; 
        10'b0001001100: data <= 12'h000; 
        10'b0001001101: data <= 12'hfff; 
        10'b0001001110: data <= 12'hffb; 
        10'b0001001111: data <= 12'hffe; 
        10'b0001010000: data <= 12'h000; 
        10'b0001010001: data <= 12'h001; 
        10'b0001010010: data <= 12'hfff; 
        10'b0001010011: data <= 12'hffe; 
        10'b0001010100: data <= 12'hffe; 
        10'b0001010101: data <= 12'hffd; 
        10'b0001010110: data <= 12'hfff; 
        10'b0001010111: data <= 12'hffe; 
        10'b0001011000: data <= 12'h001; 
        10'b0001011001: data <= 12'hffd; 
        10'b0001011010: data <= 12'hfff; 
        10'b0001011011: data <= 12'h000; 
        10'b0001011100: data <= 12'h001; 
        10'b0001011101: data <= 12'h007; 
        10'b0001011110: data <= 12'h00c; 
        10'b0001011111: data <= 12'h00b; 
        10'b0001100000: data <= 12'h00b; 
        10'b0001100001: data <= 12'h010; 
        10'b0001100010: data <= 12'h009; 
        10'b0001100011: data <= 12'h004; 
        10'b0001100100: data <= 12'h007; 
        10'b0001100101: data <= 12'h003; 
        10'b0001100110: data <= 12'hffd; 
        10'b0001100111: data <= 12'hfff; 
        10'b0001101000: data <= 12'hffc; 
        10'b0001101001: data <= 12'hffc; 
        10'b0001101010: data <= 12'hffb; 
        10'b0001101011: data <= 12'hffd; 
        10'b0001101100: data <= 12'h000; 
        10'b0001101101: data <= 12'h001; 
        10'b0001101110: data <= 12'hffd; 
        10'b0001101111: data <= 12'hfff; 
        10'b0001110000: data <= 12'hffd; 
        10'b0001110001: data <= 12'hffe; 
        10'b0001110010: data <= 12'h001; 
        10'b0001110011: data <= 12'hffc; 
        10'b0001110100: data <= 12'hffd; 
        10'b0001110101: data <= 12'hfff; 
        10'b0001110110: data <= 12'h002; 
        10'b0001110111: data <= 12'h002; 
        10'b0001111000: data <= 12'h005; 
        10'b0001111001: data <= 12'h00e; 
        10'b0001111010: data <= 12'h00e; 
        10'b0001111011: data <= 12'h012; 
        10'b0001111100: data <= 12'h00f; 
        10'b0001111101: data <= 12'h00c; 
        10'b0001111110: data <= 12'h00b; 
        10'b0001111111: data <= 12'h005; 
        10'b0010000000: data <= 12'h006; 
        10'b0010000001: data <= 12'h006; 
        10'b0010000010: data <= 12'hffe; 
        10'b0010000011: data <= 12'hffd; 
        10'b0010000100: data <= 12'hffe; 
        10'b0010000101: data <= 12'hff9; 
        10'b0010000110: data <= 12'hff7; 
        10'b0010000111: data <= 12'hff8; 
        10'b0010001000: data <= 12'hfff; 
        10'b0010001001: data <= 12'hfff; 
        10'b0010001010: data <= 12'hffd; 
        10'b0010001011: data <= 12'hfff; 
        10'b0010001100: data <= 12'h000; 
        10'b0010001101: data <= 12'hfff; 
        10'b0010001110: data <= 12'hffd; 
        10'b0010001111: data <= 12'hffc; 
        10'b0010010000: data <= 12'hffd; 
        10'b0010010001: data <= 12'hffd; 
        10'b0010010010: data <= 12'h002; 
        10'b0010010011: data <= 12'h007; 
        10'b0010010100: data <= 12'h00a; 
        10'b0010010101: data <= 12'h010; 
        10'b0010010110: data <= 12'h012; 
        10'b0010010111: data <= 12'h013; 
        10'b0010011000: data <= 12'h011; 
        10'b0010011001: data <= 12'h013; 
        10'b0010011010: data <= 12'h012; 
        10'b0010011011: data <= 12'h011; 
        10'b0010011100: data <= 12'h012; 
        10'b0010011101: data <= 12'h00f; 
        10'b0010011110: data <= 12'h00b; 
        10'b0010011111: data <= 12'hffc; 
        10'b0010100000: data <= 12'hffc; 
        10'b0010100001: data <= 12'hff9; 
        10'b0010100010: data <= 12'hff9; 
        10'b0010100011: data <= 12'hff5; 
        10'b0010100100: data <= 12'hffb; 
        10'b0010100101: data <= 12'hffd; 
        10'b0010100110: data <= 12'h000; 
        10'b0010100111: data <= 12'hffe; 
        10'b0010101000: data <= 12'hfff; 
        10'b0010101001: data <= 12'hffd; 
        10'b0010101010: data <= 12'h001; 
        10'b0010101011: data <= 12'hfff; 
        10'b0010101100: data <= 12'hffe; 
        10'b0010101101: data <= 12'h001; 
        10'b0010101110: data <= 12'h007; 
        10'b0010101111: data <= 12'h00d; 
        10'b0010110000: data <= 12'h00a; 
        10'b0010110001: data <= 12'h00b; 
        10'b0010110010: data <= 12'h00f; 
        10'b0010110011: data <= 12'h00a; 
        10'b0010110100: data <= 12'h00a; 
        10'b0010110101: data <= 12'h00d; 
        10'b0010110110: data <= 12'h00c; 
        10'b0010110111: data <= 12'h006; 
        10'b0010111000: data <= 12'h007; 
        10'b0010111001: data <= 12'h002; 
        10'b0010111010: data <= 12'h001; 
        10'b0010111011: data <= 12'hffc; 
        10'b0010111100: data <= 12'hffd; 
        10'b0010111101: data <= 12'hff7; 
        10'b0010111110: data <= 12'hff7; 
        10'b0010111111: data <= 12'hff4; 
        10'b0011000000: data <= 12'hff9; 
        10'b0011000001: data <= 12'hffc; 
        10'b0011000010: data <= 12'h001; 
        10'b0011000011: data <= 12'h000; 
        10'b0011000100: data <= 12'hffe; 
        10'b0011000101: data <= 12'h000; 
        10'b0011000110: data <= 12'h000; 
        10'b0011000111: data <= 12'hffe; 
        10'b0011001000: data <= 12'h000; 
        10'b0011001001: data <= 12'h004; 
        10'b0011001010: data <= 12'h009; 
        10'b0011001011: data <= 12'h00d; 
        10'b0011001100: data <= 12'h00a; 
        10'b0011001101: data <= 12'h00a; 
        10'b0011001110: data <= 12'h004; 
        10'b0011001111: data <= 12'h004; 
        10'b0011010000: data <= 12'h001; 
        10'b0011010001: data <= 12'h007; 
        10'b0011010010: data <= 12'h008; 
        10'b0011010011: data <= 12'h002; 
        10'b0011010100: data <= 12'h001; 
        10'b0011010101: data <= 12'hff5; 
        10'b0011010110: data <= 12'hffc; 
        10'b0011010111: data <= 12'hffd; 
        10'b0011011000: data <= 12'hffd; 
        10'b0011011001: data <= 12'hffc; 
        10'b0011011010: data <= 12'hffd; 
        10'b0011011011: data <= 12'hff6; 
        10'b0011011100: data <= 12'hff9; 
        10'b0011011101: data <= 12'hffe; 
        10'b0011011110: data <= 12'hffd; 
        10'b0011011111: data <= 12'hffd; 
        10'b0011100000: data <= 12'hfff; 
        10'b0011100001: data <= 12'h000; 
        10'b0011100010: data <= 12'hfff; 
        10'b0011100011: data <= 12'h000; 
        10'b0011100100: data <= 12'h002; 
        10'b0011100101: data <= 12'h006; 
        10'b0011100110: data <= 12'h004; 
        10'b0011100111: data <= 12'h006; 
        10'b0011101000: data <= 12'h006; 
        10'b0011101001: data <= 12'h007; 
        10'b0011101010: data <= 12'h007; 
        10'b0011101011: data <= 12'h008; 
        10'b0011101100: data <= 12'h005; 
        10'b0011101101: data <= 12'h006; 
        10'b0011101110: data <= 12'h00f; 
        10'b0011101111: data <= 12'h008; 
        10'b0011110000: data <= 12'hfff; 
        10'b0011110001: data <= 12'hffc; 
        10'b0011110010: data <= 12'h000; 
        10'b0011110011: data <= 12'h003; 
        10'b0011110100: data <= 12'h000; 
        10'b0011110101: data <= 12'hffe; 
        10'b0011110110: data <= 12'hffa; 
        10'b0011110111: data <= 12'hff4; 
        10'b0011111000: data <= 12'hff7; 
        10'b0011111001: data <= 12'hffc; 
        10'b0011111010: data <= 12'hffe; 
        10'b0011111011: data <= 12'hffd; 
        10'b0011111100: data <= 12'hffd; 
        10'b0011111101: data <= 12'hfff; 
        10'b0011111110: data <= 12'h000; 
        10'b0011111111: data <= 12'h002; 
        10'b0100000000: data <= 12'h003; 
        10'b0100000001: data <= 12'h007; 
        10'b0100000010: data <= 12'h002; 
        10'b0100000011: data <= 12'h000; 
        10'b0100000100: data <= 12'hffe; 
        10'b0100000101: data <= 12'h004; 
        10'b0100000110: data <= 12'h003; 
        10'b0100000111: data <= 12'h004; 
        10'b0100001000: data <= 12'h001; 
        10'b0100001001: data <= 12'h000; 
        10'b0100001010: data <= 12'h009; 
        10'b0100001011: data <= 12'h00a; 
        10'b0100001100: data <= 12'h004; 
        10'b0100001101: data <= 12'h000; 
        10'b0100001110: data <= 12'hfff; 
        10'b0100001111: data <= 12'h000; 
        10'b0100010000: data <= 12'h000; 
        10'b0100010001: data <= 12'h000; 
        10'b0100010010: data <= 12'hffc; 
        10'b0100010011: data <= 12'hff6; 
        10'b0100010100: data <= 12'hff7; 
        10'b0100010101: data <= 12'hffd; 
        10'b0100010110: data <= 12'h000; 
        10'b0100010111: data <= 12'hffd; 
        10'b0100011000: data <= 12'h001; 
        10'b0100011001: data <= 12'hfff; 
        10'b0100011010: data <= 12'hfff; 
        10'b0100011011: data <= 12'hffe; 
        10'b0100011100: data <= 12'h000; 
        10'b0100011101: data <= 12'hffe; 
        10'b0100011110: data <= 12'hffd; 
        10'b0100011111: data <= 12'hff0; 
        10'b0100100000: data <= 12'hff2; 
        10'b0100100001: data <= 12'hff5; 
        10'b0100100010: data <= 12'hfef; 
        10'b0100100011: data <= 12'hfee; 
        10'b0100100100: data <= 12'hfeb; 
        10'b0100100101: data <= 12'hfe8; 
        10'b0100100110: data <= 12'hff6; 
        10'b0100100111: data <= 12'h002; 
        10'b0100101000: data <= 12'h003; 
        10'b0100101001: data <= 12'h000; 
        10'b0100101010: data <= 12'h001; 
        10'b0100101011: data <= 12'hffe; 
        10'b0100101100: data <= 12'hfff; 
        10'b0100101101: data <= 12'hffe; 
        10'b0100101110: data <= 12'hffb; 
        10'b0100101111: data <= 12'hff4; 
        10'b0100110000: data <= 12'hffa; 
        10'b0100110001: data <= 12'h000; 
        10'b0100110010: data <= 12'h000; 
        10'b0100110011: data <= 12'hffd; 
        10'b0100110100: data <= 12'hffd; 
        10'b0100110101: data <= 12'h001; 
        10'b0100110110: data <= 12'h000; 
        10'b0100110111: data <= 12'hffd; 
        10'b0100111000: data <= 12'hffa; 
        10'b0100111001: data <= 12'hff3; 
        10'b0100111010: data <= 12'hfea; 
        10'b0100111011: data <= 12'hfe0; 
        10'b0100111100: data <= 12'hfe2; 
        10'b0100111101: data <= 12'hfdc; 
        10'b0100111110: data <= 12'hfdc; 
        10'b0100111111: data <= 12'hfdf; 
        10'b0101000000: data <= 12'hfdd; 
        10'b0101000001: data <= 12'hfd6; 
        10'b0101000010: data <= 12'hfdf; 
        10'b0101000011: data <= 12'hff0; 
        10'b0101000100: data <= 12'hffb; 
        10'b0101000101: data <= 12'hffb; 
        10'b0101000110: data <= 12'hffc; 
        10'b0101000111: data <= 12'hfff; 
        10'b0101001000: data <= 12'hffd; 
        10'b0101001001: data <= 12'hffd; 
        10'b0101001010: data <= 12'hff9; 
        10'b0101001011: data <= 12'hffb; 
        10'b0101001100: data <= 12'hfff; 
        10'b0101001101: data <= 12'hffe; 
        10'b0101001110: data <= 12'hffd; 
        10'b0101001111: data <= 12'hfff; 
        10'b0101010000: data <= 12'hfff; 
        10'b0101010001: data <= 12'hfff; 
        10'b0101010010: data <= 12'h000; 
        10'b0101010011: data <= 12'hfff; 
        10'b0101010100: data <= 12'hffa; 
        10'b0101010101: data <= 12'hfed; 
        10'b0101010110: data <= 12'hfda; 
        10'b0101010111: data <= 12'hfd2; 
        10'b0101011000: data <= 12'hfd5; 
        10'b0101011001: data <= 12'hfd7; 
        10'b0101011010: data <= 12'hfdb; 
        10'b0101011011: data <= 12'hfdd; 
        10'b0101011100: data <= 12'hfdd; 
        10'b0101011101: data <= 12'hfdc; 
        10'b0101011110: data <= 12'hfe2; 
        10'b0101011111: data <= 12'hfec; 
        10'b0101100000: data <= 12'hff2; 
        10'b0101100001: data <= 12'hff4; 
        10'b0101100010: data <= 12'hffa; 
        10'b0101100011: data <= 12'h000; 
        10'b0101100100: data <= 12'h000; 
        10'b0101100101: data <= 12'hffd; 
        10'b0101100110: data <= 12'hff8; 
        10'b0101100111: data <= 12'hff4; 
        10'b0101101000: data <= 12'hfff; 
        10'b0101101001: data <= 12'hffe; 
        10'b0101101010: data <= 12'h001; 
        10'b0101101011: data <= 12'hfff; 
        10'b0101101100: data <= 12'hffe; 
        10'b0101101101: data <= 12'hffe; 
        10'b0101101110: data <= 12'h001; 
        10'b0101101111: data <= 12'hffe; 
        10'b0101110000: data <= 12'hff6; 
        10'b0101110001: data <= 12'hfe7; 
        10'b0101110010: data <= 12'hfd9; 
        10'b0101110011: data <= 12'hfdc; 
        10'b0101110100: data <= 12'hfdf; 
        10'b0101110101: data <= 12'hfe9; 
        10'b0101110110: data <= 12'hff0; 
        10'b0101110111: data <= 12'hff8; 
        10'b0101111000: data <= 12'hff4; 
        10'b0101111001: data <= 12'hffb; 
        10'b0101111010: data <= 12'hff2; 
        10'b0101111011: data <= 12'hff2; 
        10'b0101111100: data <= 12'hfef; 
        10'b0101111101: data <= 12'hff4; 
        10'b0101111110: data <= 12'hff9; 
        10'b0101111111: data <= 12'hfff; 
        10'b0110000000: data <= 12'hffe; 
        10'b0110000001: data <= 12'hffc; 
        10'b0110000010: data <= 12'hff6; 
        10'b0110000011: data <= 12'hff7; 
        10'b0110000100: data <= 12'hffb; 
        10'b0110000101: data <= 12'h001; 
        10'b0110000110: data <= 12'hffe; 
        10'b0110000111: data <= 12'h000; 
        10'b0110001000: data <= 12'h001; 
        10'b0110001001: data <= 12'hfff; 
        10'b0110001010: data <= 12'h000; 
        10'b0110001011: data <= 12'hffe; 
        10'b0110001100: data <= 12'hffc; 
        10'b0110001101: data <= 12'hfef; 
        10'b0110001110: data <= 12'hfeb; 
        10'b0110001111: data <= 12'hfef; 
        10'b0110010000: data <= 12'hff9; 
        10'b0110010001: data <= 12'hfff; 
        10'b0110010010: data <= 12'h004; 
        10'b0110010011: data <= 12'h006; 
        10'b0110010100: data <= 12'h007; 
        10'b0110010101: data <= 12'h00a; 
        10'b0110010110: data <= 12'h001; 
        10'b0110010111: data <= 12'hff9; 
        10'b0110011000: data <= 12'hffb; 
        10'b0110011001: data <= 12'hff7; 
        10'b0110011010: data <= 12'hfff; 
        10'b0110011011: data <= 12'hffa; 
        10'b0110011100: data <= 12'hffe; 
        10'b0110011101: data <= 12'hffa; 
        10'b0110011110: data <= 12'hff5; 
        10'b0110011111: data <= 12'hff8; 
        10'b0110100000: data <= 12'hffe; 
        10'b0110100001: data <= 12'h004; 
        10'b0110100010: data <= 12'h005; 
        10'b0110100011: data <= 12'hffd; 
        10'b0110100100: data <= 12'hffe; 
        10'b0110100101: data <= 12'hfff; 
        10'b0110100110: data <= 12'hffe; 
        10'b0110100111: data <= 12'h004; 
        10'b0110101000: data <= 12'h002; 
        10'b0110101001: data <= 12'h001; 
        10'b0110101010: data <= 12'h004; 
        10'b0110101011: data <= 12'h005; 
        10'b0110101100: data <= 12'h00a; 
        10'b0110101101: data <= 12'h007; 
        10'b0110101110: data <= 12'h008; 
        10'b0110101111: data <= 12'h005; 
        10'b0110110000: data <= 12'h004; 
        10'b0110110001: data <= 12'h00a; 
        10'b0110110010: data <= 12'h001; 
        10'b0110110011: data <= 12'h004; 
        10'b0110110100: data <= 12'h001; 
        10'b0110110101: data <= 12'hff8; 
        10'b0110110110: data <= 12'hff8; 
        10'b0110110111: data <= 12'hffb; 
        10'b0110111000: data <= 12'hffd; 
        10'b0110111001: data <= 12'hffb; 
        10'b0110111010: data <= 12'hff6; 
        10'b0110111011: data <= 12'hffb; 
        10'b0110111100: data <= 12'h003; 
        10'b0110111101: data <= 12'h005; 
        10'b0110111110: data <= 12'h003; 
        10'b0110111111: data <= 12'hffd; 
        10'b0111000000: data <= 12'hffe; 
        10'b0111000001: data <= 12'hffd; 
        10'b0111000010: data <= 12'hffc; 
        10'b0111000011: data <= 12'h004; 
        10'b0111000100: data <= 12'h008; 
        10'b0111000101: data <= 12'h00e; 
        10'b0111000110: data <= 12'h00e; 
        10'b0111000111: data <= 12'h008; 
        10'b0111001000: data <= 12'h003; 
        10'b0111001001: data <= 12'h007; 
        10'b0111001010: data <= 12'h007; 
        10'b0111001011: data <= 12'h006; 
        10'b0111001100: data <= 12'h00d; 
        10'b0111001101: data <= 12'h00b; 
        10'b0111001110: data <= 12'h002; 
        10'b0111001111: data <= 12'hfff; 
        10'b0111010000: data <= 12'h000; 
        10'b0111010001: data <= 12'hffb; 
        10'b0111010010: data <= 12'hffb; 
        10'b0111010011: data <= 12'hff8; 
        10'b0111010100: data <= 12'hffd; 
        10'b0111010101: data <= 12'h000; 
        10'b0111010110: data <= 12'h002; 
        10'b0111010111: data <= 12'h004; 
        10'b0111011000: data <= 12'h00c; 
        10'b0111011001: data <= 12'h00f; 
        10'b0111011010: data <= 12'h002; 
        10'b0111011011: data <= 12'hffe; 
        10'b0111011100: data <= 12'hffe; 
        10'b0111011101: data <= 12'h001; 
        10'b0111011110: data <= 12'hfff; 
        10'b0111011111: data <= 12'h005; 
        10'b0111100000: data <= 12'h00e; 
        10'b0111100001: data <= 12'h014; 
        10'b0111100010: data <= 12'h012; 
        10'b0111100011: data <= 12'h00d; 
        10'b0111100100: data <= 12'h009; 
        10'b0111100101: data <= 12'h00b; 
        10'b0111100110: data <= 12'h010; 
        10'b0111100111: data <= 12'h00d; 
        10'b0111101000: data <= 12'h00f; 
        10'b0111101001: data <= 12'h007; 
        10'b0111101010: data <= 12'h004; 
        10'b0111101011: data <= 12'h005; 
        10'b0111101100: data <= 12'h005; 
        10'b0111101101: data <= 12'hfff; 
        10'b0111101110: data <= 12'h003; 
        10'b0111101111: data <= 12'hffe; 
        10'b0111110000: data <= 12'h006; 
        10'b0111110001: data <= 12'h006; 
        10'b0111110010: data <= 12'h005; 
        10'b0111110011: data <= 12'h007; 
        10'b0111110100: data <= 12'h013; 
        10'b0111110101: data <= 12'h010; 
        10'b0111110110: data <= 12'h004; 
        10'b0111110111: data <= 12'h000; 
        10'b0111111000: data <= 12'h000; 
        10'b0111111001: data <= 12'h000; 
        10'b0111111010: data <= 12'hffb; 
        10'b0111111011: data <= 12'h001; 
        10'b0111111100: data <= 12'h010; 
        10'b0111111101: data <= 12'h01a; 
        10'b0111111110: data <= 12'h019; 
        10'b0111111111: data <= 12'h012; 
        10'b1000000000: data <= 12'h00c; 
        10'b1000000001: data <= 12'h00d; 
        10'b1000000010: data <= 12'h014; 
        10'b1000000011: data <= 12'h012; 
        10'b1000000100: data <= 12'h01d; 
        10'b1000000101: data <= 12'h015; 
        10'b1000000110: data <= 12'h013; 
        10'b1000000111: data <= 12'h009; 
        10'b1000001000: data <= 12'h006; 
        10'b1000001001: data <= 12'h00b; 
        10'b1000001010: data <= 12'h007; 
        10'b1000001011: data <= 12'h005; 
        10'b1000001100: data <= 12'h00e; 
        10'b1000001101: data <= 12'h00e; 
        10'b1000001110: data <= 12'h00f; 
        10'b1000001111: data <= 12'h014; 
        10'b1000010000: data <= 12'h019; 
        10'b1000010001: data <= 12'h00e; 
        10'b1000010010: data <= 12'hfff; 
        10'b1000010011: data <= 12'hffd; 
        10'b1000010100: data <= 12'hffd; 
        10'b1000010101: data <= 12'hffe; 
        10'b1000010110: data <= 12'hffd; 
        10'b1000010111: data <= 12'h000; 
        10'b1000011000: data <= 12'h009; 
        10'b1000011001: data <= 12'h010; 
        10'b1000011010: data <= 12'h014; 
        10'b1000011011: data <= 12'h012; 
        10'b1000011100: data <= 12'h010; 
        10'b1000011101: data <= 12'h011; 
        10'b1000011110: data <= 12'h010; 
        10'b1000011111: data <= 12'h012; 
        10'b1000100000: data <= 12'h014; 
        10'b1000100001: data <= 12'h00f; 
        10'b1000100010: data <= 12'h00a; 
        10'b1000100011: data <= 12'h005; 
        10'b1000100100: data <= 12'h007; 
        10'b1000100101: data <= 12'h00c; 
        10'b1000100110: data <= 12'h006; 
        10'b1000100111: data <= 12'h006; 
        10'b1000101000: data <= 12'h00a; 
        10'b1000101001: data <= 12'h00d; 
        10'b1000101010: data <= 12'h010; 
        10'b1000101011: data <= 12'h012; 
        10'b1000101100: data <= 12'h00f; 
        10'b1000101101: data <= 12'h008; 
        10'b1000101110: data <= 12'h001; 
        10'b1000101111: data <= 12'h000; 
        10'b1000110000: data <= 12'hffd; 
        10'b1000110001: data <= 12'h000; 
        10'b1000110010: data <= 12'hfff; 
        10'b1000110011: data <= 12'hffc; 
        10'b1000110100: data <= 12'h008; 
        10'b1000110101: data <= 12'h009; 
        10'b1000110110: data <= 12'h00f; 
        10'b1000110111: data <= 12'h014; 
        10'b1000111000: data <= 12'h013; 
        10'b1000111001: data <= 12'h00d; 
        10'b1000111010: data <= 12'h00c; 
        10'b1000111011: data <= 12'h015; 
        10'b1000111100: data <= 12'h00b; 
        10'b1000111101: data <= 12'h004; 
        10'b1000111110: data <= 12'h003; 
        10'b1000111111: data <= 12'h003; 
        10'b1001000000: data <= 12'h004; 
        10'b1001000001: data <= 12'h000; 
        10'b1001000010: data <= 12'h009; 
        10'b1001000011: data <= 12'h00e; 
        10'b1001000100: data <= 12'h009; 
        10'b1001000101: data <= 12'h00d; 
        10'b1001000110: data <= 12'h013; 
        10'b1001000111: data <= 12'h010; 
        10'b1001001000: data <= 12'h00c; 
        10'b1001001001: data <= 12'h006; 
        10'b1001001010: data <= 12'h000; 
        10'b1001001011: data <= 12'hfff; 
        10'b1001001100: data <= 12'hfff; 
        10'b1001001101: data <= 12'hffd; 
        10'b1001001110: data <= 12'hfff; 
        10'b1001001111: data <= 12'hffe; 
        10'b1001010000: data <= 12'h002; 
        10'b1001010001: data <= 12'h004; 
        10'b1001010010: data <= 12'h00a; 
        10'b1001010011: data <= 12'h00b; 
        10'b1001010100: data <= 12'h00a; 
        10'b1001010101: data <= 12'h00d; 
        10'b1001010110: data <= 12'h00b; 
        10'b1001010111: data <= 12'h00b; 
        10'b1001011000: data <= 12'h004; 
        10'b1001011001: data <= 12'h002; 
        10'b1001011010: data <= 12'hfff; 
        10'b1001011011: data <= 12'h000; 
        10'b1001011100: data <= 12'h005; 
        10'b1001011101: data <= 12'h006; 
        10'b1001011110: data <= 12'h00d; 
        10'b1001011111: data <= 12'h00e; 
        10'b1001100000: data <= 12'h006; 
        10'b1001100001: data <= 12'h00d; 
        10'b1001100010: data <= 12'h011; 
        10'b1001100011: data <= 12'h013; 
        10'b1001100100: data <= 12'h009; 
        10'b1001100101: data <= 12'h004; 
        10'b1001100110: data <= 12'h001; 
        10'b1001100111: data <= 12'h000; 
        10'b1001101000: data <= 12'hffd; 
        10'b1001101001: data <= 12'hfff; 
        10'b1001101010: data <= 12'hffd; 
        10'b1001101011: data <= 12'h001; 
        10'b1001101100: data <= 12'h003; 
        10'b1001101101: data <= 12'h001; 
        10'b1001101110: data <= 12'h007; 
        10'b1001101111: data <= 12'h006; 
        10'b1001110000: data <= 12'h006; 
        10'b1001110001: data <= 12'h008; 
        10'b1001110010: data <= 12'h008; 
        10'b1001110011: data <= 12'h009; 
        10'b1001110100: data <= 12'h001; 
        10'b1001110101: data <= 12'hff9; 
        10'b1001110110: data <= 12'hff7; 
        10'b1001110111: data <= 12'hffb; 
        10'b1001111000: data <= 12'hffb; 
        10'b1001111001: data <= 12'h004; 
        10'b1001111010: data <= 12'h00c; 
        10'b1001111011: data <= 12'h00f; 
        10'b1001111100: data <= 12'h00e; 
        10'b1001111101: data <= 12'h00d; 
        10'b1001111110: data <= 12'h00c; 
        10'b1001111111: data <= 12'h00d; 
        10'b1010000000: data <= 12'h005; 
        10'b1010000001: data <= 12'hfff; 
        10'b1010000010: data <= 12'hfff; 
        10'b1010000011: data <= 12'hffe; 
        10'b1010000100: data <= 12'hfff; 
        10'b1010000101: data <= 12'hfff; 
        10'b1010000110: data <= 12'hfff; 
        10'b1010000111: data <= 12'hffe; 
        10'b1010001000: data <= 12'hffe; 
        10'b1010001001: data <= 12'hffc; 
        10'b1010001010: data <= 12'hffc; 
        10'b1010001011: data <= 12'hffc; 
        10'b1010001100: data <= 12'hffa; 
        10'b1010001101: data <= 12'hffc; 
        10'b1010001110: data <= 12'hffe; 
        10'b1010001111: data <= 12'h003; 
        10'b1010010000: data <= 12'h000; 
        10'b1010010001: data <= 12'hffb; 
        10'b1010010010: data <= 12'hff9; 
        10'b1010010011: data <= 12'hff7; 
        10'b1010010100: data <= 12'hff7; 
        10'b1010010101: data <= 12'hffb; 
        10'b1010010110: data <= 12'h002; 
        10'b1010010111: data <= 12'h00c; 
        10'b1010011000: data <= 12'h00b; 
        10'b1010011001: data <= 12'h00d; 
        10'b1010011010: data <= 12'h009; 
        10'b1010011011: data <= 12'h004; 
        10'b1010011100: data <= 12'h002; 
        10'b1010011101: data <= 12'h001; 
        10'b1010011110: data <= 12'h000; 
        10'b1010011111: data <= 12'hffe; 
        10'b1010100000: data <= 12'hfff; 
        10'b1010100001: data <= 12'hffe; 
        10'b1010100010: data <= 12'h000; 
        10'b1010100011: data <= 12'h000; 
        10'b1010100100: data <= 12'hffd; 
        10'b1010100101: data <= 12'hff9; 
        10'b1010100110: data <= 12'hff3; 
        10'b1010100111: data <= 12'hff6; 
        10'b1010101000: data <= 12'hff6; 
        10'b1010101001: data <= 12'hff5; 
        10'b1010101010: data <= 12'hff5; 
        10'b1010101011: data <= 12'hff8; 
        10'b1010101100: data <= 12'hff8; 
        10'b1010101101: data <= 12'hffc; 
        10'b1010101110: data <= 12'hffa; 
        10'b1010101111: data <= 12'hff8; 
        10'b1010110000: data <= 12'hff8; 
        10'b1010110001: data <= 12'hffa; 
        10'b1010110010: data <= 12'hff8; 
        10'b1010110011: data <= 12'hffc; 
        10'b1010110100: data <= 12'hffc; 
        10'b1010110101: data <= 12'hffc; 
        10'b1010110110: data <= 12'hffe; 
        10'b1010110111: data <= 12'hffe; 
        10'b1010111000: data <= 12'h000; 
        10'b1010111001: data <= 12'h001; 
        10'b1010111010: data <= 12'hffd; 
        10'b1010111011: data <= 12'hffd; 
        10'b1010111100: data <= 12'h000; 
        10'b1010111101: data <= 12'hffc; 
        10'b1010111110: data <= 12'hffe; 
        10'b1010111111: data <= 12'hffe; 
        10'b1011000000: data <= 12'hffd; 
        10'b1011000001: data <= 12'hffb; 
        10'b1011000010: data <= 12'hffa; 
        10'b1011000011: data <= 12'hff6; 
        10'b1011000100: data <= 12'hff5; 
        10'b1011000101: data <= 12'hff6; 
        10'b1011000110: data <= 12'hff7; 
        10'b1011000111: data <= 12'hff5; 
        10'b1011001000: data <= 12'hff8; 
        10'b1011001001: data <= 12'hff9; 
        10'b1011001010: data <= 12'hff6; 
        10'b1011001011: data <= 12'hff8; 
        10'b1011001100: data <= 12'hffa; 
        10'b1011001101: data <= 12'hffb; 
        10'b1011001110: data <= 12'hffe; 
        10'b1011001111: data <= 12'hffb; 
        10'b1011010000: data <= 12'hffe; 
        10'b1011010001: data <= 12'hffe; 
        10'b1011010010: data <= 12'h000; 
        10'b1011010011: data <= 12'hffd; 
        10'b1011010100: data <= 12'hfff; 
        10'b1011010101: data <= 12'hffd; 
        10'b1011010110: data <= 12'hffd; 
        10'b1011010111: data <= 12'hffd; 
        10'b1011011000: data <= 12'hffd; 
        10'b1011011001: data <= 12'hffe; 
        10'b1011011010: data <= 12'hffe; 
        10'b1011011011: data <= 12'h000; 
        10'b1011011100: data <= 12'hfff; 
        10'b1011011101: data <= 12'hffe; 
        10'b1011011110: data <= 12'hfff; 
        10'b1011011111: data <= 12'h000; 
        10'b1011100000: data <= 12'hffe; 
        10'b1011100001: data <= 12'h000; 
        10'b1011100010: data <= 12'h000; 
        10'b1011100011: data <= 12'h000; 
        10'b1011100100: data <= 12'h000; 
        10'b1011100101: data <= 12'hfff; 
        10'b1011100110: data <= 12'hffe; 
        10'b1011100111: data <= 12'hffc; 
        10'b1011101000: data <= 12'hffe; 
        10'b1011101001: data <= 12'hfff; 
        10'b1011101010: data <= 12'hfff; 
        10'b1011101011: data <= 12'hffd; 
        10'b1011101100: data <= 12'h000; 
        10'b1011101101: data <= 12'h000; 
        10'b1011101110: data <= 12'hffd; 
        10'b1011101111: data <= 12'hffe; 
        10'b1011110000: data <= 12'hffd; 
        10'b1011110001: data <= 12'h000; 
        10'b1011110010: data <= 12'h000; 
        10'b1011110011: data <= 12'h000; 
        10'b1011110100: data <= 12'h000; 
        10'b1011110101: data <= 12'hffe; 
        10'b1011110110: data <= 12'hffd; 
        10'b1011110111: data <= 12'hfff; 
        10'b1011111000: data <= 12'hffd; 
        10'b1011111001: data <= 12'h001; 
        10'b1011111010: data <= 12'h001; 
        10'b1011111011: data <= 12'hffe; 
        10'b1011111100: data <= 12'h000; 
        10'b1011111101: data <= 12'hffd; 
        10'b1011111110: data <= 12'h000; 
        10'b1011111111: data <= 12'hffd; 
        10'b1100000000: data <= 12'h000; 
        10'b1100000001: data <= 12'hffe; 
        10'b1100000010: data <= 12'hfff; 
        10'b1100000011: data <= 12'hffd; 
        10'b1100000100: data <= 12'hfff; 
        10'b1100000101: data <= 12'hffe; 
        10'b1100000110: data <= 12'hfff; 
        10'b1100000111: data <= 12'hfff; 
        10'b1100001000: data <= 12'h000; 
        10'b1100001001: data <= 12'hffc; 
        10'b1100001010: data <= 12'hffe; 
        10'b1100001011: data <= 12'h000; 
        10'b1100001100: data <= 12'hffc; 
        10'b1100001101: data <= 12'hfff; 
        10'b1100001110: data <= 12'hfff; 
        10'b1100001111: data <= 12'hffe; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 7) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 13'h1ffa; 
        10'b0000000001: data <= 13'h0000; 
        10'b0000000010: data <= 13'h1ffd; 
        10'b0000000011: data <= 13'h1ffb; 
        10'b0000000100: data <= 13'h1ffd; 
        10'b0000000101: data <= 13'h1ffb; 
        10'b0000000110: data <= 13'h1ffe; 
        10'b0000000111: data <= 13'h1ffe; 
        10'b0000001000: data <= 13'h1ff9; 
        10'b0000001001: data <= 13'h1ffd; 
        10'b0000001010: data <= 13'h1ffa; 
        10'b0000001011: data <= 13'h1ffc; 
        10'b0000001100: data <= 13'h0001; 
        10'b0000001101: data <= 13'h0001; 
        10'b0000001110: data <= 13'h1ffa; 
        10'b0000001111: data <= 13'h1ffe; 
        10'b0000010000: data <= 13'h1ffa; 
        10'b0000010001: data <= 13'h1ffa; 
        10'b0000010010: data <= 13'h0002; 
        10'b0000010011: data <= 13'h0000; 
        10'b0000010100: data <= 13'h1ffb; 
        10'b0000010101: data <= 13'h1ffe; 
        10'b0000010110: data <= 13'h1ffc; 
        10'b0000010111: data <= 13'h1ff9; 
        10'b0000011000: data <= 13'h1ffa; 
        10'b0000011001: data <= 13'h1ffe; 
        10'b0000011010: data <= 13'h0000; 
        10'b0000011011: data <= 13'h1ffe; 
        10'b0000011100: data <= 13'h1ffd; 
        10'b0000011101: data <= 13'h1ffd; 
        10'b0000011110: data <= 13'h0002; 
        10'b0000011111: data <= 13'h1ffe; 
        10'b0000100000: data <= 13'h1ffa; 
        10'b0000100001: data <= 13'h1ffa; 
        10'b0000100010: data <= 13'h1ff9; 
        10'b0000100011: data <= 13'h1ffb; 
        10'b0000100100: data <= 13'h1ffb; 
        10'b0000100101: data <= 13'h1ffe; 
        10'b0000100110: data <= 13'h0000; 
        10'b0000100111: data <= 13'h1ffa; 
        10'b0000101000: data <= 13'h1ffc; 
        10'b0000101001: data <= 13'h1ffa; 
        10'b0000101010: data <= 13'h1ffe; 
        10'b0000101011: data <= 13'h1ff9; 
        10'b0000101100: data <= 13'h1ffe; 
        10'b0000101101: data <= 13'h1ffa; 
        10'b0000101110: data <= 13'h1ffc; 
        10'b0000101111: data <= 13'h1ffb; 
        10'b0000110000: data <= 13'h1ffe; 
        10'b0000110001: data <= 13'h1ffa; 
        10'b0000110010: data <= 13'h1ff9; 
        10'b0000110011: data <= 13'h1ff9; 
        10'b0000110100: data <= 13'h0000; 
        10'b0000110101: data <= 13'h1ffe; 
        10'b0000110110: data <= 13'h0000; 
        10'b0000110111: data <= 13'h1ffc; 
        10'b0000111000: data <= 13'h1ffd; 
        10'b0000111001: data <= 13'h1ff9; 
        10'b0000111010: data <= 13'h1ffa; 
        10'b0000111011: data <= 13'h0000; 
        10'b0000111100: data <= 13'h1ff9; 
        10'b0000111101: data <= 13'h1ffa; 
        10'b0000111110: data <= 13'h1ffd; 
        10'b0000111111: data <= 13'h1ffe; 
        10'b0001000000: data <= 13'h1fff; 
        10'b0001000001: data <= 13'h1ffc; 
        10'b0001000010: data <= 13'h0004; 
        10'b0001000011: data <= 13'h0003; 
        10'b0001000100: data <= 13'h0009; 
        10'b0001000101: data <= 13'h0007; 
        10'b0001000110: data <= 13'h0007; 
        10'b0001000111: data <= 13'h0003; 
        10'b0001001000: data <= 13'h0009; 
        10'b0001001001: data <= 13'h0003; 
        10'b0001001010: data <= 13'h0003; 
        10'b0001001011: data <= 13'h1ffb; 
        10'b0001001100: data <= 13'h0000; 
        10'b0001001101: data <= 13'h1ffe; 
        10'b0001001110: data <= 13'h1ff7; 
        10'b0001001111: data <= 13'h1ffd; 
        10'b0001010000: data <= 13'h1fff; 
        10'b0001010001: data <= 13'h0002; 
        10'b0001010010: data <= 13'h1ffd; 
        10'b0001010011: data <= 13'h1ffc; 
        10'b0001010100: data <= 13'h1ffb; 
        10'b0001010101: data <= 13'h1ffb; 
        10'b0001010110: data <= 13'h1fff; 
        10'b0001010111: data <= 13'h1ffb; 
        10'b0001011000: data <= 13'h0001; 
        10'b0001011001: data <= 13'h1ffa; 
        10'b0001011010: data <= 13'h1ffe; 
        10'b0001011011: data <= 13'h0000; 
        10'b0001011100: data <= 13'h0002; 
        10'b0001011101: data <= 13'h000f; 
        10'b0001011110: data <= 13'h0017; 
        10'b0001011111: data <= 13'h0017; 
        10'b0001100000: data <= 13'h0016; 
        10'b0001100001: data <= 13'h0020; 
        10'b0001100010: data <= 13'h0012; 
        10'b0001100011: data <= 13'h0008; 
        10'b0001100100: data <= 13'h000f; 
        10'b0001100101: data <= 13'h0007; 
        10'b0001100110: data <= 13'h1ffa; 
        10'b0001100111: data <= 13'h1ffe; 
        10'b0001101000: data <= 13'h1ff9; 
        10'b0001101001: data <= 13'h1ff7; 
        10'b0001101010: data <= 13'h1ff6; 
        10'b0001101011: data <= 13'h1ffb; 
        10'b0001101100: data <= 13'h0001; 
        10'b0001101101: data <= 13'h0002; 
        10'b0001101110: data <= 13'h1ffa; 
        10'b0001101111: data <= 13'h1fff; 
        10'b0001110000: data <= 13'h1ffb; 
        10'b0001110001: data <= 13'h1ffc; 
        10'b0001110010: data <= 13'h0002; 
        10'b0001110011: data <= 13'h1ff8; 
        10'b0001110100: data <= 13'h1ff9; 
        10'b0001110101: data <= 13'h1ffe; 
        10'b0001110110: data <= 13'h0003; 
        10'b0001110111: data <= 13'h0003; 
        10'b0001111000: data <= 13'h0009; 
        10'b0001111001: data <= 13'h001c; 
        10'b0001111010: data <= 13'h001c; 
        10'b0001111011: data <= 13'h0024; 
        10'b0001111100: data <= 13'h001e; 
        10'b0001111101: data <= 13'h0018; 
        10'b0001111110: data <= 13'h0016; 
        10'b0001111111: data <= 13'h000a; 
        10'b0010000000: data <= 13'h000d; 
        10'b0010000001: data <= 13'h000c; 
        10'b0010000010: data <= 13'h1ffc; 
        10'b0010000011: data <= 13'h1ffa; 
        10'b0010000100: data <= 13'h1ffb; 
        10'b0010000101: data <= 13'h1ff2; 
        10'b0010000110: data <= 13'h1fef; 
        10'b0010000111: data <= 13'h1ff0; 
        10'b0010001000: data <= 13'h1ffe; 
        10'b0010001001: data <= 13'h1ffe; 
        10'b0010001010: data <= 13'h1ff9; 
        10'b0010001011: data <= 13'h1fff; 
        10'b0010001100: data <= 13'h0001; 
        10'b0010001101: data <= 13'h1ffe; 
        10'b0010001110: data <= 13'h1ffb; 
        10'b0010001111: data <= 13'h1ff9; 
        10'b0010010000: data <= 13'h1ffa; 
        10'b0010010001: data <= 13'h1ffb; 
        10'b0010010010: data <= 13'h0003; 
        10'b0010010011: data <= 13'h000e; 
        10'b0010010100: data <= 13'h0013; 
        10'b0010010101: data <= 13'h0021; 
        10'b0010010110: data <= 13'h0024; 
        10'b0010010111: data <= 13'h0026; 
        10'b0010011000: data <= 13'h0023; 
        10'b0010011001: data <= 13'h0027; 
        10'b0010011010: data <= 13'h0024; 
        10'b0010011011: data <= 13'h0021; 
        10'b0010011100: data <= 13'h0024; 
        10'b0010011101: data <= 13'h001d; 
        10'b0010011110: data <= 13'h0015; 
        10'b0010011111: data <= 13'h1ff7; 
        10'b0010100000: data <= 13'h1ff7; 
        10'b0010100001: data <= 13'h1ff2; 
        10'b0010100010: data <= 13'h1ff2; 
        10'b0010100011: data <= 13'h1fea; 
        10'b0010100100: data <= 13'h1ff6; 
        10'b0010100101: data <= 13'h1ffb; 
        10'b0010100110: data <= 13'h0001; 
        10'b0010100111: data <= 13'h1ffc; 
        10'b0010101000: data <= 13'h1ffd; 
        10'b0010101001: data <= 13'h1ffb; 
        10'b0010101010: data <= 13'h0001; 
        10'b0010101011: data <= 13'h1ffd; 
        10'b0010101100: data <= 13'h1ffc; 
        10'b0010101101: data <= 13'h0002; 
        10'b0010101110: data <= 13'h000d; 
        10'b0010101111: data <= 13'h001a; 
        10'b0010110000: data <= 13'h0014; 
        10'b0010110001: data <= 13'h0017; 
        10'b0010110010: data <= 13'h001f; 
        10'b0010110011: data <= 13'h0013; 
        10'b0010110100: data <= 13'h0014; 
        10'b0010110101: data <= 13'h001a; 
        10'b0010110110: data <= 13'h0017; 
        10'b0010110111: data <= 13'h000d; 
        10'b0010111000: data <= 13'h000e; 
        10'b0010111001: data <= 13'h0004; 
        10'b0010111010: data <= 13'h0003; 
        10'b0010111011: data <= 13'h1ff8; 
        10'b0010111100: data <= 13'h1ffb; 
        10'b0010111101: data <= 13'h1fee; 
        10'b0010111110: data <= 13'h1fee; 
        10'b0010111111: data <= 13'h1fe7; 
        10'b0011000000: data <= 13'h1ff1; 
        10'b0011000001: data <= 13'h1ff8; 
        10'b0011000010: data <= 13'h0001; 
        10'b0011000011: data <= 13'h1fff; 
        10'b0011000100: data <= 13'h1ffc; 
        10'b0011000101: data <= 13'h0001; 
        10'b0011000110: data <= 13'h0001; 
        10'b0011000111: data <= 13'h1ffd; 
        10'b0011001000: data <= 13'h0000; 
        10'b0011001001: data <= 13'h0007; 
        10'b0011001010: data <= 13'h0011; 
        10'b0011001011: data <= 13'h0019; 
        10'b0011001100: data <= 13'h0015; 
        10'b0011001101: data <= 13'h0013; 
        10'b0011001110: data <= 13'h0007; 
        10'b0011001111: data <= 13'h0009; 
        10'b0011010000: data <= 13'h0001; 
        10'b0011010001: data <= 13'h000d; 
        10'b0011010010: data <= 13'h0011; 
        10'b0011010011: data <= 13'h0003; 
        10'b0011010100: data <= 13'h0002; 
        10'b0011010101: data <= 13'h1feb; 
        10'b0011010110: data <= 13'h1ff9; 
        10'b0011010111: data <= 13'h1ffa; 
        10'b0011011000: data <= 13'h1ff9; 
        10'b0011011001: data <= 13'h1ff8; 
        10'b0011011010: data <= 13'h1ffa; 
        10'b0011011011: data <= 13'h1fec; 
        10'b0011011100: data <= 13'h1ff2; 
        10'b0011011101: data <= 13'h1ffc; 
        10'b0011011110: data <= 13'h1ffb; 
        10'b0011011111: data <= 13'h1ff9; 
        10'b0011100000: data <= 13'h1ffe; 
        10'b0011100001: data <= 13'h0001; 
        10'b0011100010: data <= 13'h1ffd; 
        10'b0011100011: data <= 13'h0001; 
        10'b0011100100: data <= 13'h0004; 
        10'b0011100101: data <= 13'h000c; 
        10'b0011100110: data <= 13'h0009; 
        10'b0011100111: data <= 13'h000c; 
        10'b0011101000: data <= 13'h000c; 
        10'b0011101001: data <= 13'h000e; 
        10'b0011101010: data <= 13'h000e; 
        10'b0011101011: data <= 13'h0010; 
        10'b0011101100: data <= 13'h0009; 
        10'b0011101101: data <= 13'h000b; 
        10'b0011101110: data <= 13'h001d; 
        10'b0011101111: data <= 13'h0010; 
        10'b0011110000: data <= 13'h1ffe; 
        10'b0011110001: data <= 13'h1ff8; 
        10'b0011110010: data <= 13'h0000; 
        10'b0011110011: data <= 13'h0006; 
        10'b0011110100: data <= 13'h0000; 
        10'b0011110101: data <= 13'h1ffc; 
        10'b0011110110: data <= 13'h1ff4; 
        10'b0011110111: data <= 13'h1fe8; 
        10'b0011111000: data <= 13'h1fee; 
        10'b0011111001: data <= 13'h1ff8; 
        10'b0011111010: data <= 13'h1ffc; 
        10'b0011111011: data <= 13'h1ffa; 
        10'b0011111100: data <= 13'h1ffb; 
        10'b0011111101: data <= 13'h1fff; 
        10'b0011111110: data <= 13'h0000; 
        10'b0011111111: data <= 13'h0003; 
        10'b0100000000: data <= 13'h0006; 
        10'b0100000001: data <= 13'h000d; 
        10'b0100000010: data <= 13'h0005; 
        10'b0100000011: data <= 13'h0001; 
        10'b0100000100: data <= 13'h1ffb; 
        10'b0100000101: data <= 13'h0007; 
        10'b0100000110: data <= 13'h0006; 
        10'b0100000111: data <= 13'h0007; 
        10'b0100001000: data <= 13'h0002; 
        10'b0100001001: data <= 13'h1fff; 
        10'b0100001010: data <= 13'h0013; 
        10'b0100001011: data <= 13'h0015; 
        10'b0100001100: data <= 13'h0007; 
        10'b0100001101: data <= 13'h0001; 
        10'b0100001110: data <= 13'h1ffe; 
        10'b0100001111: data <= 13'h0000; 
        10'b0100010000: data <= 13'h1fff; 
        10'b0100010001: data <= 13'h0000; 
        10'b0100010010: data <= 13'h1ff8; 
        10'b0100010011: data <= 13'h1fec; 
        10'b0100010100: data <= 13'h1fef; 
        10'b0100010101: data <= 13'h1ffa; 
        10'b0100010110: data <= 13'h0001; 
        10'b0100010111: data <= 13'h1ff9; 
        10'b0100011000: data <= 13'h0001; 
        10'b0100011001: data <= 13'h1fff; 
        10'b0100011010: data <= 13'h1ffd; 
        10'b0100011011: data <= 13'h1ffc; 
        10'b0100011100: data <= 13'h0001; 
        10'b0100011101: data <= 13'h1ffd; 
        10'b0100011110: data <= 13'h1ff9; 
        10'b0100011111: data <= 13'h1fe0; 
        10'b0100100000: data <= 13'h1fe3; 
        10'b0100100001: data <= 13'h1fea; 
        10'b0100100010: data <= 13'h1fdf; 
        10'b0100100011: data <= 13'h1fdb; 
        10'b0100100100: data <= 13'h1fd5; 
        10'b0100100101: data <= 13'h1fd0; 
        10'b0100100110: data <= 13'h1fec; 
        10'b0100100111: data <= 13'h0004; 
        10'b0100101000: data <= 13'h0005; 
        10'b0100101001: data <= 13'h0001; 
        10'b0100101010: data <= 13'h0003; 
        10'b0100101011: data <= 13'h1ffc; 
        10'b0100101100: data <= 13'h1ffd; 
        10'b0100101101: data <= 13'h1ffc; 
        10'b0100101110: data <= 13'h1ff6; 
        10'b0100101111: data <= 13'h1fe9; 
        10'b0100110000: data <= 13'h1ff3; 
        10'b0100110001: data <= 13'h1fff; 
        10'b0100110010: data <= 13'h1fff; 
        10'b0100110011: data <= 13'h1ffb; 
        10'b0100110100: data <= 13'h1ff9; 
        10'b0100110101: data <= 13'h0002; 
        10'b0100110110: data <= 13'h1fff; 
        10'b0100110111: data <= 13'h1ffa; 
        10'b0100111000: data <= 13'h1ff4; 
        10'b0100111001: data <= 13'h1fe6; 
        10'b0100111010: data <= 13'h1fd3; 
        10'b0100111011: data <= 13'h1fc1; 
        10'b0100111100: data <= 13'h1fc3; 
        10'b0100111101: data <= 13'h1fb8; 
        10'b0100111110: data <= 13'h1fb8; 
        10'b0100111111: data <= 13'h1fbe; 
        10'b0101000000: data <= 13'h1fba; 
        10'b0101000001: data <= 13'h1fab; 
        10'b0101000010: data <= 13'h1fbf; 
        10'b0101000011: data <= 13'h1fe1; 
        10'b0101000100: data <= 13'h1ff5; 
        10'b0101000101: data <= 13'h1ff7; 
        10'b0101000110: data <= 13'h1ff7; 
        10'b0101000111: data <= 13'h1ffe; 
        10'b0101001000: data <= 13'h1ffb; 
        10'b0101001001: data <= 13'h1ffa; 
        10'b0101001010: data <= 13'h1ff1; 
        10'b0101001011: data <= 13'h1ff6; 
        10'b0101001100: data <= 13'h1ffe; 
        10'b0101001101: data <= 13'h1ffc; 
        10'b0101001110: data <= 13'h1ffa; 
        10'b0101001111: data <= 13'h1ffe; 
        10'b0101010000: data <= 13'h1ffe; 
        10'b0101010001: data <= 13'h1ffe; 
        10'b0101010010: data <= 13'h0001; 
        10'b0101010011: data <= 13'h1ffd; 
        10'b0101010100: data <= 13'h1ff3; 
        10'b0101010101: data <= 13'h1fd9; 
        10'b0101010110: data <= 13'h1fb4; 
        10'b0101010111: data <= 13'h1fa3; 
        10'b0101011000: data <= 13'h1fa9; 
        10'b0101011001: data <= 13'h1fae; 
        10'b0101011010: data <= 13'h1fb5; 
        10'b0101011011: data <= 13'h1fba; 
        10'b0101011100: data <= 13'h1fba; 
        10'b0101011101: data <= 13'h1fb7; 
        10'b0101011110: data <= 13'h1fc4; 
        10'b0101011111: data <= 13'h1fd8; 
        10'b0101100000: data <= 13'h1fe5; 
        10'b0101100001: data <= 13'h1fe7; 
        10'b0101100010: data <= 13'h1ff4; 
        10'b0101100011: data <= 13'h0000; 
        10'b0101100100: data <= 13'h0000; 
        10'b0101100101: data <= 13'h1ff9; 
        10'b0101100110: data <= 13'h1ff0; 
        10'b0101100111: data <= 13'h1fe8; 
        10'b0101101000: data <= 13'h1ffd; 
        10'b0101101001: data <= 13'h1ffc; 
        10'b0101101010: data <= 13'h0002; 
        10'b0101101011: data <= 13'h1ffe; 
        10'b0101101100: data <= 13'h1ffb; 
        10'b0101101101: data <= 13'h1ffd; 
        10'b0101101110: data <= 13'h0002; 
        10'b0101101111: data <= 13'h1ffb; 
        10'b0101110000: data <= 13'h1feb; 
        10'b0101110001: data <= 13'h1fcf; 
        10'b0101110010: data <= 13'h1fb2; 
        10'b0101110011: data <= 13'h1fb8; 
        10'b0101110100: data <= 13'h1fbd; 
        10'b0101110101: data <= 13'h1fd2; 
        10'b0101110110: data <= 13'h1fdf; 
        10'b0101110111: data <= 13'h1ff1; 
        10'b0101111000: data <= 13'h1fe8; 
        10'b0101111001: data <= 13'h1ff5; 
        10'b0101111010: data <= 13'h1fe4; 
        10'b0101111011: data <= 13'h1fe4; 
        10'b0101111100: data <= 13'h1fdf; 
        10'b0101111101: data <= 13'h1fe8; 
        10'b0101111110: data <= 13'h1ff3; 
        10'b0101111111: data <= 13'h1ffd; 
        10'b0110000000: data <= 13'h1ffc; 
        10'b0110000001: data <= 13'h1ff7; 
        10'b0110000010: data <= 13'h1fec; 
        10'b0110000011: data <= 13'h1fee; 
        10'b0110000100: data <= 13'h1ff7; 
        10'b0110000101: data <= 13'h0002; 
        10'b0110000110: data <= 13'h1ffd; 
        10'b0110000111: data <= 13'h0000; 
        10'b0110001000: data <= 13'h0001; 
        10'b0110001001: data <= 13'h1ffe; 
        10'b0110001010: data <= 13'h0000; 
        10'b0110001011: data <= 13'h1ffc; 
        10'b0110001100: data <= 13'h1ff8; 
        10'b0110001101: data <= 13'h1fdf; 
        10'b0110001110: data <= 13'h1fd6; 
        10'b0110001111: data <= 13'h1fde; 
        10'b0110010000: data <= 13'h1ff2; 
        10'b0110010001: data <= 13'h1ffe; 
        10'b0110010010: data <= 13'h0009; 
        10'b0110010011: data <= 13'h000b; 
        10'b0110010100: data <= 13'h000d; 
        10'b0110010101: data <= 13'h0015; 
        10'b0110010110: data <= 13'h0001; 
        10'b0110010111: data <= 13'h1ff3; 
        10'b0110011000: data <= 13'h1ff6; 
        10'b0110011001: data <= 13'h1fef; 
        10'b0110011010: data <= 13'h1ffd; 
        10'b0110011011: data <= 13'h1ff5; 
        10'b0110011100: data <= 13'h1ffc; 
        10'b0110011101: data <= 13'h1ff3; 
        10'b0110011110: data <= 13'h1fe9; 
        10'b0110011111: data <= 13'h1fef; 
        10'b0110100000: data <= 13'h1ffd; 
        10'b0110100001: data <= 13'h0008; 
        10'b0110100010: data <= 13'h0009; 
        10'b0110100011: data <= 13'h1ffb; 
        10'b0110100100: data <= 13'h1ffc; 
        10'b0110100101: data <= 13'h1ffd; 
        10'b0110100110: data <= 13'h1ffc; 
        10'b0110100111: data <= 13'h0008; 
        10'b0110101000: data <= 13'h0004; 
        10'b0110101001: data <= 13'h0002; 
        10'b0110101010: data <= 13'h0009; 
        10'b0110101011: data <= 13'h000b; 
        10'b0110101100: data <= 13'h0014; 
        10'b0110101101: data <= 13'h000e; 
        10'b0110101110: data <= 13'h0011; 
        10'b0110101111: data <= 13'h000a; 
        10'b0110110000: data <= 13'h0009; 
        10'b0110110001: data <= 13'h0014; 
        10'b0110110010: data <= 13'h0002; 
        10'b0110110011: data <= 13'h0008; 
        10'b0110110100: data <= 13'h0001; 
        10'b0110110101: data <= 13'h1ff0; 
        10'b0110110110: data <= 13'h1ff1; 
        10'b0110110111: data <= 13'h1ff7; 
        10'b0110111000: data <= 13'h1ff9; 
        10'b0110111001: data <= 13'h1ff6; 
        10'b0110111010: data <= 13'h1feb; 
        10'b0110111011: data <= 13'h1ff5; 
        10'b0110111100: data <= 13'h0006; 
        10'b0110111101: data <= 13'h000b; 
        10'b0110111110: data <= 13'h0006; 
        10'b0110111111: data <= 13'h1ffa; 
        10'b0111000000: data <= 13'h1ffc; 
        10'b0111000001: data <= 13'h1ff9; 
        10'b0111000010: data <= 13'h1ff8; 
        10'b0111000011: data <= 13'h0008; 
        10'b0111000100: data <= 13'h0011; 
        10'b0111000101: data <= 13'h001c; 
        10'b0111000110: data <= 13'h001c; 
        10'b0111000111: data <= 13'h0011; 
        10'b0111001000: data <= 13'h0007; 
        10'b0111001001: data <= 13'h000e; 
        10'b0111001010: data <= 13'h000d; 
        10'b0111001011: data <= 13'h000c; 
        10'b0111001100: data <= 13'h0019; 
        10'b0111001101: data <= 13'h0016; 
        10'b0111001110: data <= 13'h0005; 
        10'b0111001111: data <= 13'h1ffd; 
        10'b0111010000: data <= 13'h0000; 
        10'b0111010001: data <= 13'h1ff6; 
        10'b0111010010: data <= 13'h1ff7; 
        10'b0111010011: data <= 13'h1ff0; 
        10'b0111010100: data <= 13'h1ffa; 
        10'b0111010101: data <= 13'h0001; 
        10'b0111010110: data <= 13'h0004; 
        10'b0111010111: data <= 13'h0007; 
        10'b0111011000: data <= 13'h0018; 
        10'b0111011001: data <= 13'h001d; 
        10'b0111011010: data <= 13'h0005; 
        10'b0111011011: data <= 13'h1ffb; 
        10'b0111011100: data <= 13'h1ffc; 
        10'b0111011101: data <= 13'h0001; 
        10'b0111011110: data <= 13'h1ffd; 
        10'b0111011111: data <= 13'h000a; 
        10'b0111100000: data <= 13'h001d; 
        10'b0111100001: data <= 13'h0028; 
        10'b0111100010: data <= 13'h0025; 
        10'b0111100011: data <= 13'h0019; 
        10'b0111100100: data <= 13'h0012; 
        10'b0111100101: data <= 13'h0015; 
        10'b0111100110: data <= 13'h0021; 
        10'b0111100111: data <= 13'h001b; 
        10'b0111101000: data <= 13'h001f; 
        10'b0111101001: data <= 13'h000e; 
        10'b0111101010: data <= 13'h0007; 
        10'b0111101011: data <= 13'h000a; 
        10'b0111101100: data <= 13'h000a; 
        10'b0111101101: data <= 13'h1ffe; 
        10'b0111101110: data <= 13'h0007; 
        10'b0111101111: data <= 13'h1ffc; 
        10'b0111110000: data <= 13'h000c; 
        10'b0111110001: data <= 13'h000d; 
        10'b0111110010: data <= 13'h000a; 
        10'b0111110011: data <= 13'h000d; 
        10'b0111110100: data <= 13'h0026; 
        10'b0111110101: data <= 13'h0021; 
        10'b0111110110: data <= 13'h0007; 
        10'b0111110111: data <= 13'h0001; 
        10'b0111111000: data <= 13'h1fff; 
        10'b0111111001: data <= 13'h0000; 
        10'b0111111010: data <= 13'h1ff6; 
        10'b0111111011: data <= 13'h0003; 
        10'b0111111100: data <= 13'h001f; 
        10'b0111111101: data <= 13'h0035; 
        10'b0111111110: data <= 13'h0032; 
        10'b0111111111: data <= 13'h0024; 
        10'b1000000000: data <= 13'h0018; 
        10'b1000000001: data <= 13'h001b; 
        10'b1000000010: data <= 13'h0029; 
        10'b1000000011: data <= 13'h0025; 
        10'b1000000100: data <= 13'h003b; 
        10'b1000000101: data <= 13'h002b; 
        10'b1000000110: data <= 13'h0025; 
        10'b1000000111: data <= 13'h0012; 
        10'b1000001000: data <= 13'h000c; 
        10'b1000001001: data <= 13'h0017; 
        10'b1000001010: data <= 13'h000f; 
        10'b1000001011: data <= 13'h000a; 
        10'b1000001100: data <= 13'h001b; 
        10'b1000001101: data <= 13'h001c; 
        10'b1000001110: data <= 13'h001e; 
        10'b1000001111: data <= 13'h0028; 
        10'b1000010000: data <= 13'h0032; 
        10'b1000010001: data <= 13'h001d; 
        10'b1000010010: data <= 13'h1ffd; 
        10'b1000010011: data <= 13'h1ffa; 
        10'b1000010100: data <= 13'h1ffb; 
        10'b1000010101: data <= 13'h1ffb; 
        10'b1000010110: data <= 13'h1ff9; 
        10'b1000010111: data <= 13'h0000; 
        10'b1000011000: data <= 13'h0011; 
        10'b1000011001: data <= 13'h0020; 
        10'b1000011010: data <= 13'h0029; 
        10'b1000011011: data <= 13'h0023; 
        10'b1000011100: data <= 13'h0021; 
        10'b1000011101: data <= 13'h0022; 
        10'b1000011110: data <= 13'h0021; 
        10'b1000011111: data <= 13'h0023; 
        10'b1000100000: data <= 13'h0027; 
        10'b1000100001: data <= 13'h001e; 
        10'b1000100010: data <= 13'h0014; 
        10'b1000100011: data <= 13'h0009; 
        10'b1000100100: data <= 13'h000e; 
        10'b1000100101: data <= 13'h0019; 
        10'b1000100110: data <= 13'h000c; 
        10'b1000100111: data <= 13'h000c; 
        10'b1000101000: data <= 13'h0014; 
        10'b1000101001: data <= 13'h0019; 
        10'b1000101010: data <= 13'h0021; 
        10'b1000101011: data <= 13'h0023; 
        10'b1000101100: data <= 13'h001e; 
        10'b1000101101: data <= 13'h0010; 
        10'b1000101110: data <= 13'h0001; 
        10'b1000101111: data <= 13'h0000; 
        10'b1000110000: data <= 13'h1ffa; 
        10'b1000110001: data <= 13'h0000; 
        10'b1000110010: data <= 13'h1ffe; 
        10'b1000110011: data <= 13'h1ff7; 
        10'b1000110100: data <= 13'h000f; 
        10'b1000110101: data <= 13'h0013; 
        10'b1000110110: data <= 13'h001d; 
        10'b1000110111: data <= 13'h0029; 
        10'b1000111000: data <= 13'h0027; 
        10'b1000111001: data <= 13'h001a; 
        10'b1000111010: data <= 13'h0019; 
        10'b1000111011: data <= 13'h0029; 
        10'b1000111100: data <= 13'h0017; 
        10'b1000111101: data <= 13'h0008; 
        10'b1000111110: data <= 13'h0005; 
        10'b1000111111: data <= 13'h0006; 
        10'b1001000000: data <= 13'h0008; 
        10'b1001000001: data <= 13'h0000; 
        10'b1001000010: data <= 13'h0012; 
        10'b1001000011: data <= 13'h001c; 
        10'b1001000100: data <= 13'h0013; 
        10'b1001000101: data <= 13'h001b; 
        10'b1001000110: data <= 13'h0025; 
        10'b1001000111: data <= 13'h0021; 
        10'b1001001000: data <= 13'h0017; 
        10'b1001001001: data <= 13'h000b; 
        10'b1001001010: data <= 13'h0000; 
        10'b1001001011: data <= 13'h1fff; 
        10'b1001001100: data <= 13'h1ffe; 
        10'b1001001101: data <= 13'h1ffa; 
        10'b1001001110: data <= 13'h1fff; 
        10'b1001001111: data <= 13'h1ffd; 
        10'b1001010000: data <= 13'h0003; 
        10'b1001010001: data <= 13'h0008; 
        10'b1001010010: data <= 13'h0014; 
        10'b1001010011: data <= 13'h0017; 
        10'b1001010100: data <= 13'h0014; 
        10'b1001010101: data <= 13'h0019; 
        10'b1001010110: data <= 13'h0016; 
        10'b1001010111: data <= 13'h0016; 
        10'b1001011000: data <= 13'h0009; 
        10'b1001011001: data <= 13'h0004; 
        10'b1001011010: data <= 13'h1ffe; 
        10'b1001011011: data <= 13'h0001; 
        10'b1001011100: data <= 13'h000b; 
        10'b1001011101: data <= 13'h000c; 
        10'b1001011110: data <= 13'h001a; 
        10'b1001011111: data <= 13'h001b; 
        10'b1001100000: data <= 13'h000c; 
        10'b1001100001: data <= 13'h001b; 
        10'b1001100010: data <= 13'h0021; 
        10'b1001100011: data <= 13'h0026; 
        10'b1001100100: data <= 13'h0013; 
        10'b1001100101: data <= 13'h0007; 
        10'b1001100110: data <= 13'h0002; 
        10'b1001100111: data <= 13'h1fff; 
        10'b1001101000: data <= 13'h1ffa; 
        10'b1001101001: data <= 13'h1ffe; 
        10'b1001101010: data <= 13'h1ffb; 
        10'b1001101011: data <= 13'h0002; 
        10'b1001101100: data <= 13'h0006; 
        10'b1001101101: data <= 13'h0002; 
        10'b1001101110: data <= 13'h000e; 
        10'b1001101111: data <= 13'h000c; 
        10'b1001110000: data <= 13'h000b; 
        10'b1001110001: data <= 13'h0010; 
        10'b1001110010: data <= 13'h0010; 
        10'b1001110011: data <= 13'h0013; 
        10'b1001110100: data <= 13'h0002; 
        10'b1001110101: data <= 13'h1ff1; 
        10'b1001110110: data <= 13'h1fed; 
        10'b1001110111: data <= 13'h1ff5; 
        10'b1001111000: data <= 13'h1ff6; 
        10'b1001111001: data <= 13'h0008; 
        10'b1001111010: data <= 13'h0018; 
        10'b1001111011: data <= 13'h001f; 
        10'b1001111100: data <= 13'h001c; 
        10'b1001111101: data <= 13'h001b; 
        10'b1001111110: data <= 13'h0017; 
        10'b1001111111: data <= 13'h001a; 
        10'b1010000000: data <= 13'h000a; 
        10'b1010000001: data <= 13'h1fff; 
        10'b1010000010: data <= 13'h1ffe; 
        10'b1010000011: data <= 13'h1ffc; 
        10'b1010000100: data <= 13'h1ffe; 
        10'b1010000101: data <= 13'h1fff; 
        10'b1010000110: data <= 13'h1ffd; 
        10'b1010000111: data <= 13'h1ffd; 
        10'b1010001000: data <= 13'h1ffc; 
        10'b1010001001: data <= 13'h1ff9; 
        10'b1010001010: data <= 13'h1ff7; 
        10'b1010001011: data <= 13'h1ff8; 
        10'b1010001100: data <= 13'h1ff3; 
        10'b1010001101: data <= 13'h1ff9; 
        10'b1010001110: data <= 13'h1ffb; 
        10'b1010001111: data <= 13'h0006; 
        10'b1010010000: data <= 13'h0001; 
        10'b1010010001: data <= 13'h1ff6; 
        10'b1010010010: data <= 13'h1ff3; 
        10'b1010010011: data <= 13'h1fee; 
        10'b1010010100: data <= 13'h1fed; 
        10'b1010010101: data <= 13'h1ff6; 
        10'b1010010110: data <= 13'h0004; 
        10'b1010010111: data <= 13'h0018; 
        10'b1010011000: data <= 13'h0015; 
        10'b1010011001: data <= 13'h001a; 
        10'b1010011010: data <= 13'h0013; 
        10'b1010011011: data <= 13'h0007; 
        10'b1010011100: data <= 13'h0004; 
        10'b1010011101: data <= 13'h0003; 
        10'b1010011110: data <= 13'h1fff; 
        10'b1010011111: data <= 13'h1ffd; 
        10'b1010100000: data <= 13'h1ffe; 
        10'b1010100001: data <= 13'h1ffb; 
        10'b1010100010: data <= 13'h0000; 
        10'b1010100011: data <= 13'h1fff; 
        10'b1010100100: data <= 13'h1ffb; 
        10'b1010100101: data <= 13'h1ff2; 
        10'b1010100110: data <= 13'h1fe6; 
        10'b1010100111: data <= 13'h1fec; 
        10'b1010101000: data <= 13'h1fec; 
        10'b1010101001: data <= 13'h1fea; 
        10'b1010101010: data <= 13'h1feb; 
        10'b1010101011: data <= 13'h1ff0; 
        10'b1010101100: data <= 13'h1ff0; 
        10'b1010101101: data <= 13'h1ff7; 
        10'b1010101110: data <= 13'h1ff4; 
        10'b1010101111: data <= 13'h1fef; 
        10'b1010110000: data <= 13'h1ff0; 
        10'b1010110001: data <= 13'h1ff4; 
        10'b1010110010: data <= 13'h1ff1; 
        10'b1010110011: data <= 13'h1ff8; 
        10'b1010110100: data <= 13'h1ff9; 
        10'b1010110101: data <= 13'h1ff9; 
        10'b1010110110: data <= 13'h1ffc; 
        10'b1010110111: data <= 13'h1ffd; 
        10'b1010111000: data <= 13'h0000; 
        10'b1010111001: data <= 13'h0003; 
        10'b1010111010: data <= 13'h1ffa; 
        10'b1010111011: data <= 13'h1ffb; 
        10'b1010111100: data <= 13'h0000; 
        10'b1010111101: data <= 13'h1ff9; 
        10'b1010111110: data <= 13'h1ffc; 
        10'b1010111111: data <= 13'h1ffc; 
        10'b1011000000: data <= 13'h1ffa; 
        10'b1011000001: data <= 13'h1ff6; 
        10'b1011000010: data <= 13'h1ff3; 
        10'b1011000011: data <= 13'h1fed; 
        10'b1011000100: data <= 13'h1feb; 
        10'b1011000101: data <= 13'h1fec; 
        10'b1011000110: data <= 13'h1fee; 
        10'b1011000111: data <= 13'h1fe9; 
        10'b1011001000: data <= 13'h1ff1; 
        10'b1011001001: data <= 13'h1ff2; 
        10'b1011001010: data <= 13'h1fed; 
        10'b1011001011: data <= 13'h1ff0; 
        10'b1011001100: data <= 13'h1ff4; 
        10'b1011001101: data <= 13'h1ff5; 
        10'b1011001110: data <= 13'h1ffc; 
        10'b1011001111: data <= 13'h1ff6; 
        10'b1011010000: data <= 13'h1ffc; 
        10'b1011010001: data <= 13'h1ffc; 
        10'b1011010010: data <= 13'h0000; 
        10'b1011010011: data <= 13'h1ffb; 
        10'b1011010100: data <= 13'h1ffe; 
        10'b1011010101: data <= 13'h1ffb; 
        10'b1011010110: data <= 13'h1ff9; 
        10'b1011010111: data <= 13'h1ffb; 
        10'b1011011000: data <= 13'h1ff9; 
        10'b1011011001: data <= 13'h1ffc; 
        10'b1011011010: data <= 13'h1ffd; 
        10'b1011011011: data <= 13'h0000; 
        10'b1011011100: data <= 13'h1fff; 
        10'b1011011101: data <= 13'h1ffd; 
        10'b1011011110: data <= 13'h1fff; 
        10'b1011011111: data <= 13'h0000; 
        10'b1011100000: data <= 13'h1ffd; 
        10'b1011100001: data <= 13'h0000; 
        10'b1011100010: data <= 13'h0000; 
        10'b1011100011: data <= 13'h0000; 
        10'b1011100100: data <= 13'h0001; 
        10'b1011100101: data <= 13'h1ffe; 
        10'b1011100110: data <= 13'h1ffb; 
        10'b1011100111: data <= 13'h1ff8; 
        10'b1011101000: data <= 13'h1ffc; 
        10'b1011101001: data <= 13'h1ffe; 
        10'b1011101010: data <= 13'h1ffd; 
        10'b1011101011: data <= 13'h1ffb; 
        10'b1011101100: data <= 13'h0001; 
        10'b1011101101: data <= 13'h0000; 
        10'b1011101110: data <= 13'h1ffb; 
        10'b1011101111: data <= 13'h1ffc; 
        10'b1011110000: data <= 13'h1ff9; 
        10'b1011110001: data <= 13'h0000; 
        10'b1011110010: data <= 13'h0000; 
        10'b1011110011: data <= 13'h0000; 
        10'b1011110100: data <= 13'h1fff; 
        10'b1011110101: data <= 13'h1ffb; 
        10'b1011110110: data <= 13'h1ffa; 
        10'b1011110111: data <= 13'h1ffe; 
        10'b1011111000: data <= 13'h1ff9; 
        10'b1011111001: data <= 13'h0001; 
        10'b1011111010: data <= 13'h0001; 
        10'b1011111011: data <= 13'h1ffc; 
        10'b1011111100: data <= 13'h0000; 
        10'b1011111101: data <= 13'h1ffb; 
        10'b1011111110: data <= 13'h0001; 
        10'b1011111111: data <= 13'h1ff9; 
        10'b1100000000: data <= 13'h0000; 
        10'b1100000001: data <= 13'h1ffd; 
        10'b1100000010: data <= 13'h1ffe; 
        10'b1100000011: data <= 13'h1ffa; 
        10'b1100000100: data <= 13'h1ffe; 
        10'b1100000101: data <= 13'h1ffc; 
        10'b1100000110: data <= 13'h1ffe; 
        10'b1100000111: data <= 13'h1ffd; 
        10'b1100001000: data <= 13'h1fff; 
        10'b1100001001: data <= 13'h1ff9; 
        10'b1100001010: data <= 13'h1ffd; 
        10'b1100001011: data <= 13'h0000; 
        10'b1100001100: data <= 13'h1ff9; 
        10'b1100001101: data <= 13'h1ffd; 
        10'b1100001110: data <= 13'h1fff; 
        10'b1100001111: data <= 13'h1ffc; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 8) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 14'h3ff3; 
        10'b0000000001: data <= 14'h0000; 
        10'b0000000010: data <= 14'h3ffa; 
        10'b0000000011: data <= 14'h3ff5; 
        10'b0000000100: data <= 14'h3ff9; 
        10'b0000000101: data <= 14'h3ff6; 
        10'b0000000110: data <= 14'h3ffc; 
        10'b0000000111: data <= 14'h3ffc; 
        10'b0000001000: data <= 14'h3ff3; 
        10'b0000001001: data <= 14'h3ffb; 
        10'b0000001010: data <= 14'h3ff4; 
        10'b0000001011: data <= 14'h3ff8; 
        10'b0000001100: data <= 14'h0002; 
        10'b0000001101: data <= 14'h0002; 
        10'b0000001110: data <= 14'h3ff3; 
        10'b0000001111: data <= 14'h3ffb; 
        10'b0000010000: data <= 14'h3ff4; 
        10'b0000010001: data <= 14'h3ff5; 
        10'b0000010010: data <= 14'h0003; 
        10'b0000010011: data <= 14'h0001; 
        10'b0000010100: data <= 14'h3ff6; 
        10'b0000010101: data <= 14'h3ffc; 
        10'b0000010110: data <= 14'h3ff8; 
        10'b0000010111: data <= 14'h3ff2; 
        10'b0000011000: data <= 14'h3ff3; 
        10'b0000011001: data <= 14'h3ffb; 
        10'b0000011010: data <= 14'h3fff; 
        10'b0000011011: data <= 14'h3ffc; 
        10'b0000011100: data <= 14'h3ffb; 
        10'b0000011101: data <= 14'h3ffa; 
        10'b0000011110: data <= 14'h0003; 
        10'b0000011111: data <= 14'h3ffd; 
        10'b0000100000: data <= 14'h3ff4; 
        10'b0000100001: data <= 14'h3ff3; 
        10'b0000100010: data <= 14'h3ff3; 
        10'b0000100011: data <= 14'h3ff6; 
        10'b0000100100: data <= 14'h3ff6; 
        10'b0000100101: data <= 14'h3ffb; 
        10'b0000100110: data <= 14'h0000; 
        10'b0000100111: data <= 14'h3ff4; 
        10'b0000101000: data <= 14'h3ff8; 
        10'b0000101001: data <= 14'h3ff4; 
        10'b0000101010: data <= 14'h3ffc; 
        10'b0000101011: data <= 14'h3ff2; 
        10'b0000101100: data <= 14'h3ffc; 
        10'b0000101101: data <= 14'h3ff4; 
        10'b0000101110: data <= 14'h3ff8; 
        10'b0000101111: data <= 14'h3ff5; 
        10'b0000110000: data <= 14'h3ffc; 
        10'b0000110001: data <= 14'h3ff5; 
        10'b0000110010: data <= 14'h3ff3; 
        10'b0000110011: data <= 14'h3ff1; 
        10'b0000110100: data <= 14'h0001; 
        10'b0000110101: data <= 14'h3ffd; 
        10'b0000110110: data <= 14'h0001; 
        10'b0000110111: data <= 14'h3ff7; 
        10'b0000111000: data <= 14'h3ffa; 
        10'b0000111001: data <= 14'h3ff2; 
        10'b0000111010: data <= 14'h3ff4; 
        10'b0000111011: data <= 14'h0000; 
        10'b0000111100: data <= 14'h3ff3; 
        10'b0000111101: data <= 14'h3ff4; 
        10'b0000111110: data <= 14'h3ff9; 
        10'b0000111111: data <= 14'h3ffb; 
        10'b0001000000: data <= 14'h3fff; 
        10'b0001000001: data <= 14'h3ff8; 
        10'b0001000010: data <= 14'h0007; 
        10'b0001000011: data <= 14'h0006; 
        10'b0001000100: data <= 14'h0012; 
        10'b0001000101: data <= 14'h000f; 
        10'b0001000110: data <= 14'h000d; 
        10'b0001000111: data <= 14'h0005; 
        10'b0001001000: data <= 14'h0012; 
        10'b0001001001: data <= 14'h0006; 
        10'b0001001010: data <= 14'h0005; 
        10'b0001001011: data <= 14'h3ff7; 
        10'b0001001100: data <= 14'h0000; 
        10'b0001001101: data <= 14'h3ffc; 
        10'b0001001110: data <= 14'h3fed; 
        10'b0001001111: data <= 14'h3ff9; 
        10'b0001010000: data <= 14'h3ffe; 
        10'b0001010001: data <= 14'h0005; 
        10'b0001010010: data <= 14'h3ffb; 
        10'b0001010011: data <= 14'h3ff8; 
        10'b0001010100: data <= 14'h3ff7; 
        10'b0001010101: data <= 14'h3ff6; 
        10'b0001010110: data <= 14'h3ffd; 
        10'b0001010111: data <= 14'h3ff6; 
        10'b0001011000: data <= 14'h0003; 
        10'b0001011001: data <= 14'h3ff4; 
        10'b0001011010: data <= 14'h3ffc; 
        10'b0001011011: data <= 14'h0000; 
        10'b0001011100: data <= 14'h0003; 
        10'b0001011101: data <= 14'h001d; 
        10'b0001011110: data <= 14'h002e; 
        10'b0001011111: data <= 14'h002e; 
        10'b0001100000: data <= 14'h002c; 
        10'b0001100001: data <= 14'h0040; 
        10'b0001100010: data <= 14'h0023; 
        10'b0001100011: data <= 14'h0010; 
        10'b0001100100: data <= 14'h001e; 
        10'b0001100101: data <= 14'h000e; 
        10'b0001100110: data <= 14'h3ff3; 
        10'b0001100111: data <= 14'h3ffd; 
        10'b0001101000: data <= 14'h3ff1; 
        10'b0001101001: data <= 14'h3fef; 
        10'b0001101010: data <= 14'h3feb; 
        10'b0001101011: data <= 14'h3ff6; 
        10'b0001101100: data <= 14'h0002; 
        10'b0001101101: data <= 14'h0005; 
        10'b0001101110: data <= 14'h3ff4; 
        10'b0001101111: data <= 14'h3ffe; 
        10'b0001110000: data <= 14'h3ff6; 
        10'b0001110001: data <= 14'h3ff9; 
        10'b0001110010: data <= 14'h0004; 
        10'b0001110011: data <= 14'h3ff1; 
        10'b0001110100: data <= 14'h3ff3; 
        10'b0001110101: data <= 14'h3ffc; 
        10'b0001110110: data <= 14'h0007; 
        10'b0001110111: data <= 14'h0007; 
        10'b0001111000: data <= 14'h0013; 
        10'b0001111001: data <= 14'h0038; 
        10'b0001111010: data <= 14'h0039; 
        10'b0001111011: data <= 14'h0048; 
        10'b0001111100: data <= 14'h003d; 
        10'b0001111101: data <= 14'h0030; 
        10'b0001111110: data <= 14'h002c; 
        10'b0001111111: data <= 14'h0013; 
        10'b0010000000: data <= 14'h001a; 
        10'b0010000001: data <= 14'h0018; 
        10'b0010000010: data <= 14'h3ff9; 
        10'b0010000011: data <= 14'h3ff4; 
        10'b0010000100: data <= 14'h3ff7; 
        10'b0010000101: data <= 14'h3fe4; 
        10'b0010000110: data <= 14'h3fde; 
        10'b0010000111: data <= 14'h3fdf; 
        10'b0010001000: data <= 14'h3ffc; 
        10'b0010001001: data <= 14'h3ffc; 
        10'b0010001010: data <= 14'h3ff2; 
        10'b0010001011: data <= 14'h3ffd; 
        10'b0010001100: data <= 14'h0001; 
        10'b0010001101: data <= 14'h3ffc; 
        10'b0010001110: data <= 14'h3ff5; 
        10'b0010001111: data <= 14'h3ff1; 
        10'b0010010000: data <= 14'h3ff4; 
        10'b0010010001: data <= 14'h3ff6; 
        10'b0010010010: data <= 14'h0006; 
        10'b0010010011: data <= 14'h001c; 
        10'b0010010100: data <= 14'h0026; 
        10'b0010010101: data <= 14'h0041; 
        10'b0010010110: data <= 14'h0048; 
        10'b0010010111: data <= 14'h004c; 
        10'b0010011000: data <= 14'h0045; 
        10'b0010011001: data <= 14'h004e; 
        10'b0010011010: data <= 14'h0048; 
        10'b0010011011: data <= 14'h0043; 
        10'b0010011100: data <= 14'h0048; 
        10'b0010011101: data <= 14'h003b; 
        10'b0010011110: data <= 14'h002a; 
        10'b0010011111: data <= 14'h3fee; 
        10'b0010100000: data <= 14'h3fef; 
        10'b0010100001: data <= 14'h3fe4; 
        10'b0010100010: data <= 14'h3fe3; 
        10'b0010100011: data <= 14'h3fd4; 
        10'b0010100100: data <= 14'h3fed; 
        10'b0010100101: data <= 14'h3ff5; 
        10'b0010100110: data <= 14'h0002; 
        10'b0010100111: data <= 14'h3ff8; 
        10'b0010101000: data <= 14'h3ffa; 
        10'b0010101001: data <= 14'h3ff6; 
        10'b0010101010: data <= 14'h0002; 
        10'b0010101011: data <= 14'h3ffa; 
        10'b0010101100: data <= 14'h3ff9; 
        10'b0010101101: data <= 14'h0005; 
        10'b0010101110: data <= 14'h001b; 
        10'b0010101111: data <= 14'h0034; 
        10'b0010110000: data <= 14'h0028; 
        10'b0010110001: data <= 14'h002d; 
        10'b0010110010: data <= 14'h003d; 
        10'b0010110011: data <= 14'h0026; 
        10'b0010110100: data <= 14'h0029; 
        10'b0010110101: data <= 14'h0035; 
        10'b0010110110: data <= 14'h002e; 
        10'b0010110111: data <= 14'h0019; 
        10'b0010111000: data <= 14'h001c; 
        10'b0010111001: data <= 14'h0007; 
        10'b0010111010: data <= 14'h0005; 
        10'b0010111011: data <= 14'h3ff0; 
        10'b0010111100: data <= 14'h3ff5; 
        10'b0010111101: data <= 14'h3fdc; 
        10'b0010111110: data <= 14'h3fdc; 
        10'b0010111111: data <= 14'h3fce; 
        10'b0011000000: data <= 14'h3fe2; 
        10'b0011000001: data <= 14'h3fef; 
        10'b0011000010: data <= 14'h0002; 
        10'b0011000011: data <= 14'h3ffe; 
        10'b0011000100: data <= 14'h3ff8; 
        10'b0011000101: data <= 14'h0002; 
        10'b0011000110: data <= 14'h0002; 
        10'b0011000111: data <= 14'h3ff9; 
        10'b0011001000: data <= 14'h0001; 
        10'b0011001001: data <= 14'h000e; 
        10'b0011001010: data <= 14'h0023; 
        10'b0011001011: data <= 14'h0032; 
        10'b0011001100: data <= 14'h0029; 
        10'b0011001101: data <= 14'h0026; 
        10'b0011001110: data <= 14'h000f; 
        10'b0011001111: data <= 14'h0011; 
        10'b0011010000: data <= 14'h0003; 
        10'b0011010001: data <= 14'h001b; 
        10'b0011010010: data <= 14'h0021; 
        10'b0011010011: data <= 14'h0007; 
        10'b0011010100: data <= 14'h0004; 
        10'b0011010101: data <= 14'h3fd6; 
        10'b0011010110: data <= 14'h3ff2; 
        10'b0011010111: data <= 14'h3ff4; 
        10'b0011011000: data <= 14'h3ff3; 
        10'b0011011001: data <= 14'h3ff0; 
        10'b0011011010: data <= 14'h3ff4; 
        10'b0011011011: data <= 14'h3fd7; 
        10'b0011011100: data <= 14'h3fe4; 
        10'b0011011101: data <= 14'h3ff7; 
        10'b0011011110: data <= 14'h3ff5; 
        10'b0011011111: data <= 14'h3ff3; 
        10'b0011100000: data <= 14'h3ffd; 
        10'b0011100001: data <= 14'h0002; 
        10'b0011100010: data <= 14'h3ffa; 
        10'b0011100011: data <= 14'h0002; 
        10'b0011100100: data <= 14'h0008; 
        10'b0011100101: data <= 14'h0018; 
        10'b0011100110: data <= 14'h0011; 
        10'b0011100111: data <= 14'h0018; 
        10'b0011101000: data <= 14'h0018; 
        10'b0011101001: data <= 14'h001b; 
        10'b0011101010: data <= 14'h001b; 
        10'b0011101011: data <= 14'h001f; 
        10'b0011101100: data <= 14'h0012; 
        10'b0011101101: data <= 14'h0016; 
        10'b0011101110: data <= 14'h003a; 
        10'b0011101111: data <= 14'h0021; 
        10'b0011110000: data <= 14'h3ffc; 
        10'b0011110001: data <= 14'h3ff0; 
        10'b0011110010: data <= 14'h0000; 
        10'b0011110011: data <= 14'h000d; 
        10'b0011110100: data <= 14'h0000; 
        10'b0011110101: data <= 14'h3ff7; 
        10'b0011110110: data <= 14'h3fe8; 
        10'b0011110111: data <= 14'h3fd0; 
        10'b0011111000: data <= 14'h3fdb; 
        10'b0011111001: data <= 14'h3ff1; 
        10'b0011111010: data <= 14'h3ff9; 
        10'b0011111011: data <= 14'h3ff4; 
        10'b0011111100: data <= 14'h3ff6; 
        10'b0011111101: data <= 14'h3ffe; 
        10'b0011111110: data <= 14'h3fff; 
        10'b0011111111: data <= 14'h0006; 
        10'b0100000000: data <= 14'h000c; 
        10'b0100000001: data <= 14'h001a; 
        10'b0100000010: data <= 14'h0009; 
        10'b0100000011: data <= 14'h0002; 
        10'b0100000100: data <= 14'h3ff7; 
        10'b0100000101: data <= 14'h000e; 
        10'b0100000110: data <= 14'h000b; 
        10'b0100000111: data <= 14'h000e; 
        10'b0100001000: data <= 14'h0004; 
        10'b0100001001: data <= 14'h3fff; 
        10'b0100001010: data <= 14'h0026; 
        10'b0100001011: data <= 14'h0029; 
        10'b0100001100: data <= 14'h000e; 
        10'b0100001101: data <= 14'h0001; 
        10'b0100001110: data <= 14'h3ffc; 
        10'b0100001111: data <= 14'h0000; 
        10'b0100010000: data <= 14'h3ffe; 
        10'b0100010001: data <= 14'h3fff; 
        10'b0100010010: data <= 14'h3ff1; 
        10'b0100010011: data <= 14'h3fd7; 
        10'b0100010100: data <= 14'h3fdd; 
        10'b0100010101: data <= 14'h3ff5; 
        10'b0100010110: data <= 14'h0002; 
        10'b0100010111: data <= 14'h3ff3; 
        10'b0100011000: data <= 14'h0003; 
        10'b0100011001: data <= 14'h3ffd; 
        10'b0100011010: data <= 14'h3ffa; 
        10'b0100011011: data <= 14'h3ff7; 
        10'b0100011100: data <= 14'h0002; 
        10'b0100011101: data <= 14'h3ffa; 
        10'b0100011110: data <= 14'h3ff3; 
        10'b0100011111: data <= 14'h3fc0; 
        10'b0100100000: data <= 14'h3fc7; 
        10'b0100100001: data <= 14'h3fd5; 
        10'b0100100010: data <= 14'h3fbe; 
        10'b0100100011: data <= 14'h3fb7; 
        10'b0100100100: data <= 14'h3fab; 
        10'b0100100101: data <= 14'h3fa0; 
        10'b0100100110: data <= 14'h3fd8; 
        10'b0100100111: data <= 14'h0007; 
        10'b0100101000: data <= 14'h000a; 
        10'b0100101001: data <= 14'h0002; 
        10'b0100101010: data <= 14'h0005; 
        10'b0100101011: data <= 14'h3ff8; 
        10'b0100101100: data <= 14'h3ffa; 
        10'b0100101101: data <= 14'h3ff8; 
        10'b0100101110: data <= 14'h3fec; 
        10'b0100101111: data <= 14'h3fd1; 
        10'b0100110000: data <= 14'h3fe6; 
        10'b0100110001: data <= 14'h3fff; 
        10'b0100110010: data <= 14'h3fff; 
        10'b0100110011: data <= 14'h3ff5; 
        10'b0100110100: data <= 14'h3ff3; 
        10'b0100110101: data <= 14'h0003; 
        10'b0100110110: data <= 14'h3fff; 
        10'b0100110111: data <= 14'h3ff4; 
        10'b0100111000: data <= 14'h3fe8; 
        10'b0100111001: data <= 14'h3fcc; 
        10'b0100111010: data <= 14'h3fa6; 
        10'b0100111011: data <= 14'h3f81; 
        10'b0100111100: data <= 14'h3f86; 
        10'b0100111101: data <= 14'h3f71; 
        10'b0100111110: data <= 14'h3f70; 
        10'b0100111111: data <= 14'h3f7d; 
        10'b0101000000: data <= 14'h3f75; 
        10'b0101000001: data <= 14'h3f56; 
        10'b0101000010: data <= 14'h3f7d; 
        10'b0101000011: data <= 14'h3fc2; 
        10'b0101000100: data <= 14'h3fea; 
        10'b0101000101: data <= 14'h3fed; 
        10'b0101000110: data <= 14'h3fee; 
        10'b0101000111: data <= 14'h3ffc; 
        10'b0101001000: data <= 14'h3ff5; 
        10'b0101001001: data <= 14'h3ff5; 
        10'b0101001010: data <= 14'h3fe2; 
        10'b0101001011: data <= 14'h3fec; 
        10'b0101001100: data <= 14'h3ffc; 
        10'b0101001101: data <= 14'h3ff9; 
        10'b0101001110: data <= 14'h3ff5; 
        10'b0101001111: data <= 14'h3ffd; 
        10'b0101010000: data <= 14'h3ffb; 
        10'b0101010001: data <= 14'h3ffc; 
        10'b0101010010: data <= 14'h0001; 
        10'b0101010011: data <= 14'h3ffa; 
        10'b0101010100: data <= 14'h3fe6; 
        10'b0101010101: data <= 14'h3fb2; 
        10'b0101010110: data <= 14'h3f68; 
        10'b0101010111: data <= 14'h3f46; 
        10'b0101011000: data <= 14'h3f53; 
        10'b0101011001: data <= 14'h3f5c; 
        10'b0101011010: data <= 14'h3f6a; 
        10'b0101011011: data <= 14'h3f74; 
        10'b0101011100: data <= 14'h3f74; 
        10'b0101011101: data <= 14'h3f6e; 
        10'b0101011110: data <= 14'h3f88; 
        10'b0101011111: data <= 14'h3fb0; 
        10'b0101100000: data <= 14'h3fc9; 
        10'b0101100001: data <= 14'h3fcf; 
        10'b0101100010: data <= 14'h3fe7; 
        10'b0101100011: data <= 14'h0000; 
        10'b0101100100: data <= 14'h0000; 
        10'b0101100101: data <= 14'h3ff2; 
        10'b0101100110: data <= 14'h3fe0; 
        10'b0101100111: data <= 14'h3fd0; 
        10'b0101101000: data <= 14'h3ffa; 
        10'b0101101001: data <= 14'h3ff8; 
        10'b0101101010: data <= 14'h0004; 
        10'b0101101011: data <= 14'h3ffc; 
        10'b0101101100: data <= 14'h3ff6; 
        10'b0101101101: data <= 14'h3ffa; 
        10'b0101101110: data <= 14'h0003; 
        10'b0101101111: data <= 14'h3ff6; 
        10'b0101110000: data <= 14'h3fd6; 
        10'b0101110001: data <= 14'h3f9e; 
        10'b0101110010: data <= 14'h3f64; 
        10'b0101110011: data <= 14'h3f71; 
        10'b0101110100: data <= 14'h3f7a; 
        10'b0101110101: data <= 14'h3fa4; 
        10'b0101110110: data <= 14'h3fbf; 
        10'b0101110111: data <= 14'h3fe1; 
        10'b0101111000: data <= 14'h3fd0; 
        10'b0101111001: data <= 14'h3fea; 
        10'b0101111010: data <= 14'h3fc9; 
        10'b0101111011: data <= 14'h3fc8; 
        10'b0101111100: data <= 14'h3fbd; 
        10'b0101111101: data <= 14'h3fd0; 
        10'b0101111110: data <= 14'h3fe5; 
        10'b0101111111: data <= 14'h3ffb; 
        10'b0110000000: data <= 14'h3ff8; 
        10'b0110000001: data <= 14'h3fef; 
        10'b0110000010: data <= 14'h3fd8; 
        10'b0110000011: data <= 14'h3fdc; 
        10'b0110000100: data <= 14'h3fee; 
        10'b0110000101: data <= 14'h0005; 
        10'b0110000110: data <= 14'h3ffa; 
        10'b0110000111: data <= 14'h0000; 
        10'b0110001000: data <= 14'h0002; 
        10'b0110001001: data <= 14'h3ffd; 
        10'b0110001010: data <= 14'h0000; 
        10'b0110001011: data <= 14'h3ff8; 
        10'b0110001100: data <= 14'h3ff0; 
        10'b0110001101: data <= 14'h3fbe; 
        10'b0110001110: data <= 14'h3fac; 
        10'b0110001111: data <= 14'h3fbb; 
        10'b0110010000: data <= 14'h3fe5; 
        10'b0110010001: data <= 14'h3ffb; 
        10'b0110010010: data <= 14'h0011; 
        10'b0110010011: data <= 14'h0017; 
        10'b0110010100: data <= 14'h001b; 
        10'b0110010101: data <= 14'h002a; 
        10'b0110010110: data <= 14'h0003; 
        10'b0110010111: data <= 14'h3fe5; 
        10'b0110011000: data <= 14'h3fec; 
        10'b0110011001: data <= 14'h3fdd; 
        10'b0110011010: data <= 14'h3ffa; 
        10'b0110011011: data <= 14'h3fea; 
        10'b0110011100: data <= 14'h3ff9; 
        10'b0110011101: data <= 14'h3fe6; 
        10'b0110011110: data <= 14'h3fd2; 
        10'b0110011111: data <= 14'h3fdf; 
        10'b0110100000: data <= 14'h3ff9; 
        10'b0110100001: data <= 14'h0010; 
        10'b0110100010: data <= 14'h0012; 
        10'b0110100011: data <= 14'h3ff6; 
        10'b0110100100: data <= 14'h3ff9; 
        10'b0110100101: data <= 14'h3ffa; 
        10'b0110100110: data <= 14'h3ff9; 
        10'b0110100111: data <= 14'h000f; 
        10'b0110101000: data <= 14'h0007; 
        10'b0110101001: data <= 14'h0003; 
        10'b0110101010: data <= 14'h0012; 
        10'b0110101011: data <= 14'h0015; 
        10'b0110101100: data <= 14'h0027; 
        10'b0110101101: data <= 14'h001c; 
        10'b0110101110: data <= 14'h0021; 
        10'b0110101111: data <= 14'h0013; 
        10'b0110110000: data <= 14'h0011; 
        10'b0110110001: data <= 14'h0028; 
        10'b0110110010: data <= 14'h0003; 
        10'b0110110011: data <= 14'h0010; 
        10'b0110110100: data <= 14'h0002; 
        10'b0110110101: data <= 14'h3fe0; 
        10'b0110110110: data <= 14'h3fe1; 
        10'b0110110111: data <= 14'h3fed; 
        10'b0110111000: data <= 14'h3ff2; 
        10'b0110111001: data <= 14'h3feb; 
        10'b0110111010: data <= 14'h3fd6; 
        10'b0110111011: data <= 14'h3feb; 
        10'b0110111100: data <= 14'h000d; 
        10'b0110111101: data <= 14'h0016; 
        10'b0110111110: data <= 14'h000c; 
        10'b0110111111: data <= 14'h3ff4; 
        10'b0111000000: data <= 14'h3ff7; 
        10'b0111000001: data <= 14'h3ff2; 
        10'b0111000010: data <= 14'h3ff0; 
        10'b0111000011: data <= 14'h0010; 
        10'b0111000100: data <= 14'h0022; 
        10'b0111000101: data <= 14'h0037; 
        10'b0111000110: data <= 14'h0038; 
        10'b0111000111: data <= 14'h0022; 
        10'b0111001000: data <= 14'h000e; 
        10'b0111001001: data <= 14'h001d; 
        10'b0111001010: data <= 14'h001b; 
        10'b0111001011: data <= 14'h0019; 
        10'b0111001100: data <= 14'h0033; 
        10'b0111001101: data <= 14'h002d; 
        10'b0111001110: data <= 14'h0009; 
        10'b0111001111: data <= 14'h3ffb; 
        10'b0111010000: data <= 14'h0000; 
        10'b0111010001: data <= 14'h3feb; 
        10'b0111010010: data <= 14'h3fee; 
        10'b0111010011: data <= 14'h3fe0; 
        10'b0111010100: data <= 14'h3ff5; 
        10'b0111010101: data <= 14'h0002; 
        10'b0111010110: data <= 14'h0007; 
        10'b0111010111: data <= 14'h000f; 
        10'b0111011000: data <= 14'h002f; 
        10'b0111011001: data <= 14'h003a; 
        10'b0111011010: data <= 14'h000a; 
        10'b0111011011: data <= 14'h3ff7; 
        10'b0111011100: data <= 14'h3ff8; 
        10'b0111011101: data <= 14'h0003; 
        10'b0111011110: data <= 14'h3ffa; 
        10'b0111011111: data <= 14'h0014; 
        10'b0111100000: data <= 14'h003a; 
        10'b0111100001: data <= 14'h0051; 
        10'b0111100010: data <= 14'h004a; 
        10'b0111100011: data <= 14'h0032; 
        10'b0111100100: data <= 14'h0023; 
        10'b0111100101: data <= 14'h002b; 
        10'b0111100110: data <= 14'h0041; 
        10'b0111100111: data <= 14'h0036; 
        10'b0111101000: data <= 14'h003e; 
        10'b0111101001: data <= 14'h001d; 
        10'b0111101010: data <= 14'h000f; 
        10'b0111101011: data <= 14'h0014; 
        10'b0111101100: data <= 14'h0014; 
        10'b0111101101: data <= 14'h3ffd; 
        10'b0111101110: data <= 14'h000d; 
        10'b0111101111: data <= 14'h3ff8; 
        10'b0111110000: data <= 14'h0018; 
        10'b0111110001: data <= 14'h001a; 
        10'b0111110010: data <= 14'h0013; 
        10'b0111110011: data <= 14'h001b; 
        10'b0111110100: data <= 14'h004c; 
        10'b0111110101: data <= 14'h0042; 
        10'b0111110110: data <= 14'h000f; 
        10'b0111110111: data <= 14'h0002; 
        10'b0111111000: data <= 14'h3ffe; 
        10'b0111111001: data <= 14'h3fff; 
        10'b0111111010: data <= 14'h3fec; 
        10'b0111111011: data <= 14'h0005; 
        10'b0111111100: data <= 14'h003f; 
        10'b0111111101: data <= 14'h006a; 
        10'b0111111110: data <= 14'h0064; 
        10'b0111111111: data <= 14'h0048; 
        10'b1000000000: data <= 14'h0030; 
        10'b1000000001: data <= 14'h0035; 
        10'b1000000010: data <= 14'h0051; 
        10'b1000000011: data <= 14'h0049; 
        10'b1000000100: data <= 14'h0075; 
        10'b1000000101: data <= 14'h0055; 
        10'b1000000110: data <= 14'h004b; 
        10'b1000000111: data <= 14'h0024; 
        10'b1000001000: data <= 14'h0019; 
        10'b1000001001: data <= 14'h002e; 
        10'b1000001010: data <= 14'h001e; 
        10'b1000001011: data <= 14'h0014; 
        10'b1000001100: data <= 14'h0036; 
        10'b1000001101: data <= 14'h0038; 
        10'b1000001110: data <= 14'h003d; 
        10'b1000001111: data <= 14'h0051; 
        10'b1000010000: data <= 14'h0064; 
        10'b1000010001: data <= 14'h003a; 
        10'b1000010010: data <= 14'h3ffa; 
        10'b1000010011: data <= 14'h3ff4; 
        10'b1000010100: data <= 14'h3ff6; 
        10'b1000010101: data <= 14'h3ff7; 
        10'b1000010110: data <= 14'h3ff2; 
        10'b1000010111: data <= 14'h0000; 
        10'b1000011000: data <= 14'h0022; 
        10'b1000011001: data <= 14'h0040; 
        10'b1000011010: data <= 14'h0051; 
        10'b1000011011: data <= 14'h0046; 
        10'b1000011100: data <= 14'h0041; 
        10'b1000011101: data <= 14'h0045; 
        10'b1000011110: data <= 14'h0042; 
        10'b1000011111: data <= 14'h0046; 
        10'b1000100000: data <= 14'h004e; 
        10'b1000100001: data <= 14'h003c; 
        10'b1000100010: data <= 14'h0027; 
        10'b1000100011: data <= 14'h0013; 
        10'b1000100100: data <= 14'h001d; 
        10'b1000100101: data <= 14'h0032; 
        10'b1000100110: data <= 14'h0018; 
        10'b1000100111: data <= 14'h0018; 
        10'b1000101000: data <= 14'h0028; 
        10'b1000101001: data <= 14'h0032; 
        10'b1000101010: data <= 14'h0042; 
        10'b1000101011: data <= 14'h0046; 
        10'b1000101100: data <= 14'h003d; 
        10'b1000101101: data <= 14'h0020; 
        10'b1000101110: data <= 14'h0003; 
        10'b1000101111: data <= 14'h0001; 
        10'b1000110000: data <= 14'h3ff3; 
        10'b1000110001: data <= 14'h3fff; 
        10'b1000110010: data <= 14'h3ffd; 
        10'b1000110011: data <= 14'h3fef; 
        10'b1000110100: data <= 14'h001f; 
        10'b1000110101: data <= 14'h0026; 
        10'b1000110110: data <= 14'h003b; 
        10'b1000110111: data <= 14'h0052; 
        10'b1000111000: data <= 14'h004d; 
        10'b1000111001: data <= 14'h0033; 
        10'b1000111010: data <= 14'h0031; 
        10'b1000111011: data <= 14'h0053; 
        10'b1000111100: data <= 14'h002e; 
        10'b1000111101: data <= 14'h000f; 
        10'b1000111110: data <= 14'h000a; 
        10'b1000111111: data <= 14'h000d; 
        10'b1001000000: data <= 14'h0010; 
        10'b1001000001: data <= 14'h0001; 
        10'b1001000010: data <= 14'h0024; 
        10'b1001000011: data <= 14'h0038; 
        10'b1001000100: data <= 14'h0026; 
        10'b1001000101: data <= 14'h0036; 
        10'b1001000110: data <= 14'h004b; 
        10'b1001000111: data <= 14'h0041; 
        10'b1001001000: data <= 14'h002f; 
        10'b1001001001: data <= 14'h0016; 
        10'b1001001010: data <= 14'h0000; 
        10'b1001001011: data <= 14'h3ffe; 
        10'b1001001100: data <= 14'h3ffb; 
        10'b1001001101: data <= 14'h3ff4; 
        10'b1001001110: data <= 14'h3ffe; 
        10'b1001001111: data <= 14'h3ff9; 
        10'b1001010000: data <= 14'h0006; 
        10'b1001010001: data <= 14'h0010; 
        10'b1001010010: data <= 14'h0029; 
        10'b1001010011: data <= 14'h002e; 
        10'b1001010100: data <= 14'h0028; 
        10'b1001010101: data <= 14'h0032; 
        10'b1001010110: data <= 14'h002c; 
        10'b1001010111: data <= 14'h002c; 
        10'b1001011000: data <= 14'h0011; 
        10'b1001011001: data <= 14'h0008; 
        10'b1001011010: data <= 14'h3ffc; 
        10'b1001011011: data <= 14'h0002; 
        10'b1001011100: data <= 14'h0016; 
        10'b1001011101: data <= 14'h0018; 
        10'b1001011110: data <= 14'h0034; 
        10'b1001011111: data <= 14'h0037; 
        10'b1001100000: data <= 14'h0018; 
        10'b1001100001: data <= 14'h0036; 
        10'b1001100010: data <= 14'h0042; 
        10'b1001100011: data <= 14'h004c; 
        10'b1001100100: data <= 14'h0025; 
        10'b1001100101: data <= 14'h000f; 
        10'b1001100110: data <= 14'h0003; 
        10'b1001100111: data <= 14'h3ffe; 
        10'b1001101000: data <= 14'h3ff3; 
        10'b1001101001: data <= 14'h3ffd; 
        10'b1001101010: data <= 14'h3ff5; 
        10'b1001101011: data <= 14'h0004; 
        10'b1001101100: data <= 14'h000d; 
        10'b1001101101: data <= 14'h0005; 
        10'b1001101110: data <= 14'h001c; 
        10'b1001101111: data <= 14'h0018; 
        10'b1001110000: data <= 14'h0017; 
        10'b1001110001: data <= 14'h0020; 
        10'b1001110010: data <= 14'h0020; 
        10'b1001110011: data <= 14'h0025; 
        10'b1001110100: data <= 14'h0004; 
        10'b1001110101: data <= 14'h3fe2; 
        10'b1001110110: data <= 14'h3fdb; 
        10'b1001110111: data <= 14'h3feb; 
        10'b1001111000: data <= 14'h3fec; 
        10'b1001111001: data <= 14'h000f; 
        10'b1001111010: data <= 14'h0030; 
        10'b1001111011: data <= 14'h003e; 
        10'b1001111100: data <= 14'h0038; 
        10'b1001111101: data <= 14'h0036; 
        10'b1001111110: data <= 14'h002f; 
        10'b1001111111: data <= 14'h0034; 
        10'b1010000000: data <= 14'h0013; 
        10'b1010000001: data <= 14'h3ffe; 
        10'b1010000010: data <= 14'h3ffd; 
        10'b1010000011: data <= 14'h3ff7; 
        10'b1010000100: data <= 14'h3ffd; 
        10'b1010000101: data <= 14'h3ffd; 
        10'b1010000110: data <= 14'h3ffa; 
        10'b1010000111: data <= 14'h3ffa; 
        10'b1010001000: data <= 14'h3ff9; 
        10'b1010001001: data <= 14'h3ff2; 
        10'b1010001010: data <= 14'h3fee; 
        10'b1010001011: data <= 14'h3ff1; 
        10'b1010001100: data <= 14'h3fe7; 
        10'b1010001101: data <= 14'h3ff1; 
        10'b1010001110: data <= 14'h3ff6; 
        10'b1010001111: data <= 14'h000d; 
        10'b1010010000: data <= 14'h0001; 
        10'b1010010001: data <= 14'h3fec; 
        10'b1010010010: data <= 14'h3fe5; 
        10'b1010010011: data <= 14'h3fdd; 
        10'b1010010100: data <= 14'h3fda; 
        10'b1010010101: data <= 14'h3fec; 
        10'b1010010110: data <= 14'h0008; 
        10'b1010010111: data <= 14'h0030; 
        10'b1010011000: data <= 14'h002a; 
        10'b1010011001: data <= 14'h0034; 
        10'b1010011010: data <= 14'h0025; 
        10'b1010011011: data <= 14'h000e; 
        10'b1010011100: data <= 14'h0009; 
        10'b1010011101: data <= 14'h0005; 
        10'b1010011110: data <= 14'h3fff; 
        10'b1010011111: data <= 14'h3ff9; 
        10'b1010100000: data <= 14'h3ffb; 
        10'b1010100001: data <= 14'h3ff6; 
        10'b1010100010: data <= 14'h0000; 
        10'b1010100011: data <= 14'h3ffe; 
        10'b1010100100: data <= 14'h3ff6; 
        10'b1010100101: data <= 14'h3fe5; 
        10'b1010100110: data <= 14'h3fcc; 
        10'b1010100111: data <= 14'h3fd9; 
        10'b1010101000: data <= 14'h3fd8; 
        10'b1010101001: data <= 14'h3fd5; 
        10'b1010101010: data <= 14'h3fd5; 
        10'b1010101011: data <= 14'h3fdf; 
        10'b1010101100: data <= 14'h3fdf; 
        10'b1010101101: data <= 14'h3fee; 
        10'b1010101110: data <= 14'h3fe9; 
        10'b1010101111: data <= 14'h3fdf; 
        10'b1010110000: data <= 14'h3fe0; 
        10'b1010110001: data <= 14'h3fe7; 
        10'b1010110010: data <= 14'h3fe2; 
        10'b1010110011: data <= 14'h3ff0; 
        10'b1010110100: data <= 14'h3ff2; 
        10'b1010110101: data <= 14'h3ff2; 
        10'b1010110110: data <= 14'h3ff8; 
        10'b1010110111: data <= 14'h3ff9; 
        10'b1010111000: data <= 14'h3fff; 
        10'b1010111001: data <= 14'h0005; 
        10'b1010111010: data <= 14'h3ff5; 
        10'b1010111011: data <= 14'h3ff5; 
        10'b1010111100: data <= 14'h0000; 
        10'b1010111101: data <= 14'h3ff2; 
        10'b1010111110: data <= 14'h3ff9; 
        10'b1010111111: data <= 14'h3ff7; 
        10'b1011000000: data <= 14'h3ff5; 
        10'b1011000001: data <= 14'h3fed; 
        10'b1011000010: data <= 14'h3fe7; 
        10'b1011000011: data <= 14'h3fd9; 
        10'b1011000100: data <= 14'h3fd5; 
        10'b1011000101: data <= 14'h3fd8; 
        10'b1011000110: data <= 14'h3fdc; 
        10'b1011000111: data <= 14'h3fd2; 
        10'b1011001000: data <= 14'h3fe1; 
        10'b1011001001: data <= 14'h3fe3; 
        10'b1011001010: data <= 14'h3fda; 
        10'b1011001011: data <= 14'h3fe0; 
        10'b1011001100: data <= 14'h3fe9; 
        10'b1011001101: data <= 14'h3fea; 
        10'b1011001110: data <= 14'h3ff8; 
        10'b1011001111: data <= 14'h3fec; 
        10'b1011010000: data <= 14'h3ff9; 
        10'b1011010001: data <= 14'h3ff8; 
        10'b1011010010: data <= 14'h0000; 
        10'b1011010011: data <= 14'h3ff5; 
        10'b1011010100: data <= 14'h3ffc; 
        10'b1011010101: data <= 14'h3ff5; 
        10'b1011010110: data <= 14'h3ff2; 
        10'b1011010111: data <= 14'h3ff6; 
        10'b1011011000: data <= 14'h3ff3; 
        10'b1011011001: data <= 14'h3ff8; 
        10'b1011011010: data <= 14'h3ffa; 
        10'b1011011011: data <= 14'h0001; 
        10'b1011011100: data <= 14'h3ffe; 
        10'b1011011101: data <= 14'h3ff9; 
        10'b1011011110: data <= 14'h3ffd; 
        10'b1011011111: data <= 14'h0000; 
        10'b1011100000: data <= 14'h3ff9; 
        10'b1011100001: data <= 14'h0001; 
        10'b1011100010: data <= 14'h0000; 
        10'b1011100011: data <= 14'h0000; 
        10'b1011100100: data <= 14'h0001; 
        10'b1011100101: data <= 14'h3ffc; 
        10'b1011100110: data <= 14'h3ff7; 
        10'b1011100111: data <= 14'h3ff1; 
        10'b1011101000: data <= 14'h3ff8; 
        10'b1011101001: data <= 14'h3ffc; 
        10'b1011101010: data <= 14'h3ffb; 
        10'b1011101011: data <= 14'h3ff5; 
        10'b1011101100: data <= 14'h0001; 
        10'b1011101101: data <= 14'h0000; 
        10'b1011101110: data <= 14'h3ff5; 
        10'b1011101111: data <= 14'h3ff8; 
        10'b1011110000: data <= 14'h3ff3; 
        10'b1011110001: data <= 14'h0001; 
        10'b1011110010: data <= 14'h0000; 
        10'b1011110011: data <= 14'h3fff; 
        10'b1011110100: data <= 14'h3fff; 
        10'b1011110101: data <= 14'h3ff6; 
        10'b1011110110: data <= 14'h3ff4; 
        10'b1011110111: data <= 14'h3ffb; 
        10'b1011111000: data <= 14'h3ff2; 
        10'b1011111001: data <= 14'h0003; 
        10'b1011111010: data <= 14'h0003; 
        10'b1011111011: data <= 14'h3ff8; 
        10'b1011111100: data <= 14'h3fff; 
        10'b1011111101: data <= 14'h3ff5; 
        10'b1011111110: data <= 14'h0002; 
        10'b1011111111: data <= 14'h3ff2; 
        10'b1100000000: data <= 14'h3fff; 
        10'b1100000001: data <= 14'h3ff9; 
        10'b1100000010: data <= 14'h3ffd; 
        10'b1100000011: data <= 14'h3ff4; 
        10'b1100000100: data <= 14'h3ffb; 
        10'b1100000101: data <= 14'h3ff9; 
        10'b1100000110: data <= 14'h3ffc; 
        10'b1100000111: data <= 14'h3ffb; 
        10'b1100001000: data <= 14'h3ffe; 
        10'b1100001001: data <= 14'h3ff1; 
        10'b1100001010: data <= 14'h3ffa; 
        10'b1100001011: data <= 14'h0000; 
        10'b1100001100: data <= 14'h3ff1; 
        10'b1100001101: data <= 14'h3ffb; 
        10'b1100001110: data <= 14'h3ffe; 
        10'b1100001111: data <= 14'h3ff8; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 9) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 15'h7fe6; 
        10'b0000000001: data <= 15'h0001; 
        10'b0000000010: data <= 15'h7ff3; 
        10'b0000000011: data <= 15'h7feb; 
        10'b0000000100: data <= 15'h7ff3; 
        10'b0000000101: data <= 15'h7fec; 
        10'b0000000110: data <= 15'h7ff7; 
        10'b0000000111: data <= 15'h7ff9; 
        10'b0000001000: data <= 15'h7fe6; 
        10'b0000001001: data <= 15'h7ff5; 
        10'b0000001010: data <= 15'h7fe7; 
        10'b0000001011: data <= 15'h7ff0; 
        10'b0000001100: data <= 15'h0005; 
        10'b0000001101: data <= 15'h0004; 
        10'b0000001110: data <= 15'h7fe7; 
        10'b0000001111: data <= 15'h7ff7; 
        10'b0000010000: data <= 15'h7fe9; 
        10'b0000010001: data <= 15'h7fe9; 
        10'b0000010010: data <= 15'h0007; 
        10'b0000010011: data <= 15'h0002; 
        10'b0000010100: data <= 15'h7fed; 
        10'b0000010101: data <= 15'h7ff8; 
        10'b0000010110: data <= 15'h7fef; 
        10'b0000010111: data <= 15'h7fe4; 
        10'b0000011000: data <= 15'h7fe6; 
        10'b0000011001: data <= 15'h7ff6; 
        10'b0000011010: data <= 15'h7fff; 
        10'b0000011011: data <= 15'h7ff9; 
        10'b0000011100: data <= 15'h7ff5; 
        10'b0000011101: data <= 15'h7ff3; 
        10'b0000011110: data <= 15'h0006; 
        10'b0000011111: data <= 15'h7ffa; 
        10'b0000100000: data <= 15'h7fe8; 
        10'b0000100001: data <= 15'h7fe7; 
        10'b0000100010: data <= 15'h7fe6; 
        10'b0000100011: data <= 15'h7fec; 
        10'b0000100100: data <= 15'h7fec; 
        10'b0000100101: data <= 15'h7ff7; 
        10'b0000100110: data <= 15'h0000; 
        10'b0000100111: data <= 15'h7fe9; 
        10'b0000101000: data <= 15'h7ff1; 
        10'b0000101001: data <= 15'h7fe8; 
        10'b0000101010: data <= 15'h7ff7; 
        10'b0000101011: data <= 15'h7fe4; 
        10'b0000101100: data <= 15'h7ff9; 
        10'b0000101101: data <= 15'h7fe9; 
        10'b0000101110: data <= 15'h7ff0; 
        10'b0000101111: data <= 15'h7fea; 
        10'b0000110000: data <= 15'h7ff7; 
        10'b0000110001: data <= 15'h7fe9; 
        10'b0000110010: data <= 15'h7fe5; 
        10'b0000110011: data <= 15'h7fe3; 
        10'b0000110100: data <= 15'h0001; 
        10'b0000110101: data <= 15'h7ffa; 
        10'b0000110110: data <= 15'h0002; 
        10'b0000110111: data <= 15'h7fee; 
        10'b0000111000: data <= 15'h7ff4; 
        10'b0000111001: data <= 15'h7fe4; 
        10'b0000111010: data <= 15'h7fe7; 
        10'b0000111011: data <= 15'h0000; 
        10'b0000111100: data <= 15'h7fe5; 
        10'b0000111101: data <= 15'h7fe8; 
        10'b0000111110: data <= 15'h7ff2; 
        10'b0000111111: data <= 15'h7ff6; 
        10'b0001000000: data <= 15'h7ffd; 
        10'b0001000001: data <= 15'h7ff1; 
        10'b0001000010: data <= 15'h000e; 
        10'b0001000011: data <= 15'h000c; 
        10'b0001000100: data <= 15'h0025; 
        10'b0001000101: data <= 15'h001d; 
        10'b0001000110: data <= 15'h001b; 
        10'b0001000111: data <= 15'h000b; 
        10'b0001001000: data <= 15'h0024; 
        10'b0001001001: data <= 15'h000c; 
        10'b0001001010: data <= 15'h000b; 
        10'b0001001011: data <= 15'h7fee; 
        10'b0001001100: data <= 15'h7fff; 
        10'b0001001101: data <= 15'h7ff7; 
        10'b0001001110: data <= 15'h7fda; 
        10'b0001001111: data <= 15'h7ff3; 
        10'b0001010000: data <= 15'h7ffc; 
        10'b0001010001: data <= 15'h0009; 
        10'b0001010010: data <= 15'h7ff5; 
        10'b0001010011: data <= 15'h7ff1; 
        10'b0001010100: data <= 15'h7fee; 
        10'b0001010101: data <= 15'h7feb; 
        10'b0001010110: data <= 15'h7ffa; 
        10'b0001010111: data <= 15'h7fed; 
        10'b0001011000: data <= 15'h0005; 
        10'b0001011001: data <= 15'h7fe9; 
        10'b0001011010: data <= 15'h7ff8; 
        10'b0001011011: data <= 15'h0000; 
        10'b0001011100: data <= 15'h0007; 
        10'b0001011101: data <= 15'h003b; 
        10'b0001011110: data <= 15'h005c; 
        10'b0001011111: data <= 15'h005c; 
        10'b0001100000: data <= 15'h0058; 
        10'b0001100001: data <= 15'h0081; 
        10'b0001100010: data <= 15'h0046; 
        10'b0001100011: data <= 15'h001f; 
        10'b0001100100: data <= 15'h003b; 
        10'b0001100101: data <= 15'h001b; 
        10'b0001100110: data <= 15'h7fe6; 
        10'b0001100111: data <= 15'h7ffa; 
        10'b0001101000: data <= 15'h7fe3; 
        10'b0001101001: data <= 15'h7fde; 
        10'b0001101010: data <= 15'h7fd6; 
        10'b0001101011: data <= 15'h7feb; 
        10'b0001101100: data <= 15'h0003; 
        10'b0001101101: data <= 15'h000a; 
        10'b0001101110: data <= 15'h7fe9; 
        10'b0001101111: data <= 15'h7ffb; 
        10'b0001110000: data <= 15'h7fec; 
        10'b0001110001: data <= 15'h7ff2; 
        10'b0001110010: data <= 15'h0007; 
        10'b0001110011: data <= 15'h7fe2; 
        10'b0001110100: data <= 15'h7fe5; 
        10'b0001110101: data <= 15'h7ff8; 
        10'b0001110110: data <= 15'h000e; 
        10'b0001110111: data <= 15'h000d; 
        10'b0001111000: data <= 15'h0026; 
        10'b0001111001: data <= 15'h0071; 
        10'b0001111010: data <= 15'h0072; 
        10'b0001111011: data <= 15'h008f; 
        10'b0001111100: data <= 15'h0079; 
        10'b0001111101: data <= 15'h0060; 
        10'b0001111110: data <= 15'h0057; 
        10'b0001111111: data <= 15'h0027; 
        10'b0010000000: data <= 15'h0034; 
        10'b0010000001: data <= 15'h0030; 
        10'b0010000010: data <= 15'h7ff2; 
        10'b0010000011: data <= 15'h7fe8; 
        10'b0010000100: data <= 15'h7fed; 
        10'b0010000101: data <= 15'h7fc7; 
        10'b0010000110: data <= 15'h7fbb; 
        10'b0010000111: data <= 15'h7fbe; 
        10'b0010001000: data <= 15'h7ff8; 
        10'b0010001001: data <= 15'h7ff8; 
        10'b0010001010: data <= 15'h7fe4; 
        10'b0010001011: data <= 15'h7ffb; 
        10'b0010001100: data <= 15'h0002; 
        10'b0010001101: data <= 15'h7ff7; 
        10'b0010001110: data <= 15'h7fea; 
        10'b0010001111: data <= 15'h7fe3; 
        10'b0010010000: data <= 15'h7fe8; 
        10'b0010010001: data <= 15'h7fec; 
        10'b0010010010: data <= 15'h000d; 
        10'b0010010011: data <= 15'h0037; 
        10'b0010010100: data <= 15'h004c; 
        10'b0010010101: data <= 15'h0083; 
        10'b0010010110: data <= 15'h0091; 
        10'b0010010111: data <= 15'h0097; 
        10'b0010011000: data <= 15'h008a; 
        10'b0010011001: data <= 15'h009b; 
        10'b0010011010: data <= 15'h0090; 
        10'b0010011011: data <= 15'h0085; 
        10'b0010011100: data <= 15'h0091; 
        10'b0010011101: data <= 15'h0075; 
        10'b0010011110: data <= 15'h0055; 
        10'b0010011111: data <= 15'h7fdc; 
        10'b0010100000: data <= 15'h7fde; 
        10'b0010100001: data <= 15'h7fc8; 
        10'b0010100010: data <= 15'h7fc7; 
        10'b0010100011: data <= 15'h7fa7; 
        10'b0010100100: data <= 15'h7fda; 
        10'b0010100101: data <= 15'h7fea; 
        10'b0010100110: data <= 15'h0004; 
        10'b0010100111: data <= 15'h7fef; 
        10'b0010101000: data <= 15'h7ff4; 
        10'b0010101001: data <= 15'h7feb; 
        10'b0010101010: data <= 15'h0005; 
        10'b0010101011: data <= 15'h7ff5; 
        10'b0010101100: data <= 15'h7ff1; 
        10'b0010101101: data <= 15'h0009; 
        10'b0010101110: data <= 15'h0036; 
        10'b0010101111: data <= 15'h0068; 
        10'b0010110000: data <= 15'h0050; 
        10'b0010110001: data <= 15'h005b; 
        10'b0010110010: data <= 15'h007b; 
        10'b0010110011: data <= 15'h004d; 
        10'b0010110100: data <= 15'h0051; 
        10'b0010110101: data <= 15'h0069; 
        10'b0010110110: data <= 15'h005d; 
        10'b0010110111: data <= 15'h0033; 
        10'b0010111000: data <= 15'h0038; 
        10'b0010111001: data <= 15'h000e; 
        10'b0010111010: data <= 15'h000b; 
        10'b0010111011: data <= 15'h7fdf; 
        10'b0010111100: data <= 15'h7fea; 
        10'b0010111101: data <= 15'h7fb8; 
        10'b0010111110: data <= 15'h7fb9; 
        10'b0010111111: data <= 15'h7f9d; 
        10'b0011000000: data <= 15'h7fc5; 
        10'b0011000001: data <= 15'h7fdf; 
        10'b0011000010: data <= 15'h0004; 
        10'b0011000011: data <= 15'h7ffd; 
        10'b0011000100: data <= 15'h7ff1; 
        10'b0011000101: data <= 15'h0003; 
        10'b0011000110: data <= 15'h0003; 
        10'b0011000111: data <= 15'h7ff2; 
        10'b0011001000: data <= 15'h0001; 
        10'b0011001001: data <= 15'h001d; 
        10'b0011001010: data <= 15'h0045; 
        10'b0011001011: data <= 15'h0065; 
        10'b0011001100: data <= 15'h0052; 
        10'b0011001101: data <= 15'h004d; 
        10'b0011001110: data <= 15'h001d; 
        10'b0011001111: data <= 15'h0023; 
        10'b0011010000: data <= 15'h0006; 
        10'b0011010001: data <= 15'h0036; 
        10'b0011010010: data <= 15'h0042; 
        10'b0011010011: data <= 15'h000e; 
        10'b0011010100: data <= 15'h0009; 
        10'b0011010101: data <= 15'h7fac; 
        10'b0011010110: data <= 15'h7fe3; 
        10'b0011010111: data <= 15'h7fe8; 
        10'b0011011000: data <= 15'h7fe5; 
        10'b0011011001: data <= 15'h7fe0; 
        10'b0011011010: data <= 15'h7fe8; 
        10'b0011011011: data <= 15'h7fae; 
        10'b0011011100: data <= 15'h7fc7; 
        10'b0011011101: data <= 15'h7fef; 
        10'b0011011110: data <= 15'h7fea; 
        10'b0011011111: data <= 15'h7fe5; 
        10'b0011100000: data <= 15'h7ffa; 
        10'b0011100001: data <= 15'h0004; 
        10'b0011100010: data <= 15'h7ff5; 
        10'b0011100011: data <= 15'h0004; 
        10'b0011100100: data <= 15'h000f; 
        10'b0011100101: data <= 15'h002f; 
        10'b0011100110: data <= 15'h0022; 
        10'b0011100111: data <= 15'h0030; 
        10'b0011101000: data <= 15'h0031; 
        10'b0011101001: data <= 15'h0036; 
        10'b0011101010: data <= 15'h0036; 
        10'b0011101011: data <= 15'h003e; 
        10'b0011101100: data <= 15'h0025; 
        10'b0011101101: data <= 15'h002c; 
        10'b0011101110: data <= 15'h0074; 
        10'b0011101111: data <= 15'h0041; 
        10'b0011110000: data <= 15'h7ff8; 
        10'b0011110001: data <= 15'h7fe0; 
        10'b0011110010: data <= 15'h7fff; 
        10'b0011110011: data <= 15'h001a; 
        10'b0011110100: data <= 15'h0001; 
        10'b0011110101: data <= 15'h7fee; 
        10'b0011110110: data <= 15'h7fd1; 
        10'b0011110111: data <= 15'h7fa1; 
        10'b0011111000: data <= 15'h7fb7; 
        10'b0011111001: data <= 15'h7fe2; 
        10'b0011111010: data <= 15'h7ff2; 
        10'b0011111011: data <= 15'h7fe9; 
        10'b0011111100: data <= 15'h7fec; 
        10'b0011111101: data <= 15'h7ffb; 
        10'b0011111110: data <= 15'h7fff; 
        10'b0011111111: data <= 15'h000c; 
        10'b0100000000: data <= 15'h0018; 
        10'b0100000001: data <= 15'h0035; 
        10'b0100000010: data <= 15'h0012; 
        10'b0100000011: data <= 15'h0004; 
        10'b0100000100: data <= 15'h7fee; 
        10'b0100000101: data <= 15'h001c; 
        10'b0100000110: data <= 15'h0016; 
        10'b0100000111: data <= 15'h001c; 
        10'b0100001000: data <= 15'h0007; 
        10'b0100001001: data <= 15'h7ffd; 
        10'b0100001010: data <= 15'h004c; 
        10'b0100001011: data <= 15'h0052; 
        10'b0100001100: data <= 15'h001c; 
        10'b0100001101: data <= 15'h0002; 
        10'b0100001110: data <= 15'h7ff8; 
        10'b0100001111: data <= 15'h7fff; 
        10'b0100010000: data <= 15'h7ffd; 
        10'b0100010001: data <= 15'h7ffe; 
        10'b0100010010: data <= 15'h7fe2; 
        10'b0100010011: data <= 15'h7faf; 
        10'b0100010100: data <= 15'h7fbb; 
        10'b0100010101: data <= 15'h7fe9; 
        10'b0100010110: data <= 15'h0004; 
        10'b0100010111: data <= 15'h7fe6; 
        10'b0100011000: data <= 15'h0005; 
        10'b0100011001: data <= 15'h7ffa; 
        10'b0100011010: data <= 15'h7ff4; 
        10'b0100011011: data <= 15'h7fef; 
        10'b0100011100: data <= 15'h0004; 
        10'b0100011101: data <= 15'h7ff3; 
        10'b0100011110: data <= 15'h7fe6; 
        10'b0100011111: data <= 15'h7f80; 
        10'b0100100000: data <= 15'h7f8e; 
        10'b0100100001: data <= 15'h7faa; 
        10'b0100100010: data <= 15'h7f7c; 
        10'b0100100011: data <= 15'h7f6d; 
        10'b0100100100: data <= 15'h7f56; 
        10'b0100100101: data <= 15'h7f41; 
        10'b0100100110: data <= 15'h7fb0; 
        10'b0100100111: data <= 15'h000f; 
        10'b0100101000: data <= 15'h0015; 
        10'b0100101001: data <= 15'h0003; 
        10'b0100101010: data <= 15'h000b; 
        10'b0100101011: data <= 15'h7ff0; 
        10'b0100101100: data <= 15'h7ff5; 
        10'b0100101101: data <= 15'h7ff0; 
        10'b0100101110: data <= 15'h7fd8; 
        10'b0100101111: data <= 15'h7fa3; 
        10'b0100110000: data <= 15'h7fcd; 
        10'b0100110001: data <= 15'h7ffe; 
        10'b0100110010: data <= 15'h7ffe; 
        10'b0100110011: data <= 15'h7fea; 
        10'b0100110100: data <= 15'h7fe5; 
        10'b0100110101: data <= 15'h0007; 
        10'b0100110110: data <= 15'h7ffd; 
        10'b0100110111: data <= 15'h7fe8; 
        10'b0100111000: data <= 15'h7fd0; 
        10'b0100111001: data <= 15'h7f97; 
        10'b0100111010: data <= 15'h7f4c; 
        10'b0100111011: data <= 15'h7f03; 
        10'b0100111100: data <= 15'h7f0c; 
        10'b0100111101: data <= 15'h7ee1; 
        10'b0100111110: data <= 15'h7ee0; 
        10'b0100111111: data <= 15'h7ef9; 
        10'b0101000000: data <= 15'h7ee9; 
        10'b0101000001: data <= 15'h7eac; 
        10'b0101000010: data <= 15'h7efb; 
        10'b0101000011: data <= 15'h7f83; 
        10'b0101000100: data <= 15'h7fd5; 
        10'b0101000101: data <= 15'h7fdb; 
        10'b0101000110: data <= 15'h7fdc; 
        10'b0101000111: data <= 15'h7ff9; 
        10'b0101001000: data <= 15'h7fea; 
        10'b0101001001: data <= 15'h7fea; 
        10'b0101001010: data <= 15'h7fc5; 
        10'b0101001011: data <= 15'h7fd7; 
        10'b0101001100: data <= 15'h7ff9; 
        10'b0101001101: data <= 15'h7ff2; 
        10'b0101001110: data <= 15'h7fea; 
        10'b0101001111: data <= 15'h7ffa; 
        10'b0101010000: data <= 15'h7ff7; 
        10'b0101010001: data <= 15'h7ff8; 
        10'b0101010010: data <= 15'h0003; 
        10'b0101010011: data <= 15'h7ff5; 
        10'b0101010100: data <= 15'h7fcc; 
        10'b0101010101: data <= 15'h7f64; 
        10'b0101010110: data <= 15'h7ed1; 
        10'b0101010111: data <= 15'h7e8d; 
        10'b0101011000: data <= 15'h7ea6; 
        10'b0101011001: data <= 15'h7eb8; 
        10'b0101011010: data <= 15'h7ed4; 
        10'b0101011011: data <= 15'h7ee7; 
        10'b0101011100: data <= 15'h7ee8; 
        10'b0101011101: data <= 15'h7edd; 
        10'b0101011110: data <= 15'h7f11; 
        10'b0101011111: data <= 15'h7f60; 
        10'b0101100000: data <= 15'h7f93; 
        10'b0101100001: data <= 15'h7f9e; 
        10'b0101100010: data <= 15'h7fce; 
        10'b0101100011: data <= 15'h0000; 
        10'b0101100100: data <= 15'h7fff; 
        10'b0101100101: data <= 15'h7fe4; 
        10'b0101100110: data <= 15'h7fc1; 
        10'b0101100111: data <= 15'h7fa0; 
        10'b0101101000: data <= 15'h7ff4; 
        10'b0101101001: data <= 15'h7ff0; 
        10'b0101101010: data <= 15'h0007; 
        10'b0101101011: data <= 15'h7ff8; 
        10'b0101101100: data <= 15'h7fed; 
        10'b0101101101: data <= 15'h7ff3; 
        10'b0101101110: data <= 15'h0007; 
        10'b0101101111: data <= 15'h7fec; 
        10'b0101110000: data <= 15'h7fac; 
        10'b0101110001: data <= 15'h7f3b; 
        10'b0101110010: data <= 15'h7ec8; 
        10'b0101110011: data <= 15'h7ee1; 
        10'b0101110100: data <= 15'h7ef5; 
        10'b0101110101: data <= 15'h7f48; 
        10'b0101110110: data <= 15'h7f7e; 
        10'b0101110111: data <= 15'h7fc3; 
        10'b0101111000: data <= 15'h7fa0; 
        10'b0101111001: data <= 15'h7fd4; 
        10'b0101111010: data <= 15'h7f92; 
        10'b0101111011: data <= 15'h7f90; 
        10'b0101111100: data <= 15'h7f7b; 
        10'b0101111101: data <= 15'h7fa0; 
        10'b0101111110: data <= 15'h7fcb; 
        10'b0101111111: data <= 15'h7ff6; 
        10'b0110000000: data <= 15'h7ff0; 
        10'b0110000001: data <= 15'h7fde; 
        10'b0110000010: data <= 15'h7fb1; 
        10'b0110000011: data <= 15'h7fb8; 
        10'b0110000100: data <= 15'h7fdb; 
        10'b0110000101: data <= 15'h0009; 
        10'b0110000110: data <= 15'h7ff4; 
        10'b0110000111: data <= 15'h7fff; 
        10'b0110001000: data <= 15'h0004; 
        10'b0110001001: data <= 15'h7ff9; 
        10'b0110001010: data <= 15'h0001; 
        10'b0110001011: data <= 15'h7fef; 
        10'b0110001100: data <= 15'h7fe0; 
        10'b0110001101: data <= 15'h7f7b; 
        10'b0110001110: data <= 15'h7f58; 
        10'b0110001111: data <= 15'h7f77; 
        10'b0110010000: data <= 15'h7fc9; 
        10'b0110010001: data <= 15'h7ff7; 
        10'b0110010010: data <= 15'h0022; 
        10'b0110010011: data <= 15'h002d; 
        10'b0110010100: data <= 15'h0036; 
        10'b0110010101: data <= 15'h0054; 
        10'b0110010110: data <= 15'h0006; 
        10'b0110010111: data <= 15'h7fca; 
        10'b0110011000: data <= 15'h7fd8; 
        10'b0110011001: data <= 15'h7fbb; 
        10'b0110011010: data <= 15'h7ff4; 
        10'b0110011011: data <= 15'h7fd4; 
        10'b0110011100: data <= 15'h7ff2; 
        10'b0110011101: data <= 15'h7fcd; 
        10'b0110011110: data <= 15'h7fa4; 
        10'b0110011111: data <= 15'h7fbd; 
        10'b0110100000: data <= 15'h7ff3; 
        10'b0110100001: data <= 15'h0021; 
        10'b0110100010: data <= 15'h0025; 
        10'b0110100011: data <= 15'h7feb; 
        10'b0110100100: data <= 15'h7ff2; 
        10'b0110100101: data <= 15'h7ff5; 
        10'b0110100110: data <= 15'h7ff1; 
        10'b0110100111: data <= 15'h001e; 
        10'b0110101000: data <= 15'h000f; 
        10'b0110101001: data <= 15'h0007; 
        10'b0110101010: data <= 15'h0024; 
        10'b0110101011: data <= 15'h002a; 
        10'b0110101100: data <= 15'h004e; 
        10'b0110101101: data <= 15'h0037; 
        10'b0110101110: data <= 15'h0042; 
        10'b0110101111: data <= 15'h0027; 
        10'b0110110000: data <= 15'h0022; 
        10'b0110110001: data <= 15'h0051; 
        10'b0110110010: data <= 15'h0006; 
        10'b0110110011: data <= 15'h0020; 
        10'b0110110100: data <= 15'h0005; 
        10'b0110110101: data <= 15'h7fc0; 
        10'b0110110110: data <= 15'h7fc3; 
        10'b0110110111: data <= 15'h7fdb; 
        10'b0110111000: data <= 15'h7fe5; 
        10'b0110111001: data <= 15'h7fd7; 
        10'b0110111010: data <= 15'h7fad; 
        10'b0110111011: data <= 15'h7fd5; 
        10'b0110111100: data <= 15'h001a; 
        10'b0110111101: data <= 15'h002c; 
        10'b0110111110: data <= 15'h0018; 
        10'b0110111111: data <= 15'h7fe9; 
        10'b0111000000: data <= 15'h7fee; 
        10'b0111000001: data <= 15'h7fe4; 
        10'b0111000010: data <= 15'h7fe1; 
        10'b0111000011: data <= 15'h0020; 
        10'b0111000100: data <= 15'h0044; 
        10'b0111000101: data <= 15'h006f; 
        10'b0111000110: data <= 15'h0071; 
        10'b0111000111: data <= 15'h0043; 
        10'b0111001000: data <= 15'h001c; 
        10'b0111001001: data <= 15'h003a; 
        10'b0111001010: data <= 15'h0036; 
        10'b0111001011: data <= 15'h0031; 
        10'b0111001100: data <= 15'h0065; 
        10'b0111001101: data <= 15'h0059; 
        10'b0111001110: data <= 15'h0013; 
        10'b0111001111: data <= 15'h7ff5; 
        10'b0111010000: data <= 15'h0000; 
        10'b0111010001: data <= 15'h7fd6; 
        10'b0111010010: data <= 15'h7fdc; 
        10'b0111010011: data <= 15'h7fc0; 
        10'b0111010100: data <= 15'h7fe9; 
        10'b0111010101: data <= 15'h0003; 
        10'b0111010110: data <= 15'h000e; 
        10'b0111010111: data <= 15'h001e; 
        10'b0111011000: data <= 15'h005e; 
        10'b0111011001: data <= 15'h0075; 
        10'b0111011010: data <= 15'h0014; 
        10'b0111011011: data <= 15'h7fee; 
        10'b0111011100: data <= 15'h7ff1; 
        10'b0111011101: data <= 15'h0005; 
        10'b0111011110: data <= 15'h7ff4; 
        10'b0111011111: data <= 15'h0027; 
        10'b0111100000: data <= 15'h0074; 
        10'b0111100001: data <= 15'h00a1; 
        10'b0111100010: data <= 15'h0093; 
        10'b0111100011: data <= 15'h0065; 
        10'b0111100100: data <= 15'h0046; 
        10'b0111100101: data <= 15'h0055; 
        10'b0111100110: data <= 15'h0083; 
        10'b0111100111: data <= 15'h006b; 
        10'b0111101000: data <= 15'h007b; 
        10'b0111101001: data <= 15'h003a; 
        10'b0111101010: data <= 15'h001e; 
        10'b0111101011: data <= 15'h0028; 
        10'b0111101100: data <= 15'h0028; 
        10'b0111101101: data <= 15'h7ffa; 
        10'b0111101110: data <= 15'h001a; 
        10'b0111101111: data <= 15'h7fef; 
        10'b0111110000: data <= 15'h0030; 
        10'b0111110001: data <= 15'h0034; 
        10'b0111110010: data <= 15'h0026; 
        10'b0111110011: data <= 15'h0035; 
        10'b0111110100: data <= 15'h0097; 
        10'b0111110101: data <= 15'h0083; 
        10'b0111110110: data <= 15'h001e; 
        10'b0111110111: data <= 15'h0004; 
        10'b0111111000: data <= 15'h7ffd; 
        10'b0111111001: data <= 15'h7ffe; 
        10'b0111111010: data <= 15'h7fd8; 
        10'b0111111011: data <= 15'h000b; 
        10'b0111111100: data <= 15'h007d; 
        10'b0111111101: data <= 15'h00d4; 
        10'b0111111110: data <= 15'h00c7; 
        10'b0111111111: data <= 15'h008f; 
        10'b1000000000: data <= 15'h0060; 
        10'b1000000001: data <= 15'h006a; 
        10'b1000000010: data <= 15'h00a3; 
        10'b1000000011: data <= 15'h0093; 
        10'b1000000100: data <= 15'h00ea; 
        10'b1000000101: data <= 15'h00ab; 
        10'b1000000110: data <= 15'h0095; 
        10'b1000000111: data <= 15'h0049; 
        10'b1000001000: data <= 15'h0032; 
        10'b1000001001: data <= 15'h005c; 
        10'b1000001010: data <= 15'h003b; 
        10'b1000001011: data <= 15'h0028; 
        10'b1000001100: data <= 15'h006c; 
        10'b1000001101: data <= 15'h0070; 
        10'b1000001110: data <= 15'h007a; 
        10'b1000001111: data <= 15'h00a1; 
        10'b1000010000: data <= 15'h00c8; 
        10'b1000010001: data <= 15'h0073; 
        10'b1000010010: data <= 15'h7ff5; 
        10'b1000010011: data <= 15'h7fe8; 
        10'b1000010100: data <= 15'h7fec; 
        10'b1000010101: data <= 15'h7fed; 
        10'b1000010110: data <= 15'h7fe4; 
        10'b1000010111: data <= 15'h0000; 
        10'b1000011000: data <= 15'h0045; 
        10'b1000011001: data <= 15'h0081; 
        10'b1000011010: data <= 15'h00a3; 
        10'b1000011011: data <= 15'h008d; 
        10'b1000011100: data <= 15'h0082; 
        10'b1000011101: data <= 15'h008a; 
        10'b1000011110: data <= 15'h0084; 
        10'b1000011111: data <= 15'h008c; 
        10'b1000100000: data <= 15'h009d; 
        10'b1000100001: data <= 15'h0079; 
        10'b1000100010: data <= 15'h004e; 
        10'b1000100011: data <= 15'h0025; 
        10'b1000100100: data <= 15'h0039; 
        10'b1000100101: data <= 15'h0064; 
        10'b1000100110: data <= 15'h0030; 
        10'b1000100111: data <= 15'h002f; 
        10'b1000101000: data <= 15'h0050; 
        10'b1000101001: data <= 15'h0064; 
        10'b1000101010: data <= 15'h0083; 
        10'b1000101011: data <= 15'h008d; 
        10'b1000101100: data <= 15'h0079; 
        10'b1000101101: data <= 15'h003f; 
        10'b1000101110: data <= 15'h0005; 
        10'b1000101111: data <= 15'h0001; 
        10'b1000110000: data <= 15'h7fe7; 
        10'b1000110001: data <= 15'h7ffe; 
        10'b1000110010: data <= 15'h7ff9; 
        10'b1000110011: data <= 15'h7fdd; 
        10'b1000110100: data <= 15'h003d; 
        10'b1000110101: data <= 15'h004c; 
        10'b1000110110: data <= 15'h0075; 
        10'b1000110111: data <= 15'h00a3; 
        10'b1000111000: data <= 15'h009b; 
        10'b1000111001: data <= 15'h0067; 
        10'b1000111010: data <= 15'h0063; 
        10'b1000111011: data <= 15'h00a5; 
        10'b1000111100: data <= 15'h005c; 
        10'b1000111101: data <= 15'h001e; 
        10'b1000111110: data <= 15'h0014; 
        10'b1000111111: data <= 15'h0019; 
        10'b1001000000: data <= 15'h0020; 
        10'b1001000001: data <= 15'h0001; 
        10'b1001000010: data <= 15'h0047; 
        10'b1001000011: data <= 15'h0070; 
        10'b1001000100: data <= 15'h004c; 
        10'b1001000101: data <= 15'h006c; 
        10'b1001000110: data <= 15'h0096; 
        10'b1001000111: data <= 15'h0082; 
        10'b1001001000: data <= 15'h005e; 
        10'b1001001001: data <= 15'h002c; 
        10'b1001001010: data <= 15'h7fff; 
        10'b1001001011: data <= 15'h7ffc; 
        10'b1001001100: data <= 15'h7ff6; 
        10'b1001001101: data <= 15'h7fe8; 
        10'b1001001110: data <= 15'h7ffc; 
        10'b1001001111: data <= 15'h7ff2; 
        10'b1001010000: data <= 15'h000d; 
        10'b1001010001: data <= 15'h0020; 
        10'b1001010010: data <= 15'h0051; 
        10'b1001010011: data <= 15'h005b; 
        10'b1001010100: data <= 15'h0051; 
        10'b1001010101: data <= 15'h0065; 
        10'b1001010110: data <= 15'h0059; 
        10'b1001010111: data <= 15'h0057; 
        10'b1001011000: data <= 15'h0022; 
        10'b1001011001: data <= 15'h0010; 
        10'b1001011010: data <= 15'h7ff7; 
        10'b1001011011: data <= 15'h0004; 
        10'b1001011100: data <= 15'h002b; 
        10'b1001011101: data <= 15'h0030; 
        10'b1001011110: data <= 15'h0068; 
        10'b1001011111: data <= 15'h006e; 
        10'b1001100000: data <= 15'h0030; 
        10'b1001100001: data <= 15'h006c; 
        10'b1001100010: data <= 15'h0085; 
        10'b1001100011: data <= 15'h0097; 
        10'b1001100100: data <= 15'h004b; 
        10'b1001100101: data <= 15'h001e; 
        10'b1001100110: data <= 15'h0007; 
        10'b1001100111: data <= 15'h7ffd; 
        10'b1001101000: data <= 15'h7fe7; 
        10'b1001101001: data <= 15'h7ff9; 
        10'b1001101010: data <= 15'h7fea; 
        10'b1001101011: data <= 15'h0007; 
        10'b1001101100: data <= 15'h001a; 
        10'b1001101101: data <= 15'h0009; 
        10'b1001101110: data <= 15'h0037; 
        10'b1001101111: data <= 15'h0031; 
        10'b1001110000: data <= 15'h002d; 
        10'b1001110001: data <= 15'h0040; 
        10'b1001110010: data <= 15'h003f; 
        10'b1001110011: data <= 15'h004b; 
        10'b1001110100: data <= 15'h0008; 
        10'b1001110101: data <= 15'h7fc5; 
        10'b1001110110: data <= 15'h7fb6; 
        10'b1001110111: data <= 15'h7fd6; 
        10'b1001111000: data <= 15'h7fd8; 
        10'b1001111001: data <= 15'h001f; 
        10'b1001111010: data <= 15'h0061; 
        10'b1001111011: data <= 15'h007c; 
        10'b1001111100: data <= 15'h0071; 
        10'b1001111101: data <= 15'h006c; 
        10'b1001111110: data <= 15'h005d; 
        10'b1001111111: data <= 15'h0067; 
        10'b1010000000: data <= 15'h0026; 
        10'b1010000001: data <= 15'h7ffc; 
        10'b1010000010: data <= 15'h7ff9; 
        10'b1010000011: data <= 15'h7fee; 
        10'b1010000100: data <= 15'h7ffa; 
        10'b1010000101: data <= 15'h7ffb; 
        10'b1010000110: data <= 15'h7ff5; 
        10'b1010000111: data <= 15'h7ff3; 
        10'b1010001000: data <= 15'h7ff1; 
        10'b1010001001: data <= 15'h7fe3; 
        10'b1010001010: data <= 15'h7fdd; 
        10'b1010001011: data <= 15'h7fe1; 
        10'b1010001100: data <= 15'h7fce; 
        10'b1010001101: data <= 15'h7fe2; 
        10'b1010001110: data <= 15'h7fec; 
        10'b1010001111: data <= 15'h0019; 
        10'b1010010000: data <= 15'h0002; 
        10'b1010010001: data <= 15'h7fd8; 
        10'b1010010010: data <= 15'h7fca; 
        10'b1010010011: data <= 15'h7fba; 
        10'b1010010100: data <= 15'h7fb4; 
        10'b1010010101: data <= 15'h7fd8; 
        10'b1010010110: data <= 15'h0010; 
        10'b1010010111: data <= 15'h0061; 
        10'b1010011000: data <= 15'h0055; 
        10'b1010011001: data <= 15'h0068; 
        10'b1010011010: data <= 15'h004b; 
        10'b1010011011: data <= 15'h001c; 
        10'b1010011100: data <= 15'h0011; 
        10'b1010011101: data <= 15'h000b; 
        10'b1010011110: data <= 15'h7ffe; 
        10'b1010011111: data <= 15'h7ff3; 
        10'b1010100000: data <= 15'h7ff6; 
        10'b1010100001: data <= 15'h7fec; 
        10'b1010100010: data <= 15'h7fff; 
        10'b1010100011: data <= 15'h7ffd; 
        10'b1010100100: data <= 15'h7feb; 
        10'b1010100101: data <= 15'h7fca; 
        10'b1010100110: data <= 15'h7f97; 
        10'b1010100111: data <= 15'h7fb2; 
        10'b1010101000: data <= 15'h7faf; 
        10'b1010101001: data <= 15'h7faa; 
        10'b1010101010: data <= 15'h7fab; 
        10'b1010101011: data <= 15'h7fbf; 
        10'b1010101100: data <= 15'h7fbe; 
        10'b1010101101: data <= 15'h7fdc; 
        10'b1010101110: data <= 15'h7fd1; 
        10'b1010101111: data <= 15'h7fbd; 
        10'b1010110000: data <= 15'h7fc1; 
        10'b1010110001: data <= 15'h7fce; 
        10'b1010110010: data <= 15'h7fc3; 
        10'b1010110011: data <= 15'h7fdf; 
        10'b1010110100: data <= 15'h7fe3; 
        10'b1010110101: data <= 15'h7fe3; 
        10'b1010110110: data <= 15'h7fef; 
        10'b1010110111: data <= 15'h7ff3; 
        10'b1010111000: data <= 15'h7ffe; 
        10'b1010111001: data <= 15'h000b; 
        10'b1010111010: data <= 15'h7fe9; 
        10'b1010111011: data <= 15'h7fea; 
        10'b1010111100: data <= 15'h7fff; 
        10'b1010111101: data <= 15'h7fe4; 
        10'b1010111110: data <= 15'h7ff2; 
        10'b1010111111: data <= 15'h7fef; 
        10'b1011000000: data <= 15'h7fea; 
        10'b1011000001: data <= 15'h7fda; 
        10'b1011000010: data <= 15'h7fcd; 
        10'b1011000011: data <= 15'h7fb3; 
        10'b1011000100: data <= 15'h7faa; 
        10'b1011000101: data <= 15'h7fb0; 
        10'b1011000110: data <= 15'h7fb8; 
        10'b1011000111: data <= 15'h7fa4; 
        10'b1011001000: data <= 15'h7fc2; 
        10'b1011001001: data <= 15'h7fc6; 
        10'b1011001010: data <= 15'h7fb3; 
        10'b1011001011: data <= 15'h7fc1; 
        10'b1011001100: data <= 15'h7fd1; 
        10'b1011001101: data <= 15'h7fd4; 
        10'b1011001110: data <= 15'h7fef; 
        10'b1011001111: data <= 15'h7fd8; 
        10'b1011010000: data <= 15'h7ff2; 
        10'b1011010001: data <= 15'h7ff0; 
        10'b1011010010: data <= 15'h7fff; 
        10'b1011010011: data <= 15'h7fea; 
        10'b1011010100: data <= 15'h7ff8; 
        10'b1011010101: data <= 15'h7feb; 
        10'b1011010110: data <= 15'h7fe4; 
        10'b1011010111: data <= 15'h7feb; 
        10'b1011011000: data <= 15'h7fe5; 
        10'b1011011001: data <= 15'h7fef; 
        10'b1011011010: data <= 15'h7ff4; 
        10'b1011011011: data <= 15'h0001; 
        10'b1011011100: data <= 15'h7ffc; 
        10'b1011011101: data <= 15'h7ff3; 
        10'b1011011110: data <= 15'h7ffb; 
        10'b1011011111: data <= 15'h7fff; 
        10'b1011100000: data <= 15'h7ff2; 
        10'b1011100001: data <= 15'h0002; 
        10'b1011100010: data <= 15'h0000; 
        10'b1011100011: data <= 15'h0001; 
        10'b1011100100: data <= 15'h0003; 
        10'b1011100101: data <= 15'h7ff8; 
        10'b1011100110: data <= 15'h7fee; 
        10'b1011100111: data <= 15'h7fe2; 
        10'b1011101000: data <= 15'h7ff0; 
        10'b1011101001: data <= 15'h7ff8; 
        10'b1011101010: data <= 15'h7ff6; 
        10'b1011101011: data <= 15'h7feb; 
        10'b1011101100: data <= 15'h0003; 
        10'b1011101101: data <= 15'h7fff; 
        10'b1011101110: data <= 15'h7feb; 
        10'b1011101111: data <= 15'h7fef; 
        10'b1011110000: data <= 15'h7fe5; 
        10'b1011110001: data <= 15'h0001; 
        10'b1011110010: data <= 15'h0001; 
        10'b1011110011: data <= 15'h7fff; 
        10'b1011110100: data <= 15'h7ffe; 
        10'b1011110101: data <= 15'h7fec; 
        10'b1011110110: data <= 15'h7fe8; 
        10'b1011110111: data <= 15'h7ff6; 
        10'b1011111000: data <= 15'h7fe5; 
        10'b1011111001: data <= 15'h0006; 
        10'b1011111010: data <= 15'h0005; 
        10'b1011111011: data <= 15'h7ff0; 
        10'b1011111100: data <= 15'h7ffe; 
        10'b1011111101: data <= 15'h7feb; 
        10'b1011111110: data <= 15'h0004; 
        10'b1011111111: data <= 15'h7fe4; 
        10'b1100000000: data <= 15'h7fff; 
        10'b1100000001: data <= 15'h7ff2; 
        10'b1100000010: data <= 15'h7ffa; 
        10'b1100000011: data <= 15'h7fe8; 
        10'b1100000100: data <= 15'h7ff6; 
        10'b1100000101: data <= 15'h7ff1; 
        10'b1100000110: data <= 15'h7ff8; 
        10'b1100000111: data <= 15'h7ff6; 
        10'b1100001000: data <= 15'h7ffd; 
        10'b1100001001: data <= 15'h7fe3; 
        10'b1100001010: data <= 15'h7ff4; 
        10'b1100001011: data <= 15'h0001; 
        10'b1100001100: data <= 15'h7fe3; 
        10'b1100001101: data <= 15'h7ff5; 
        10'b1100001110: data <= 15'h7ffc; 
        10'b1100001111: data <= 15'h7ff0; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 10) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 16'hffcd; 
        10'b0000000001: data <= 16'h0001; 
        10'b0000000010: data <= 16'hffe6; 
        10'b0000000011: data <= 16'hffd6; 
        10'b0000000100: data <= 16'hffe6; 
        10'b0000000101: data <= 16'hffd8; 
        10'b0000000110: data <= 16'hffef; 
        10'b0000000111: data <= 16'hfff1; 
        10'b0000001000: data <= 16'hffcb; 
        10'b0000001001: data <= 16'hffeb; 
        10'b0000001010: data <= 16'hffcf; 
        10'b0000001011: data <= 16'hffdf; 
        10'b0000001100: data <= 16'h000a; 
        10'b0000001101: data <= 16'h0009; 
        10'b0000001110: data <= 16'hffce; 
        10'b0000001111: data <= 16'hffee; 
        10'b0000010000: data <= 16'hffd1; 
        10'b0000010001: data <= 16'hffd2; 
        10'b0000010010: data <= 16'h000d; 
        10'b0000010011: data <= 16'h0004; 
        10'b0000010100: data <= 16'hffda; 
        10'b0000010101: data <= 16'hfff0; 
        10'b0000010110: data <= 16'hffde; 
        10'b0000010111: data <= 16'hffc8; 
        10'b0000011000: data <= 16'hffcd; 
        10'b0000011001: data <= 16'hffed; 
        10'b0000011010: data <= 16'hfffd; 
        10'b0000011011: data <= 16'hfff2; 
        10'b0000011100: data <= 16'hffea; 
        10'b0000011101: data <= 16'hffe7; 
        10'b0000011110: data <= 16'h000c; 
        10'b0000011111: data <= 16'hfff3; 
        10'b0000100000: data <= 16'hffcf; 
        10'b0000100001: data <= 16'hffce; 
        10'b0000100010: data <= 16'hffcc; 
        10'b0000100011: data <= 16'hffd8; 
        10'b0000100100: data <= 16'hffd9; 
        10'b0000100101: data <= 16'hffee; 
        10'b0000100110: data <= 16'h0001; 
        10'b0000100111: data <= 16'hffd1; 
        10'b0000101000: data <= 16'hffe2; 
        10'b0000101001: data <= 16'hffcf; 
        10'b0000101010: data <= 16'hffef; 
        10'b0000101011: data <= 16'hffc8; 
        10'b0000101100: data <= 16'hfff1; 
        10'b0000101101: data <= 16'hffd1; 
        10'b0000101110: data <= 16'hffe0; 
        10'b0000101111: data <= 16'hffd5; 
        10'b0000110000: data <= 16'hffee; 
        10'b0000110001: data <= 16'hffd2; 
        10'b0000110010: data <= 16'hffca; 
        10'b0000110011: data <= 16'hffc5; 
        10'b0000110100: data <= 16'h0003; 
        10'b0000110101: data <= 16'hfff3; 
        10'b0000110110: data <= 16'h0004; 
        10'b0000110111: data <= 16'hffdd; 
        10'b0000111000: data <= 16'hffe7; 
        10'b0000111001: data <= 16'hffc9; 
        10'b0000111010: data <= 16'hffce; 
        10'b0000111011: data <= 16'h0000; 
        10'b0000111100: data <= 16'hffcb; 
        10'b0000111101: data <= 16'hffcf; 
        10'b0000111110: data <= 16'hffe4; 
        10'b0000111111: data <= 16'hffed; 
        10'b0001000000: data <= 16'hfffb; 
        10'b0001000001: data <= 16'hffe2; 
        10'b0001000010: data <= 16'h001d; 
        10'b0001000011: data <= 16'h0018; 
        10'b0001000100: data <= 16'h004a; 
        10'b0001000101: data <= 16'h003b; 
        10'b0001000110: data <= 16'h0036; 
        10'b0001000111: data <= 16'h0015; 
        10'b0001001000: data <= 16'h0049; 
        10'b0001001001: data <= 16'h0019; 
        10'b0001001010: data <= 16'h0015; 
        10'b0001001011: data <= 16'hffdb; 
        10'b0001001100: data <= 16'hffff; 
        10'b0001001101: data <= 16'hffef; 
        10'b0001001110: data <= 16'hffb5; 
        10'b0001001111: data <= 16'hffe6; 
        10'b0001010000: data <= 16'hfff8; 
        10'b0001010001: data <= 16'h0012; 
        10'b0001010010: data <= 16'hffea; 
        10'b0001010011: data <= 16'hffe2; 
        10'b0001010100: data <= 16'hffdb; 
        10'b0001010101: data <= 16'hffd6; 
        10'b0001010110: data <= 16'hfff4; 
        10'b0001010111: data <= 16'hffda; 
        10'b0001011000: data <= 16'h000a; 
        10'b0001011001: data <= 16'hffd2; 
        10'b0001011010: data <= 16'hffef; 
        10'b0001011011: data <= 16'h0000; 
        10'b0001011100: data <= 16'h000d; 
        10'b0001011101: data <= 16'h0076; 
        10'b0001011110: data <= 16'h00b8; 
        10'b0001011111: data <= 16'h00b7; 
        10'b0001100000: data <= 16'h00af; 
        10'b0001100001: data <= 16'h0102; 
        10'b0001100010: data <= 16'h008d; 
        10'b0001100011: data <= 16'h003e; 
        10'b0001100100: data <= 16'h0076; 
        10'b0001100101: data <= 16'h0036; 
        10'b0001100110: data <= 16'hffcd; 
        10'b0001100111: data <= 16'hfff3; 
        10'b0001101000: data <= 16'hffc6; 
        10'b0001101001: data <= 16'hffbc; 
        10'b0001101010: data <= 16'hffad; 
        10'b0001101011: data <= 16'hffd7; 
        10'b0001101100: data <= 16'h0006; 
        10'b0001101101: data <= 16'h0014; 
        10'b0001101110: data <= 16'hffd2; 
        10'b0001101111: data <= 16'hfff7; 
        10'b0001110000: data <= 16'hffd8; 
        10'b0001110001: data <= 16'hffe4; 
        10'b0001110010: data <= 16'h000e; 
        10'b0001110011: data <= 16'hffc4; 
        10'b0001110100: data <= 16'hffcb; 
        10'b0001110101: data <= 16'hffef; 
        10'b0001110110: data <= 16'h001b; 
        10'b0001110111: data <= 16'h001a; 
        10'b0001111000: data <= 16'h004c; 
        10'b0001111001: data <= 16'h00e2; 
        10'b0001111010: data <= 16'h00e4; 
        10'b0001111011: data <= 16'h011e; 
        10'b0001111100: data <= 16'h00f2; 
        10'b0001111101: data <= 16'h00c0; 
        10'b0001111110: data <= 16'h00ae; 
        10'b0001111111: data <= 16'h004d; 
        10'b0010000000: data <= 16'h0067; 
        10'b0010000001: data <= 16'h005f; 
        10'b0010000010: data <= 16'hffe3; 
        10'b0010000011: data <= 16'hffd0; 
        10'b0010000100: data <= 16'hffdb; 
        10'b0010000101: data <= 16'hff8f; 
        10'b0010000110: data <= 16'hff77; 
        10'b0010000111: data <= 16'hff7c; 
        10'b0010001000: data <= 16'hffef; 
        10'b0010001001: data <= 16'hffef; 
        10'b0010001010: data <= 16'hffc9; 
        10'b0010001011: data <= 16'hfff6; 
        10'b0010001100: data <= 16'h0005; 
        10'b0010001101: data <= 16'hffee; 
        10'b0010001110: data <= 16'hffd5; 
        10'b0010001111: data <= 16'hffc6; 
        10'b0010010000: data <= 16'hffd0; 
        10'b0010010001: data <= 16'hffd7; 
        10'b0010010010: data <= 16'h0019; 
        10'b0010010011: data <= 16'h006e; 
        10'b0010010100: data <= 16'h0099; 
        10'b0010010101: data <= 16'h0106; 
        10'b0010010110: data <= 16'h0122; 
        10'b0010010111: data <= 16'h012e; 
        10'b0010011000: data <= 16'h0115; 
        10'b0010011001: data <= 16'h0137; 
        10'b0010011010: data <= 16'h011f; 
        10'b0010011011: data <= 16'h010b; 
        10'b0010011100: data <= 16'h0121; 
        10'b0010011101: data <= 16'h00ea; 
        10'b0010011110: data <= 16'h00a9; 
        10'b0010011111: data <= 16'hffb9; 
        10'b0010100000: data <= 16'hffbb; 
        10'b0010100001: data <= 16'hff8f; 
        10'b0010100010: data <= 16'hff8e; 
        10'b0010100011: data <= 16'hff4e; 
        10'b0010100100: data <= 16'hffb3; 
        10'b0010100101: data <= 16'hffd4; 
        10'b0010100110: data <= 16'h0007; 
        10'b0010100111: data <= 16'hffde; 
        10'b0010101000: data <= 16'hffe9; 
        10'b0010101001: data <= 16'hffd7; 
        10'b0010101010: data <= 16'h0009; 
        10'b0010101011: data <= 16'hffea; 
        10'b0010101100: data <= 16'hffe3; 
        10'b0010101101: data <= 16'h0012; 
        10'b0010101110: data <= 16'h006c; 
        10'b0010101111: data <= 16'h00d1; 
        10'b0010110000: data <= 16'h00a0; 
        10'b0010110001: data <= 16'h00b5; 
        10'b0010110010: data <= 16'h00f5; 
        10'b0010110011: data <= 16'h0099; 
        10'b0010110100: data <= 16'h00a3; 
        10'b0010110101: data <= 16'h00d2; 
        10'b0010110110: data <= 16'h00ba; 
        10'b0010110111: data <= 16'h0065; 
        10'b0010111000: data <= 16'h0070; 
        10'b0010111001: data <= 16'h001d; 
        10'b0010111010: data <= 16'h0015; 
        10'b0010111011: data <= 16'hffbe; 
        10'b0010111100: data <= 16'hffd4; 
        10'b0010111101: data <= 16'hff71; 
        10'b0010111110: data <= 16'hff72; 
        10'b0010111111: data <= 16'hff3a; 
        10'b0011000000: data <= 16'hff8a; 
        10'b0011000001: data <= 16'hffbe; 
        10'b0011000010: data <= 16'h0008; 
        10'b0011000011: data <= 16'hfff9; 
        10'b0011000100: data <= 16'hffe1; 
        10'b0011000101: data <= 16'h0006; 
        10'b0011000110: data <= 16'h0007; 
        10'b0011000111: data <= 16'hffe4; 
        10'b0011001000: data <= 16'h0003; 
        10'b0011001001: data <= 16'h003a; 
        10'b0011001010: data <= 16'h008b; 
        10'b0011001011: data <= 16'h00c9; 
        10'b0011001100: data <= 16'h00a5; 
        10'b0011001101: data <= 16'h009a; 
        10'b0011001110: data <= 16'h003b; 
        10'b0011001111: data <= 16'h0045; 
        10'b0011010000: data <= 16'h000c; 
        10'b0011010001: data <= 16'h006c; 
        10'b0011010010: data <= 16'h0085; 
        10'b0011010011: data <= 16'h001c; 
        10'b0011010100: data <= 16'h0012; 
        10'b0011010101: data <= 16'hff58; 
        10'b0011010110: data <= 16'hffc7; 
        10'b0011010111: data <= 16'hffd1; 
        10'b0011011000: data <= 16'hffca; 
        10'b0011011001: data <= 16'hffc1; 
        10'b0011011010: data <= 16'hffd1; 
        10'b0011011011: data <= 16'hff5d; 
        10'b0011011100: data <= 16'hff8f; 
        10'b0011011101: data <= 16'hffdd; 
        10'b0011011110: data <= 16'hffd4; 
        10'b0011011111: data <= 16'hffcb; 
        10'b0011100000: data <= 16'hfff4; 
        10'b0011100001: data <= 16'h0008; 
        10'b0011100010: data <= 16'hffe9; 
        10'b0011100011: data <= 16'h0007; 
        10'b0011100100: data <= 16'h001e; 
        10'b0011100101: data <= 16'h005e; 
        10'b0011100110: data <= 16'h0044; 
        10'b0011100111: data <= 16'h0060; 
        10'b0011101000: data <= 16'h0061; 
        10'b0011101001: data <= 16'h006c; 
        10'b0011101010: data <= 16'h006d; 
        10'b0011101011: data <= 16'h007c; 
        10'b0011101100: data <= 16'h004a; 
        10'b0011101101: data <= 16'h0058; 
        10'b0011101110: data <= 16'h00e8; 
        10'b0011101111: data <= 16'h0083; 
        10'b0011110000: data <= 16'hfff0; 
        10'b0011110001: data <= 16'hffc0; 
        10'b0011110010: data <= 16'hfffe; 
        10'b0011110011: data <= 16'h0034; 
        10'b0011110100: data <= 16'h0001; 
        10'b0011110101: data <= 16'hffdc; 
        10'b0011110110: data <= 16'hffa1; 
        10'b0011110111: data <= 16'hff41; 
        10'b0011111000: data <= 16'hff6e; 
        10'b0011111001: data <= 16'hffc3; 
        10'b0011111010: data <= 16'hffe3; 
        10'b0011111011: data <= 16'hffd1; 
        10'b0011111100: data <= 16'hffd8; 
        10'b0011111101: data <= 16'hfff6; 
        10'b0011111110: data <= 16'hfffe; 
        10'b0011111111: data <= 16'h0018; 
        10'b0100000000: data <= 16'h002f; 
        10'b0100000001: data <= 16'h0069; 
        10'b0100000010: data <= 16'h0025; 
        10'b0100000011: data <= 16'h0007; 
        10'b0100000100: data <= 16'hffdc; 
        10'b0100000101: data <= 16'h0039; 
        10'b0100000110: data <= 16'h002c; 
        10'b0100000111: data <= 16'h0039; 
        10'b0100001000: data <= 16'h000f; 
        10'b0100001001: data <= 16'hfffa; 
        10'b0100001010: data <= 16'h0098; 
        10'b0100001011: data <= 16'h00a4; 
        10'b0100001100: data <= 16'h0039; 
        10'b0100001101: data <= 16'h0004; 
        10'b0100001110: data <= 16'hfff1; 
        10'b0100001111: data <= 16'hffff; 
        10'b0100010000: data <= 16'hfff9; 
        10'b0100010001: data <= 16'hfffc; 
        10'b0100010010: data <= 16'hffc4; 
        10'b0100010011: data <= 16'hff5e; 
        10'b0100010100: data <= 16'hff76; 
        10'b0100010101: data <= 16'hffd3; 
        10'b0100010110: data <= 16'h0007; 
        10'b0100010111: data <= 16'hffcc; 
        10'b0100011000: data <= 16'h000a; 
        10'b0100011001: data <= 16'hfff4; 
        10'b0100011010: data <= 16'hffe8; 
        10'b0100011011: data <= 16'hffde; 
        10'b0100011100: data <= 16'h0007; 
        10'b0100011101: data <= 16'hffe6; 
        10'b0100011110: data <= 16'hffcb; 
        10'b0100011111: data <= 16'hff00; 
        10'b0100100000: data <= 16'hff1b; 
        10'b0100100001: data <= 16'hff53; 
        10'b0100100010: data <= 16'hfef8; 
        10'b0100100011: data <= 16'hfedb; 
        10'b0100100100: data <= 16'hfeab; 
        10'b0100100101: data <= 16'hfe81; 
        10'b0100100110: data <= 16'hff5f; 
        10'b0100100111: data <= 16'h001d; 
        10'b0100101000: data <= 16'h0029; 
        10'b0100101001: data <= 16'h0007; 
        10'b0100101010: data <= 16'h0015; 
        10'b0100101011: data <= 16'hffe1; 
        10'b0100101100: data <= 16'hffe9; 
        10'b0100101101: data <= 16'hffe1; 
        10'b0100101110: data <= 16'hffb0; 
        10'b0100101111: data <= 16'hff46; 
        10'b0100110000: data <= 16'hff9a; 
        10'b0100110001: data <= 16'hfffc; 
        10'b0100110010: data <= 16'hfffb; 
        10'b0100110011: data <= 16'hffd5; 
        10'b0100110100: data <= 16'hffcb; 
        10'b0100110101: data <= 16'h000d; 
        10'b0100110110: data <= 16'hfffb; 
        10'b0100110111: data <= 16'hffcf; 
        10'b0100111000: data <= 16'hffa0; 
        10'b0100111001: data <= 16'hff2e; 
        10'b0100111010: data <= 16'hfe98; 
        10'b0100111011: data <= 16'hfe05; 
        10'b0100111100: data <= 16'hfe19; 
        10'b0100111101: data <= 16'hfdc2; 
        10'b0100111110: data <= 16'hfdc1; 
        10'b0100111111: data <= 16'hfdf3; 
        10'b0101000000: data <= 16'hfdd3; 
        10'b0101000001: data <= 16'hfd59; 
        10'b0101000010: data <= 16'hfdf6; 
        10'b0101000011: data <= 16'hff06; 
        10'b0101000100: data <= 16'hffa9; 
        10'b0101000101: data <= 16'hffb6; 
        10'b0101000110: data <= 16'hffb8; 
        10'b0101000111: data <= 16'hfff2; 
        10'b0101001000: data <= 16'hffd5; 
        10'b0101001001: data <= 16'hffd3; 
        10'b0101001010: data <= 16'hff89; 
        10'b0101001011: data <= 16'hffaf; 
        10'b0101001100: data <= 16'hfff1; 
        10'b0101001101: data <= 16'hffe4; 
        10'b0101001110: data <= 16'hffd4; 
        10'b0101001111: data <= 16'hfff4; 
        10'b0101010000: data <= 16'hffee; 
        10'b0101010001: data <= 16'hfff1; 
        10'b0101010010: data <= 16'h0005; 
        10'b0101010011: data <= 16'hffea; 
        10'b0101010100: data <= 16'hff99; 
        10'b0101010101: data <= 16'hfec8; 
        10'b0101010110: data <= 16'hfda1; 
        10'b0101010111: data <= 16'hfd19; 
        10'b0101011000: data <= 16'hfd4b; 
        10'b0101011001: data <= 16'hfd70; 
        10'b0101011010: data <= 16'hfda8; 
        10'b0101011011: data <= 16'hfdcf; 
        10'b0101011100: data <= 16'hfdd0; 
        10'b0101011101: data <= 16'hfdba; 
        10'b0101011110: data <= 16'hfe22; 
        10'b0101011111: data <= 16'hfec1; 
        10'b0101100000: data <= 16'hff25; 
        10'b0101100001: data <= 16'hff3b; 
        10'b0101100010: data <= 16'hff9d; 
        10'b0101100011: data <= 16'h0000; 
        10'b0101100100: data <= 16'hfffe; 
        10'b0101100101: data <= 16'hffc8; 
        10'b0101100110: data <= 16'hff82; 
        10'b0101100111: data <= 16'hff40; 
        10'b0101101000: data <= 16'hffe9; 
        10'b0101101001: data <= 16'hffe0; 
        10'b0101101010: data <= 16'h000e; 
        10'b0101101011: data <= 16'hfff1; 
        10'b0101101100: data <= 16'hffd9; 
        10'b0101101101: data <= 16'hffe7; 
        10'b0101101110: data <= 16'h000d; 
        10'b0101101111: data <= 16'hffd8; 
        10'b0101110000: data <= 16'hff59; 
        10'b0101110001: data <= 16'hfe77; 
        10'b0101110010: data <= 16'hfd90; 
        10'b0101110011: data <= 16'hfdc3; 
        10'b0101110100: data <= 16'hfde9; 
        10'b0101110101: data <= 16'hfe90; 
        10'b0101110110: data <= 16'hfefb; 
        10'b0101110111: data <= 16'hff86; 
        10'b0101111000: data <= 16'hff3f; 
        10'b0101111001: data <= 16'hffa8; 
        10'b0101111010: data <= 16'hff24; 
        10'b0101111011: data <= 16'hff1f; 
        10'b0101111100: data <= 16'hfef5; 
        10'b0101111101: data <= 16'hff3f; 
        10'b0101111110: data <= 16'hff96; 
        10'b0101111111: data <= 16'hffec; 
        10'b0110000000: data <= 16'hffe1; 
        10'b0110000001: data <= 16'hffbc; 
        10'b0110000010: data <= 16'hff61; 
        10'b0110000011: data <= 16'hff6f; 
        10'b0110000100: data <= 16'hffb7; 
        10'b0110000101: data <= 16'h0012; 
        10'b0110000110: data <= 16'hffe8; 
        10'b0110000111: data <= 16'hfffe; 
        10'b0110001000: data <= 16'h0008; 
        10'b0110001001: data <= 16'hfff3; 
        10'b0110001010: data <= 16'h0001; 
        10'b0110001011: data <= 16'hffde; 
        10'b0110001100: data <= 16'hffc0; 
        10'b0110001101: data <= 16'hfef6; 
        10'b0110001110: data <= 16'hfeb0; 
        10'b0110001111: data <= 16'hfeee; 
        10'b0110010000: data <= 16'hff92; 
        10'b0110010001: data <= 16'hffed; 
        10'b0110010010: data <= 16'h0045; 
        10'b0110010011: data <= 16'h005b; 
        10'b0110010100: data <= 16'h006c; 
        10'b0110010101: data <= 16'h00a7; 
        10'b0110010110: data <= 16'h000b; 
        10'b0110010111: data <= 16'hff95; 
        10'b0110011000: data <= 16'hffb0; 
        10'b0110011001: data <= 16'hff76; 
        10'b0110011010: data <= 16'hffe9; 
        10'b0110011011: data <= 16'hffa7; 
        10'b0110011100: data <= 16'hffe4; 
        10'b0110011101: data <= 16'hff9a; 
        10'b0110011110: data <= 16'hff48; 
        10'b0110011111: data <= 16'hff7a; 
        10'b0110100000: data <= 16'hffe6; 
        10'b0110100001: data <= 16'h0041; 
        10'b0110100010: data <= 16'h004a; 
        10'b0110100011: data <= 16'hffd7; 
        10'b0110100100: data <= 16'hffe3; 
        10'b0110100101: data <= 16'hffe9; 
        10'b0110100110: data <= 16'hffe2; 
        10'b0110100111: data <= 16'h003d; 
        10'b0110101000: data <= 16'h001d; 
        10'b0110101001: data <= 16'h000d; 
        10'b0110101010: data <= 16'h0048; 
        10'b0110101011: data <= 16'h0054; 
        10'b0110101100: data <= 16'h009c; 
        10'b0110101101: data <= 16'h006f; 
        10'b0110101110: data <= 16'h0085; 
        10'b0110101111: data <= 16'h004e; 
        10'b0110110000: data <= 16'h0045; 
        10'b0110110001: data <= 16'h00a2; 
        10'b0110110010: data <= 16'h000c; 
        10'b0110110011: data <= 16'h003f; 
        10'b0110110100: data <= 16'h0009; 
        10'b0110110101: data <= 16'hff80; 
        10'b0110110110: data <= 16'hff86; 
        10'b0110110111: data <= 16'hffb5; 
        10'b0110111000: data <= 16'hffc9; 
        10'b0110111001: data <= 16'hffad; 
        10'b0110111010: data <= 16'hff59; 
        10'b0110111011: data <= 16'hffaa; 
        10'b0110111100: data <= 16'h0033; 
        10'b0110111101: data <= 16'h0057; 
        10'b0110111110: data <= 16'h002f; 
        10'b0110111111: data <= 16'hffd1; 
        10'b0111000000: data <= 16'hffdc; 
        10'b0111000001: data <= 16'hffc9; 
        10'b0111000010: data <= 16'hffc1; 
        10'b0111000011: data <= 16'h0041; 
        10'b0111000100: data <= 16'h0088; 
        10'b0111000101: data <= 16'h00dd; 
        10'b0111000110: data <= 16'h00e1; 
        10'b0111000111: data <= 16'h0086; 
        10'b0111001000: data <= 16'h0038; 
        10'b0111001001: data <= 16'h0074; 
        10'b0111001010: data <= 16'h006b; 
        10'b0111001011: data <= 16'h0062; 
        10'b0111001100: data <= 16'h00ca; 
        10'b0111001101: data <= 16'h00b2; 
        10'b0111001110: data <= 16'h0025; 
        10'b0111001111: data <= 16'hffeb; 
        10'b0111010000: data <= 16'hffff; 
        10'b0111010001: data <= 16'hffad; 
        10'b0111010010: data <= 16'hffb7; 
        10'b0111010011: data <= 16'hff80; 
        10'b0111010100: data <= 16'hffd3; 
        10'b0111010101: data <= 16'h0007; 
        10'b0111010110: data <= 16'h001c; 
        10'b0111010111: data <= 16'h003b; 
        10'b0111011000: data <= 16'h00bd; 
        10'b0111011001: data <= 16'h00ea; 
        10'b0111011010: data <= 16'h0027; 
        10'b0111011011: data <= 16'hffdb; 
        10'b0111011100: data <= 16'hffe2; 
        10'b0111011101: data <= 16'h000b; 
        10'b0111011110: data <= 16'hffe8; 
        10'b0111011111: data <= 16'h004e; 
        10'b0111100000: data <= 16'h00e7; 
        10'b0111100001: data <= 16'h0142; 
        10'b0111100010: data <= 16'h0127; 
        10'b0111100011: data <= 16'h00ca; 
        10'b0111100100: data <= 16'h008c; 
        10'b0111100101: data <= 16'h00aa; 
        10'b0111100110: data <= 16'h0106; 
        10'b0111100111: data <= 16'h00d7; 
        10'b0111101000: data <= 16'h00f6; 
        10'b0111101001: data <= 16'h0073; 
        10'b0111101010: data <= 16'h003b; 
        10'b0111101011: data <= 16'h0050; 
        10'b0111101100: data <= 16'h0051; 
        10'b0111101101: data <= 16'hfff4; 
        10'b0111101110: data <= 16'h0034; 
        10'b0111101111: data <= 16'hffdf; 
        10'b0111110000: data <= 16'h0061; 
        10'b0111110001: data <= 16'h0067; 
        10'b0111110010: data <= 16'h004d; 
        10'b0111110011: data <= 16'h006a; 
        10'b0111110100: data <= 16'h012e; 
        10'b0111110101: data <= 16'h0106; 
        10'b0111110110: data <= 16'h003c; 
        10'b0111110111: data <= 16'h0008; 
        10'b0111111000: data <= 16'hfff9; 
        10'b0111111001: data <= 16'hfffc; 
        10'b0111111010: data <= 16'hffb0; 
        10'b0111111011: data <= 16'h0015; 
        10'b0111111100: data <= 16'h00fb; 
        10'b0111111101: data <= 16'h01a8; 
        10'b0111111110: data <= 16'h018f; 
        10'b0111111111: data <= 16'h011f; 
        10'b1000000000: data <= 16'h00bf; 
        10'b1000000001: data <= 16'h00d5; 
        10'b1000000010: data <= 16'h0145; 
        10'b1000000011: data <= 16'h0126; 
        10'b1000000100: data <= 16'h01d4; 
        10'b1000000101: data <= 16'h0156; 
        10'b1000000110: data <= 16'h012a; 
        10'b1000000111: data <= 16'h0091; 
        10'b1000001000: data <= 16'h0064; 
        10'b1000001001: data <= 16'h00b8; 
        10'b1000001010: data <= 16'h0076; 
        10'b1000001011: data <= 16'h0051; 
        10'b1000001100: data <= 16'h00d9; 
        10'b1000001101: data <= 16'h00e0; 
        10'b1000001110: data <= 16'h00f4; 
        10'b1000001111: data <= 16'h0142; 
        10'b1000010000: data <= 16'h0190; 
        10'b1000010001: data <= 16'h00e7; 
        10'b1000010010: data <= 16'hffea; 
        10'b1000010011: data <= 16'hffd0; 
        10'b1000010100: data <= 16'hffd8; 
        10'b1000010101: data <= 16'hffda; 
        10'b1000010110: data <= 16'hffc8; 
        10'b1000010111: data <= 16'hffff; 
        10'b1000011000: data <= 16'h008a; 
        10'b1000011001: data <= 16'h0101; 
        10'b1000011010: data <= 16'h0145; 
        10'b1000011011: data <= 16'h011a; 
        10'b1000011100: data <= 16'h0104; 
        10'b1000011101: data <= 16'h0113; 
        10'b1000011110: data <= 16'h0108; 
        10'b1000011111: data <= 16'h0118; 
        10'b1000100000: data <= 16'h0139; 
        10'b1000100001: data <= 16'h00f1; 
        10'b1000100010: data <= 16'h009c; 
        10'b1000100011: data <= 16'h004a; 
        10'b1000100100: data <= 16'h0073; 
        10'b1000100101: data <= 16'h00c8; 
        10'b1000100110: data <= 16'h0060; 
        10'b1000100111: data <= 16'h005e; 
        10'b1000101000: data <= 16'h00a1; 
        10'b1000101001: data <= 16'h00c9; 
        10'b1000101010: data <= 16'h0106; 
        10'b1000101011: data <= 16'h0119; 
        10'b1000101100: data <= 16'h00f2; 
        10'b1000101101: data <= 16'h007f; 
        10'b1000101110: data <= 16'h000b; 
        10'b1000101111: data <= 16'h0003; 
        10'b1000110000: data <= 16'hffce; 
        10'b1000110001: data <= 16'hfffc; 
        10'b1000110010: data <= 16'hfff3; 
        10'b1000110011: data <= 16'hffbb; 
        10'b1000110100: data <= 16'h007a; 
        10'b1000110101: data <= 16'h0097; 
        10'b1000110110: data <= 16'h00ea; 
        10'b1000110111: data <= 16'h0146; 
        10'b1000111000: data <= 16'h0136; 
        10'b1000111001: data <= 16'h00cd; 
        10'b1000111010: data <= 16'h00c5; 
        10'b1000111011: data <= 16'h014a; 
        10'b1000111100: data <= 16'h00b8; 
        10'b1000111101: data <= 16'h003d; 
        10'b1000111110: data <= 16'h0029; 
        10'b1000111111: data <= 16'h0032; 
        10'b1001000000: data <= 16'h0041; 
        10'b1001000001: data <= 16'h0003; 
        10'b1001000010: data <= 16'h008f; 
        10'b1001000011: data <= 16'h00df; 
        10'b1001000100: data <= 16'h0097; 
        10'b1001000101: data <= 16'h00d7; 
        10'b1001000110: data <= 16'h012c; 
        10'b1001000111: data <= 16'h0104; 
        10'b1001001000: data <= 16'h00bb; 
        10'b1001001001: data <= 16'h0059; 
        10'b1001001010: data <= 16'hffff; 
        10'b1001001011: data <= 16'hfff8; 
        10'b1001001100: data <= 16'hffec; 
        10'b1001001101: data <= 16'hffd0; 
        10'b1001001110: data <= 16'hfff7; 
        10'b1001001111: data <= 16'hffe4; 
        10'b1001010000: data <= 16'h001a; 
        10'b1001010001: data <= 16'h0041; 
        10'b1001010010: data <= 16'h00a3; 
        10'b1001010011: data <= 16'h00b7; 
        10'b1001010100: data <= 16'h00a1; 
        10'b1001010101: data <= 16'h00c9; 
        10'b1001010110: data <= 16'h00b2; 
        10'b1001010111: data <= 16'h00af; 
        10'b1001011000: data <= 16'h0045; 
        10'b1001011001: data <= 16'h0021; 
        10'b1001011010: data <= 16'hffee; 
        10'b1001011011: data <= 16'h0008; 
        10'b1001011100: data <= 16'h0057; 
        10'b1001011101: data <= 16'h005f; 
        10'b1001011110: data <= 16'h00d1; 
        10'b1001011111: data <= 16'h00db; 
        10'b1001100000: data <= 16'h0060; 
        10'b1001100001: data <= 16'h00d7; 
        10'b1001100010: data <= 16'h010a; 
        10'b1001100011: data <= 16'h012f; 
        10'b1001100100: data <= 16'h0095; 
        10'b1001100101: data <= 16'h003b; 
        10'b1001100110: data <= 16'h000e; 
        10'b1001100111: data <= 16'hfff9; 
        10'b1001101000: data <= 16'hffcd; 
        10'b1001101001: data <= 16'hfff2; 
        10'b1001101010: data <= 16'hffd4; 
        10'b1001101011: data <= 16'h000e; 
        10'b1001101100: data <= 16'h0033; 
        10'b1001101101: data <= 16'h0012; 
        10'b1001101110: data <= 16'h006f; 
        10'b1001101111: data <= 16'h0061; 
        10'b1001110000: data <= 16'h005b; 
        10'b1001110001: data <= 16'h007f; 
        10'b1001110010: data <= 16'h007e; 
        10'b1001110011: data <= 16'h0096; 
        10'b1001110100: data <= 16'h0010; 
        10'b1001110101: data <= 16'hff8a; 
        10'b1001110110: data <= 16'hff6b; 
        10'b1001110111: data <= 16'hffac; 
        10'b1001111000: data <= 16'hffb1; 
        10'b1001111001: data <= 16'h003e; 
        10'b1001111010: data <= 16'h00c2; 
        10'b1001111011: data <= 16'h00f7; 
        10'b1001111100: data <= 16'h00e1; 
        10'b1001111101: data <= 16'h00d7; 
        10'b1001111110: data <= 16'h00bb; 
        10'b1001111111: data <= 16'h00ce; 
        10'b1010000000: data <= 16'h004d; 
        10'b1010000001: data <= 16'hfff8; 
        10'b1010000010: data <= 16'hfff3; 
        10'b1010000011: data <= 16'hffdc; 
        10'b1010000100: data <= 16'hfff4; 
        10'b1010000101: data <= 16'hfff5; 
        10'b1010000110: data <= 16'hffea; 
        10'b1010000111: data <= 16'hffe6; 
        10'b1010001000: data <= 16'hffe3; 
        10'b1010001001: data <= 16'hffc6; 
        10'b1010001010: data <= 16'hffb9; 
        10'b1010001011: data <= 16'hffc3; 
        10'b1010001100: data <= 16'hff9b; 
        10'b1010001101: data <= 16'hffc5; 
        10'b1010001110: data <= 16'hffd9; 
        10'b1010001111: data <= 16'h0033; 
        10'b1010010000: data <= 16'h0005; 
        10'b1010010001: data <= 16'hffb1; 
        10'b1010010010: data <= 16'hff95; 
        10'b1010010011: data <= 16'hff74; 
        10'b1010010100: data <= 16'hff68; 
        10'b1010010101: data <= 16'hffb1; 
        10'b1010010110: data <= 16'h001f; 
        10'b1010010111: data <= 16'h00c2; 
        10'b1010011000: data <= 16'h00aa; 
        10'b1010011001: data <= 16'h00d0; 
        10'b1010011010: data <= 16'h0095; 
        10'b1010011011: data <= 16'h0039; 
        10'b1010011100: data <= 16'h0022; 
        10'b1010011101: data <= 16'h0016; 
        10'b1010011110: data <= 16'hfffb; 
        10'b1010011111: data <= 16'hffe5; 
        10'b1010100000: data <= 16'hffed; 
        10'b1010100001: data <= 16'hffd9; 
        10'b1010100010: data <= 16'hfffe; 
        10'b1010100011: data <= 16'hfff9; 
        10'b1010100100: data <= 16'hffd6; 
        10'b1010100101: data <= 16'hff94; 
        10'b1010100110: data <= 16'hff2e; 
        10'b1010100111: data <= 16'hff63; 
        10'b1010101000: data <= 16'hff5f; 
        10'b1010101001: data <= 16'hff54; 
        10'b1010101010: data <= 16'hff55; 
        10'b1010101011: data <= 16'hff7d; 
        10'b1010101100: data <= 16'hff7c; 
        10'b1010101101: data <= 16'hffb8; 
        10'b1010101110: data <= 16'hffa3; 
        10'b1010101111: data <= 16'hff7b; 
        10'b1010110000: data <= 16'hff82; 
        10'b1010110001: data <= 16'hff9d; 
        10'b1010110010: data <= 16'hff87; 
        10'b1010110011: data <= 16'hffbf; 
        10'b1010110100: data <= 16'hffc6; 
        10'b1010110101: data <= 16'hffc6; 
        10'b1010110110: data <= 16'hffde; 
        10'b1010110111: data <= 16'hffe5; 
        10'b1010111000: data <= 16'hfffc; 
        10'b1010111001: data <= 16'h0016; 
        10'b1010111010: data <= 16'hffd3; 
        10'b1010111011: data <= 16'hffd4; 
        10'b1010111100: data <= 16'hfffe; 
        10'b1010111101: data <= 16'hffc7; 
        10'b1010111110: data <= 16'hffe3; 
        10'b1010111111: data <= 16'hffdd; 
        10'b1011000000: data <= 16'hffd3; 
        10'b1011000001: data <= 16'hffb4; 
        10'b1011000010: data <= 16'hff9a; 
        10'b1011000011: data <= 16'hff65; 
        10'b1011000100: data <= 16'hff54; 
        10'b1011000101: data <= 16'hff61; 
        10'b1011000110: data <= 16'hff70; 
        10'b1011000111: data <= 16'hff48; 
        10'b1011001000: data <= 16'hff85; 
        10'b1011001001: data <= 16'hff8d; 
        10'b1011001010: data <= 16'hff67; 
        10'b1011001011: data <= 16'hff82; 
        10'b1011001100: data <= 16'hffa2; 
        10'b1011001101: data <= 16'hffa8; 
        10'b1011001110: data <= 16'hffde; 
        10'b1011001111: data <= 16'hffb0; 
        10'b1011010000: data <= 16'hffe3; 
        10'b1011010001: data <= 16'hffe1; 
        10'b1011010010: data <= 16'hffff; 
        10'b1011010011: data <= 16'hffd5; 
        10'b1011010100: data <= 16'hfff0; 
        10'b1011010101: data <= 16'hffd6; 
        10'b1011010110: data <= 16'hffc9; 
        10'b1011010111: data <= 16'hffd6; 
        10'b1011011000: data <= 16'hffcb; 
        10'b1011011001: data <= 16'hffde; 
        10'b1011011010: data <= 16'hffe8; 
        10'b1011011011: data <= 16'h0003; 
        10'b1011011100: data <= 16'hfff7; 
        10'b1011011101: data <= 16'hffe5; 
        10'b1011011110: data <= 16'hfff5; 
        10'b1011011111: data <= 16'hfffe; 
        10'b1011100000: data <= 16'hffe4; 
        10'b1011100001: data <= 16'h0003; 
        10'b1011100010: data <= 16'hffff; 
        10'b1011100011: data <= 16'h0002; 
        10'b1011100100: data <= 16'h0005; 
        10'b1011100101: data <= 16'hfff0; 
        10'b1011100110: data <= 16'hffdb; 
        10'b1011100111: data <= 16'hffc4; 
        10'b1011101000: data <= 16'hffe0; 
        10'b1011101001: data <= 16'hffef; 
        10'b1011101010: data <= 16'hffec; 
        10'b1011101011: data <= 16'hffd5; 
        10'b1011101100: data <= 16'h0006; 
        10'b1011101101: data <= 16'hffff; 
        10'b1011101110: data <= 16'hffd6; 
        10'b1011101111: data <= 16'hffdf; 
        10'b1011110000: data <= 16'hffca; 
        10'b1011110001: data <= 16'h0002; 
        10'b1011110010: data <= 16'h0002; 
        10'b1011110011: data <= 16'hfffd; 
        10'b1011110100: data <= 16'hfffb; 
        10'b1011110101: data <= 16'hffd9; 
        10'b1011110110: data <= 16'hffcf; 
        10'b1011110111: data <= 16'hffed; 
        10'b1011111000: data <= 16'hffc9; 
        10'b1011111001: data <= 16'h000b; 
        10'b1011111010: data <= 16'h000a; 
        10'b1011111011: data <= 16'hffe0; 
        10'b1011111100: data <= 16'hfffd; 
        10'b1011111101: data <= 16'hffd5; 
        10'b1011111110: data <= 16'h0007; 
        10'b1011111111: data <= 16'hffc8; 
        10'b1100000000: data <= 16'hfffd; 
        10'b1100000001: data <= 16'hffe5; 
        10'b1100000010: data <= 16'hfff3; 
        10'b1100000011: data <= 16'hffd0; 
        10'b1100000100: data <= 16'hffec; 
        10'b1100000101: data <= 16'hffe3; 
        10'b1100000110: data <= 16'hffef; 
        10'b1100000111: data <= 16'hffeb; 
        10'b1100001000: data <= 16'hfffa; 
        10'b1100001001: data <= 16'hffc6; 
        10'b1100001010: data <= 16'hffe7; 
        10'b1100001011: data <= 16'h0002; 
        10'b1100001100: data <= 16'hffc6; 
        10'b1100001101: data <= 16'hffea; 
        10'b1100001110: data <= 16'hfff8; 
        10'b1100001111: data <= 16'hffe1; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 11) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 17'h1ff99; 
        10'b0000000001: data <= 17'h00002; 
        10'b0000000010: data <= 17'h1ffcd; 
        10'b0000000011: data <= 17'h1ffab; 
        10'b0000000100: data <= 17'h1ffcb; 
        10'b0000000101: data <= 17'h1ffb1; 
        10'b0000000110: data <= 17'h1ffdd; 
        10'b0000000111: data <= 17'h1ffe3; 
        10'b0000001000: data <= 17'h1ff96; 
        10'b0000001001: data <= 17'h1ffd5; 
        10'b0000001010: data <= 17'h1ff9e; 
        10'b0000001011: data <= 17'h1ffbf; 
        10'b0000001100: data <= 17'h00014; 
        10'b0000001101: data <= 17'h00011; 
        10'b0000001110: data <= 17'h1ff9c; 
        10'b0000001111: data <= 17'h1ffdc; 
        10'b0000010000: data <= 17'h1ffa3; 
        10'b0000010001: data <= 17'h1ffa4; 
        10'b0000010010: data <= 17'h0001b; 
        10'b0000010011: data <= 17'h00008; 
        10'b0000010100: data <= 17'h1ffb4; 
        10'b0000010101: data <= 17'h1ffdf; 
        10'b0000010110: data <= 17'h1ffbc; 
        10'b0000010111: data <= 17'h1ff90; 
        10'b0000011000: data <= 17'h1ff99; 
        10'b0000011001: data <= 17'h1ffd9; 
        10'b0000011010: data <= 17'h1fffb; 
        10'b0000011011: data <= 17'h1ffe4; 
        10'b0000011100: data <= 17'h1ffd4; 
        10'b0000011101: data <= 17'h1ffcd; 
        10'b0000011110: data <= 17'h00019; 
        10'b0000011111: data <= 17'h1ffe6; 
        10'b0000100000: data <= 17'h1ff9e; 
        10'b0000100001: data <= 17'h1ff9b; 
        10'b0000100010: data <= 17'h1ff97; 
        10'b0000100011: data <= 17'h1ffb1; 
        10'b0000100100: data <= 17'h1ffb2; 
        10'b0000100101: data <= 17'h1ffdb; 
        10'b0000100110: data <= 17'h00001; 
        10'b0000100111: data <= 17'h1ffa2; 
        10'b0000101000: data <= 17'h1ffc4; 
        10'b0000101001: data <= 17'h1ff9f; 
        10'b0000101010: data <= 17'h1ffdd; 
        10'b0000101011: data <= 17'h1ff90; 
        10'b0000101100: data <= 17'h1ffe2; 
        10'b0000101101: data <= 17'h1ffa2; 
        10'b0000101110: data <= 17'h1ffc1; 
        10'b0000101111: data <= 17'h1ffa9; 
        10'b0000110000: data <= 17'h1ffdd; 
        10'b0000110001: data <= 17'h1ffa5; 
        10'b0000110010: data <= 17'h1ff95; 
        10'b0000110011: data <= 17'h1ff8b; 
        10'b0000110100: data <= 17'h00006; 
        10'b0000110101: data <= 17'h1ffe6; 
        10'b0000110110: data <= 17'h00008; 
        10'b0000110111: data <= 17'h1ffb9; 
        10'b0000111000: data <= 17'h1ffce; 
        10'b0000111001: data <= 17'h1ff92; 
        10'b0000111010: data <= 17'h1ff9c; 
        10'b0000111011: data <= 17'h1ffff; 
        10'b0000111100: data <= 17'h1ff96; 
        10'b0000111101: data <= 17'h1ff9f; 
        10'b0000111110: data <= 17'h1ffc9; 
        10'b0000111111: data <= 17'h1ffd9; 
        10'b0001000000: data <= 17'h1fff6; 
        10'b0001000001: data <= 17'h1ffc4; 
        10'b0001000010: data <= 17'h0003a; 
        10'b0001000011: data <= 17'h00030; 
        10'b0001000100: data <= 17'h00094; 
        10'b0001000101: data <= 17'h00076; 
        10'b0001000110: data <= 17'h0006c; 
        10'b0001000111: data <= 17'h0002b; 
        10'b0001001000: data <= 17'h00091; 
        10'b0001001001: data <= 17'h00032; 
        10'b0001001010: data <= 17'h0002a; 
        10'b0001001011: data <= 17'h1ffb6; 
        10'b0001001100: data <= 17'h1fffe; 
        10'b0001001101: data <= 17'h1ffde; 
        10'b0001001110: data <= 17'h1ff6a; 
        10'b0001001111: data <= 17'h1ffcb; 
        10'b0001010000: data <= 17'h1fff0; 
        10'b0001010001: data <= 17'h00024; 
        10'b0001010010: data <= 17'h1ffd5; 
        10'b0001010011: data <= 17'h1ffc3; 
        10'b0001010100: data <= 17'h1ffb7; 
        10'b0001010101: data <= 17'h1ffad; 
        10'b0001010110: data <= 17'h1ffe8; 
        10'b0001010111: data <= 17'h1ffb4; 
        10'b0001011000: data <= 17'h00015; 
        10'b0001011001: data <= 17'h1ffa3; 
        10'b0001011010: data <= 17'h1ffde; 
        10'b0001011011: data <= 17'h00000; 
        10'b0001011100: data <= 17'h0001a; 
        10'b0001011101: data <= 17'h000ec; 
        10'b0001011110: data <= 17'h00171; 
        10'b0001011111: data <= 17'h0016e; 
        10'b0001100000: data <= 17'h0015e; 
        10'b0001100001: data <= 17'h00203; 
        10'b0001100010: data <= 17'h00119; 
        10'b0001100011: data <= 17'h0007d; 
        10'b0001100100: data <= 17'h000ed; 
        10'b0001100101: data <= 17'h0006d; 
        10'b0001100110: data <= 17'h1ff99; 
        10'b0001100111: data <= 17'h1ffe7; 
        10'b0001101000: data <= 17'h1ff8c; 
        10'b0001101001: data <= 17'h1ff78; 
        10'b0001101010: data <= 17'h1ff59; 
        10'b0001101011: data <= 17'h1ffad; 
        10'b0001101100: data <= 17'h0000c; 
        10'b0001101101: data <= 17'h00027; 
        10'b0001101110: data <= 17'h1ffa4; 
        10'b0001101111: data <= 17'h1ffed; 
        10'b0001110000: data <= 17'h1ffaf; 
        10'b0001110001: data <= 17'h1ffc8; 
        10'b0001110010: data <= 17'h0001c; 
        10'b0001110011: data <= 17'h1ff88; 
        10'b0001110100: data <= 17'h1ff96; 
        10'b0001110101: data <= 17'h1ffde; 
        10'b0001110110: data <= 17'h00037; 
        10'b0001110111: data <= 17'h00035; 
        10'b0001111000: data <= 17'h00098; 
        10'b0001111001: data <= 17'h001c3; 
        10'b0001111010: data <= 17'h001c8; 
        10'b0001111011: data <= 17'h0023d; 
        10'b0001111100: data <= 17'h001e4; 
        10'b0001111101: data <= 17'h00180; 
        10'b0001111110: data <= 17'h0015d; 
        10'b0001111111: data <= 17'h0009a; 
        10'b0010000000: data <= 17'h000ce; 
        10'b0010000001: data <= 17'h000bf; 
        10'b0010000010: data <= 17'h1ffc7; 
        10'b0010000011: data <= 17'h1ffa0; 
        10'b0010000100: data <= 17'h1ffb6; 
        10'b0010000101: data <= 17'h1ff1d; 
        10'b0010000110: data <= 17'h1feee; 
        10'b0010000111: data <= 17'h1fef8; 
        10'b0010001000: data <= 17'h1ffde; 
        10'b0010001001: data <= 17'h1ffde; 
        10'b0010001010: data <= 17'h1ff92; 
        10'b0010001011: data <= 17'h1ffeb; 
        10'b0010001100: data <= 17'h00009; 
        10'b0010001101: data <= 17'h1ffdc; 
        10'b0010001110: data <= 17'h1ffa9; 
        10'b0010001111: data <= 17'h1ff8c; 
        10'b0010010000: data <= 17'h1ffa1; 
        10'b0010010001: data <= 17'h1ffae; 
        10'b0010010010: data <= 17'h00033; 
        10'b0010010011: data <= 17'h000dd; 
        10'b0010010100: data <= 17'h00132; 
        10'b0010010101: data <= 17'h0020b; 
        10'b0010010110: data <= 17'h00244; 
        10'b0010010111: data <= 17'h0025d; 
        10'b0010011000: data <= 17'h0022a; 
        10'b0010011001: data <= 17'h0026d; 
        10'b0010011010: data <= 17'h0023f; 
        10'b0010011011: data <= 17'h00215; 
        10'b0010011100: data <= 17'h00243; 
        10'b0010011101: data <= 17'h001d4; 
        10'b0010011110: data <= 17'h00152; 
        10'b0010011111: data <= 17'h1ff71; 
        10'b0010100000: data <= 17'h1ff76; 
        10'b0010100001: data <= 17'h1ff1f; 
        10'b0010100010: data <= 17'h1ff1b; 
        10'b0010100011: data <= 17'h1fe9d; 
        10'b0010100100: data <= 17'h1ff67; 
        10'b0010100101: data <= 17'h1ffa9; 
        10'b0010100110: data <= 17'h0000e; 
        10'b0010100111: data <= 17'h1ffbc; 
        10'b0010101000: data <= 17'h1ffd2; 
        10'b0010101001: data <= 17'h1ffad; 
        10'b0010101010: data <= 17'h00013; 
        10'b0010101011: data <= 17'h1ffd3; 
        10'b0010101100: data <= 17'h1ffc6; 
        10'b0010101101: data <= 17'h00025; 
        10'b0010101110: data <= 17'h000d8; 
        10'b0010101111: data <= 17'h001a1; 
        10'b0010110000: data <= 17'h0013f; 
        10'b0010110001: data <= 17'h0016a; 
        10'b0010110010: data <= 17'h001ea; 
        10'b0010110011: data <= 17'h00133; 
        10'b0010110100: data <= 17'h00146; 
        10'b0010110101: data <= 17'h001a5; 
        10'b0010110110: data <= 17'h00174; 
        10'b0010110111: data <= 17'h000ca; 
        10'b0010111000: data <= 17'h000e0; 
        10'b0010111001: data <= 17'h0003a; 
        10'b0010111010: data <= 17'h0002b; 
        10'b0010111011: data <= 17'h1ff7d; 
        10'b0010111100: data <= 17'h1ffa9; 
        10'b0010111101: data <= 17'h1fee1; 
        10'b0010111110: data <= 17'h1fee4; 
        10'b0010111111: data <= 17'h1fe73; 
        10'b0011000000: data <= 17'h1ff14; 
        10'b0011000001: data <= 17'h1ff7c; 
        10'b0011000010: data <= 17'h00011; 
        10'b0011000011: data <= 17'h1fff3; 
        10'b0011000100: data <= 17'h1ffc3; 
        10'b0011000101: data <= 17'h0000c; 
        10'b0011000110: data <= 17'h0000d; 
        10'b0011000111: data <= 17'h1ffc8; 
        10'b0011001000: data <= 17'h00006; 
        10'b0011001001: data <= 17'h00074; 
        10'b0011001010: data <= 17'h00116; 
        10'b0011001011: data <= 17'h00192; 
        10'b0011001100: data <= 17'h00149; 
        10'b0011001101: data <= 17'h00133; 
        10'b0011001110: data <= 17'h00075; 
        10'b0011001111: data <= 17'h0008b; 
        10'b0011010000: data <= 17'h00018; 
        10'b0011010001: data <= 17'h000d8; 
        10'b0011010010: data <= 17'h0010a; 
        10'b0011010011: data <= 17'h00038; 
        10'b0011010100: data <= 17'h00024; 
        10'b0011010101: data <= 17'h1feaf; 
        10'b0011010110: data <= 17'h1ff8e; 
        10'b0011010111: data <= 17'h1ffa1; 
        10'b0011011000: data <= 17'h1ff94; 
        10'b0011011001: data <= 17'h1ff82; 
        10'b0011011010: data <= 17'h1ffa2; 
        10'b0011011011: data <= 17'h1feb9; 
        10'b0011011100: data <= 17'h1ff1e; 
        10'b0011011101: data <= 17'h1ffbb; 
        10'b0011011110: data <= 17'h1ffa9; 
        10'b0011011111: data <= 17'h1ff96; 
        10'b0011100000: data <= 17'h1ffe8; 
        10'b0011100001: data <= 17'h00010; 
        10'b0011100010: data <= 17'h1ffd3; 
        10'b0011100011: data <= 17'h0000f; 
        10'b0011100100: data <= 17'h0003d; 
        10'b0011100101: data <= 17'h000bc; 
        10'b0011100110: data <= 17'h00088; 
        10'b0011100111: data <= 17'h000c0; 
        10'b0011101000: data <= 17'h000c3; 
        10'b0011101001: data <= 17'h000d8; 
        10'b0011101010: data <= 17'h000d9; 
        10'b0011101011: data <= 17'h000f8; 
        10'b0011101100: data <= 17'h00094; 
        10'b0011101101: data <= 17'h000b0; 
        10'b0011101110: data <= 17'h001d1; 
        10'b0011101111: data <= 17'h00105; 
        10'b0011110000: data <= 17'h1ffe0; 
        10'b0011110001: data <= 17'h1ff80; 
        10'b0011110010: data <= 17'h1fffd; 
        10'b0011110011: data <= 17'h00067; 
        10'b0011110100: data <= 17'h00002; 
        10'b0011110101: data <= 17'h1ffb9; 
        10'b0011110110: data <= 17'h1ff43; 
        10'b0011110111: data <= 17'h1fe83; 
        10'b0011111000: data <= 17'h1fedc; 
        10'b0011111001: data <= 17'h1ff86; 
        10'b0011111010: data <= 17'h1ffc7; 
        10'b0011111011: data <= 17'h1ffa2; 
        10'b0011111100: data <= 17'h1ffb0; 
        10'b0011111101: data <= 17'h1ffec; 
        10'b0011111110: data <= 17'h1fffc; 
        10'b0011111111: data <= 17'h00031; 
        10'b0100000000: data <= 17'h0005f; 
        10'b0100000001: data <= 17'h000d3; 
        10'b0100000010: data <= 17'h0004a; 
        10'b0100000011: data <= 17'h0000e; 
        10'b0100000100: data <= 17'h1ffb7; 
        10'b0100000101: data <= 17'h00071; 
        10'b0100000110: data <= 17'h00058; 
        10'b0100000111: data <= 17'h00072; 
        10'b0100001000: data <= 17'h0001e; 
        10'b0100001001: data <= 17'h1fff4; 
        10'b0100001010: data <= 17'h0012f; 
        10'b0100001011: data <= 17'h00148; 
        10'b0100001100: data <= 17'h00071; 
        10'b0100001101: data <= 17'h00009; 
        10'b0100001110: data <= 17'h1ffe2; 
        10'b0100001111: data <= 17'h1fffd; 
        10'b0100010000: data <= 17'h1fff2; 
        10'b0100010001: data <= 17'h1fff9; 
        10'b0100010010: data <= 17'h1ff88; 
        10'b0100010011: data <= 17'h1febc; 
        10'b0100010100: data <= 17'h1feeb; 
        10'b0100010101: data <= 17'h1ffa6; 
        10'b0100010110: data <= 17'h0000e; 
        10'b0100010111: data <= 17'h1ff98; 
        10'b0100011000: data <= 17'h00014; 
        10'b0100011001: data <= 17'h1ffe8; 
        10'b0100011010: data <= 17'h1ffd0; 
        10'b0100011011: data <= 17'h1ffbc; 
        10'b0100011100: data <= 17'h0000e; 
        10'b0100011101: data <= 17'h1ffcd; 
        10'b0100011110: data <= 17'h1ff97; 
        10'b0100011111: data <= 17'h1fe01; 
        10'b0100100000: data <= 17'h1fe36; 
        10'b0100100001: data <= 17'h1fea6; 
        10'b0100100010: data <= 17'h1fdf0; 
        10'b0100100011: data <= 17'h1fdb6; 
        10'b0100100100: data <= 17'h1fd56; 
        10'b0100100101: data <= 17'h1fd02; 
        10'b0100100110: data <= 17'h1febf; 
        10'b0100100111: data <= 17'h0003a; 
        10'b0100101000: data <= 17'h00053; 
        10'b0100101001: data <= 17'h0000e; 
        10'b0100101010: data <= 17'h0002b; 
        10'b0100101011: data <= 17'h1ffc2; 
        10'b0100101100: data <= 17'h1ffd3; 
        10'b0100101101: data <= 17'h1ffc2; 
        10'b0100101110: data <= 17'h1ff60; 
        10'b0100101111: data <= 17'h1fe8b; 
        10'b0100110000: data <= 17'h1ff33; 
        10'b0100110001: data <= 17'h1fff7; 
        10'b0100110010: data <= 17'h1fff7; 
        10'b0100110011: data <= 17'h1ffaa; 
        10'b0100110100: data <= 17'h1ff95; 
        10'b0100110101: data <= 17'h0001a; 
        10'b0100110110: data <= 17'h1fff5; 
        10'b0100110111: data <= 17'h1ff9e; 
        10'b0100111000: data <= 17'h1ff40; 
        10'b0100111001: data <= 17'h1fe5d; 
        10'b0100111010: data <= 17'h1fd31; 
        10'b0100111011: data <= 17'h1fc0a; 
        10'b0100111100: data <= 17'h1fc32; 
        10'b0100111101: data <= 17'h1fb85; 
        10'b0100111110: data <= 17'h1fb82; 
        10'b0100111111: data <= 17'h1fbe6; 
        10'b0101000000: data <= 17'h1fba5; 
        10'b0101000001: data <= 17'h1fab2; 
        10'b0101000010: data <= 17'h1fbeb; 
        10'b0101000011: data <= 17'h1fe0c; 
        10'b0101000100: data <= 17'h1ff53; 
        10'b0101000101: data <= 17'h1ff6b; 
        10'b0101000110: data <= 17'h1ff71; 
        10'b0101000111: data <= 17'h1ffe3; 
        10'b0101001000: data <= 17'h1ffaa; 
        10'b0101001001: data <= 17'h1ffa6; 
        10'b0101001010: data <= 17'h1ff13; 
        10'b0101001011: data <= 17'h1ff5e; 
        10'b0101001100: data <= 17'h1ffe3; 
        10'b0101001101: data <= 17'h1ffc8; 
        10'b0101001110: data <= 17'h1ffa7; 
        10'b0101001111: data <= 17'h1ffe7; 
        10'b0101010000: data <= 17'h1ffdb; 
        10'b0101010001: data <= 17'h1ffe2; 
        10'b0101010010: data <= 17'h0000b; 
        10'b0101010011: data <= 17'h1ffd3; 
        10'b0101010100: data <= 17'h1ff32; 
        10'b0101010101: data <= 17'h1fd90; 
        10'b0101010110: data <= 17'h1fb42; 
        10'b0101010111: data <= 17'h1fa33; 
        10'b0101011000: data <= 17'h1fa97; 
        10'b0101011001: data <= 17'h1fadf; 
        10'b0101011010: data <= 17'h1fb50; 
        10'b0101011011: data <= 17'h1fb9d; 
        10'b0101011100: data <= 17'h1fba1; 
        10'b0101011101: data <= 17'h1fb73; 
        10'b0101011110: data <= 17'h1fc43; 
        10'b0101011111: data <= 17'h1fd82; 
        10'b0101100000: data <= 17'h1fe4a; 
        10'b0101100001: data <= 17'h1fe77; 
        10'b0101100010: data <= 17'h1ff3a; 
        10'b0101100011: data <= 17'h00001; 
        10'b0101100100: data <= 17'h1fffc; 
        10'b0101100101: data <= 17'h1ff91; 
        10'b0101100110: data <= 17'h1ff03; 
        10'b0101100111: data <= 17'h1fe80; 
        10'b0101101000: data <= 17'h1ffd1; 
        10'b0101101001: data <= 17'h1ffc0; 
        10'b0101101010: data <= 17'h0001d; 
        10'b0101101011: data <= 17'h1ffe1; 
        10'b0101101100: data <= 17'h1ffb3; 
        10'b0101101101: data <= 17'h1ffcd; 
        10'b0101101110: data <= 17'h0001b; 
        10'b0101101111: data <= 17'h1ffb0; 
        10'b0101110000: data <= 17'h1feb2; 
        10'b0101110001: data <= 17'h1fced; 
        10'b0101110010: data <= 17'h1fb1f; 
        10'b0101110011: data <= 17'h1fb86; 
        10'b0101110100: data <= 17'h1fbd2; 
        10'b0101110101: data <= 17'h1fd21; 
        10'b0101110110: data <= 17'h1fdf7; 
        10'b0101110111: data <= 17'h1ff0c; 
        10'b0101111000: data <= 17'h1fe7e; 
        10'b0101111001: data <= 17'h1ff50; 
        10'b0101111010: data <= 17'h1fe47; 
        10'b0101111011: data <= 17'h1fe3e; 
        10'b0101111100: data <= 17'h1fdeb; 
        10'b0101111101: data <= 17'h1fe7f; 
        10'b0101111110: data <= 17'h1ff2c; 
        10'b0101111111: data <= 17'h1ffd7; 
        10'b0110000000: data <= 17'h1ffc2; 
        10'b0110000001: data <= 17'h1ff77; 
        10'b0110000010: data <= 17'h1fec2; 
        10'b0110000011: data <= 17'h1fedf; 
        10'b0110000100: data <= 17'h1ff6e; 
        10'b0110000101: data <= 17'h00025; 
        10'b0110000110: data <= 17'h1ffcf; 
        10'b0110000111: data <= 17'h1fffd; 
        10'b0110001000: data <= 17'h00011; 
        10'b0110001001: data <= 17'h1ffe5; 
        10'b0110001010: data <= 17'h00003; 
        10'b0110001011: data <= 17'h1ffbd; 
        10'b0110001100: data <= 17'h1ff80; 
        10'b0110001101: data <= 17'h1fded; 
        10'b0110001110: data <= 17'h1fd60; 
        10'b0110001111: data <= 17'h1fddc; 
        10'b0110010000: data <= 17'h1ff24; 
        10'b0110010001: data <= 17'h1ffda; 
        10'b0110010010: data <= 17'h00089; 
        10'b0110010011: data <= 17'h000b5; 
        10'b0110010100: data <= 17'h000d7; 
        10'b0110010101: data <= 17'h0014f; 
        10'b0110010110: data <= 17'h00017; 
        10'b0110010111: data <= 17'h1ff2a; 
        10'b0110011000: data <= 17'h1ff61; 
        10'b0110011001: data <= 17'h1feec; 
        10'b0110011010: data <= 17'h1ffd2; 
        10'b0110011011: data <= 17'h1ff4e; 
        10'b0110011100: data <= 17'h1ffc8; 
        10'b0110011101: data <= 17'h1ff33; 
        10'b0110011110: data <= 17'h1fe90; 
        10'b0110011111: data <= 17'h1fef5; 
        10'b0110100000: data <= 17'h1ffcc; 
        10'b0110100001: data <= 17'h00082; 
        10'b0110100010: data <= 17'h00094; 
        10'b0110100011: data <= 17'h1ffae; 
        10'b0110100100: data <= 17'h1ffc7; 
        10'b0110100101: data <= 17'h1ffd3; 
        10'b0110100110: data <= 17'h1ffc5; 
        10'b0110100111: data <= 17'h00079; 
        10'b0110101000: data <= 17'h0003b; 
        10'b0110101001: data <= 17'h0001b; 
        10'b0110101010: data <= 17'h00090; 
        10'b0110101011: data <= 17'h000a8; 
        10'b0110101100: data <= 17'h00139; 
        10'b0110101101: data <= 17'h000dd; 
        10'b0110101110: data <= 17'h00109; 
        10'b0110101111: data <= 17'h0009c; 
        10'b0110110000: data <= 17'h0008a; 
        10'b0110110001: data <= 17'h00144; 
        10'b0110110010: data <= 17'h00018; 
        10'b0110110011: data <= 17'h0007f; 
        10'b0110110100: data <= 17'h00012; 
        10'b0110110101: data <= 17'h1feff; 
        10'b0110110110: data <= 17'h1ff0c; 
        10'b0110110111: data <= 17'h1ff6a; 
        10'b0110111000: data <= 17'h1ff93; 
        10'b0110111001: data <= 17'h1ff5b; 
        10'b0110111010: data <= 17'h1feb3; 
        10'b0110111011: data <= 17'h1ff55; 
        10'b0110111100: data <= 17'h00066; 
        10'b0110111101: data <= 17'h000af; 
        10'b0110111110: data <= 17'h0005e; 
        10'b0110111111: data <= 17'h1ffa3; 
        10'b0111000000: data <= 17'h1ffb9; 
        10'b0111000001: data <= 17'h1ff91; 
        10'b0111000010: data <= 17'h1ff82; 
        10'b0111000011: data <= 17'h00081; 
        10'b0111000100: data <= 17'h0010f; 
        10'b0111000101: data <= 17'h001ba; 
        10'b0111000110: data <= 17'h001c3; 
        10'b0111000111: data <= 17'h0010c; 
        10'b0111001000: data <= 17'h0006f; 
        10'b0111001001: data <= 17'h000e7; 
        10'b0111001010: data <= 17'h000d7; 
        10'b0111001011: data <= 17'h000c4; 
        10'b0111001100: data <= 17'h00194; 
        10'b0111001101: data <= 17'h00164; 
        10'b0111001110: data <= 17'h0004b; 
        10'b0111001111: data <= 17'h1ffd5; 
        10'b0111010000: data <= 17'h1fffe; 
        10'b0111010001: data <= 17'h1ff59; 
        10'b0111010010: data <= 17'h1ff6e; 
        10'b0111010011: data <= 17'h1ff00; 
        10'b0111010100: data <= 17'h1ffa5; 
        10'b0111010101: data <= 17'h0000e; 
        10'b0111010110: data <= 17'h00038; 
        10'b0111010111: data <= 17'h00077; 
        10'b0111011000: data <= 17'h0017a; 
        10'b0111011001: data <= 17'h001d4; 
        10'b0111011010: data <= 17'h0004e; 
        10'b0111011011: data <= 17'h1ffb7; 
        10'b0111011100: data <= 17'h1ffc4; 
        10'b0111011101: data <= 17'h00015; 
        10'b0111011110: data <= 17'h1ffd1; 
        10'b0111011111: data <= 17'h0009d; 
        10'b0111100000: data <= 17'h001cf; 
        10'b0111100001: data <= 17'h00285; 
        10'b0111100010: data <= 17'h0024d; 
        10'b0111100011: data <= 17'h00194; 
        10'b0111100100: data <= 17'h00119; 
        10'b0111100101: data <= 17'h00155; 
        10'b0111100110: data <= 17'h0020c; 
        10'b0111100111: data <= 17'h001ad; 
        10'b0111101000: data <= 17'h001ec; 
        10'b0111101001: data <= 17'h000e6; 
        10'b0111101010: data <= 17'h00077; 
        10'b0111101011: data <= 17'h000a0; 
        10'b0111101100: data <= 17'h000a2; 
        10'b0111101101: data <= 17'h1ffe7; 
        10'b0111101110: data <= 17'h00069; 
        10'b0111101111: data <= 17'h1ffbd; 
        10'b0111110000: data <= 17'h000c1; 
        10'b0111110001: data <= 17'h000ce; 
        10'b0111110010: data <= 17'h00099; 
        10'b0111110011: data <= 17'h000d5; 
        10'b0111110100: data <= 17'h0025d; 
        10'b0111110101: data <= 17'h0020d; 
        10'b0111110110: data <= 17'h00078; 
        10'b0111110111: data <= 17'h00010; 
        10'b0111111000: data <= 17'h1fff2; 
        10'b0111111001: data <= 17'h1fff9; 
        10'b0111111010: data <= 17'h1ff61; 
        10'b0111111011: data <= 17'h0002a; 
        10'b0111111100: data <= 17'h001f6; 
        10'b0111111101: data <= 17'h00350; 
        10'b0111111110: data <= 17'h0031d; 
        10'b0111111111: data <= 17'h0023e; 
        10'b1000000000: data <= 17'h0017f; 
        10'b1000000001: data <= 17'h001aa; 
        10'b1000000010: data <= 17'h0028a; 
        10'b1000000011: data <= 17'h0024c; 
        10'b1000000100: data <= 17'h003a8; 
        10'b1000000101: data <= 17'h002ab; 
        10'b1000000110: data <= 17'h00255; 
        10'b1000000111: data <= 17'h00122; 
        10'b1000001000: data <= 17'h000c8; 
        10'b1000001001: data <= 17'h0016f; 
        10'b1000001010: data <= 17'h000ed; 
        10'b1000001011: data <= 17'h000a1; 
        10'b1000001100: data <= 17'h001b1; 
        10'b1000001101: data <= 17'h001bf; 
        10'b1000001110: data <= 17'h001e8; 
        10'b1000001111: data <= 17'h00284; 
        10'b1000010000: data <= 17'h0031f; 
        10'b1000010001: data <= 17'h001cd; 
        10'b1000010010: data <= 17'h1ffd4; 
        10'b1000010011: data <= 17'h1ffa1; 
        10'b1000010100: data <= 17'h1ffaf; 
        10'b1000010101: data <= 17'h1ffb4; 
        10'b1000010110: data <= 17'h1ff91; 
        10'b1000010111: data <= 17'h1fffe; 
        10'b1000011000: data <= 17'h00114; 
        10'b1000011001: data <= 17'h00203; 
        10'b1000011010: data <= 17'h0028a; 
        10'b1000011011: data <= 17'h00234; 
        10'b1000011100: data <= 17'h00208; 
        10'b1000011101: data <= 17'h00227; 
        10'b1000011110: data <= 17'h0020f; 
        10'b1000011111: data <= 17'h00230; 
        10'b1000100000: data <= 17'h00273; 
        10'b1000100001: data <= 17'h001e2; 
        10'b1000100010: data <= 17'h00138; 
        10'b1000100011: data <= 17'h00094; 
        10'b1000100100: data <= 17'h000e6; 
        10'b1000100101: data <= 17'h0018f; 
        10'b1000100110: data <= 17'h000c1; 
        10'b1000100111: data <= 17'h000bc; 
        10'b1000101000: data <= 17'h00142; 
        10'b1000101001: data <= 17'h00191; 
        10'b1000101010: data <= 17'h0020c; 
        10'b1000101011: data <= 17'h00232; 
        10'b1000101100: data <= 17'h001e5; 
        10'b1000101101: data <= 17'h000fe; 
        10'b1000101110: data <= 17'h00015; 
        10'b1000101111: data <= 17'h00006; 
        10'b1000110000: data <= 17'h1ff9c; 
        10'b1000110001: data <= 17'h1fff8; 
        10'b1000110010: data <= 17'h1ffe5; 
        10'b1000110011: data <= 17'h1ff76; 
        10'b1000110100: data <= 17'h000f5; 
        10'b1000110101: data <= 17'h0012e; 
        10'b1000110110: data <= 17'h001d5; 
        10'b1000110111: data <= 17'h0028c; 
        10'b1000111000: data <= 17'h0026c; 
        10'b1000111001: data <= 17'h0019a; 
        10'b1000111010: data <= 17'h0018b; 
        10'b1000111011: data <= 17'h00295; 
        10'b1000111100: data <= 17'h0016f; 
        10'b1000111101: data <= 17'h0007a; 
        10'b1000111110: data <= 17'h00051; 
        10'b1000111111: data <= 17'h00064; 
        10'b1001000000: data <= 17'h00081; 
        10'b1001000001: data <= 17'h00006; 
        10'b1001000010: data <= 17'h0011e; 
        10'b1001000011: data <= 17'h001be; 
        10'b1001000100: data <= 17'h0012f; 
        10'b1001000101: data <= 17'h001ae; 
        10'b1001000110: data <= 17'h00257; 
        10'b1001000111: data <= 17'h00208; 
        10'b1001001000: data <= 17'h00176; 
        10'b1001001001: data <= 17'h000b1; 
        10'b1001001010: data <= 17'h1fffe; 
        10'b1001001011: data <= 17'h1ffef; 
        10'b1001001100: data <= 17'h1ffd9; 
        10'b1001001101: data <= 17'h1ffa0; 
        10'b1001001110: data <= 17'h1ffef; 
        10'b1001001111: data <= 17'h1ffc9; 
        10'b1001010000: data <= 17'h00033; 
        10'b1001010001: data <= 17'h00082; 
        10'b1001010010: data <= 17'h00145; 
        10'b1001010011: data <= 17'h0016e; 
        10'b1001010100: data <= 17'h00142; 
        10'b1001010101: data <= 17'h00192; 
        10'b1001010110: data <= 17'h00164; 
        10'b1001010111: data <= 17'h0015d; 
        10'b1001011000: data <= 17'h00089; 
        10'b1001011001: data <= 17'h00041; 
        10'b1001011010: data <= 17'h1ffdd; 
        10'b1001011011: data <= 17'h0000f; 
        10'b1001011100: data <= 17'h000ae; 
        10'b1001011101: data <= 17'h000be; 
        10'b1001011110: data <= 17'h001a1; 
        10'b1001011111: data <= 17'h001b7; 
        10'b1001100000: data <= 17'h000c0; 
        10'b1001100001: data <= 17'h001ae; 
        10'b1001100010: data <= 17'h00213; 
        10'b1001100011: data <= 17'h0025d; 
        10'b1001100100: data <= 17'h0012a; 
        10'b1001100101: data <= 17'h00076; 
        10'b1001100110: data <= 17'h0001b; 
        10'b1001100111: data <= 17'h1fff3; 
        10'b1001101000: data <= 17'h1ff9b; 
        10'b1001101001: data <= 17'h1ffe5; 
        10'b1001101010: data <= 17'h1ffa9; 
        10'b1001101011: data <= 17'h0001d; 
        10'b1001101100: data <= 17'h00066; 
        10'b1001101101: data <= 17'h00025; 
        10'b1001101110: data <= 17'h000dd; 
        10'b1001101111: data <= 17'h000c2; 
        10'b1001110000: data <= 17'h000b5; 
        10'b1001110001: data <= 17'h000fe; 
        10'b1001110010: data <= 17'h000fd; 
        10'b1001110011: data <= 17'h0012b; 
        10'b1001110100: data <= 17'h00020; 
        10'b1001110101: data <= 17'h1ff13; 
        10'b1001110110: data <= 17'h1fed6; 
        10'b1001110111: data <= 17'h1ff57; 
        10'b1001111000: data <= 17'h1ff61; 
        10'b1001111001: data <= 17'h0007b; 
        10'b1001111010: data <= 17'h00184; 
        10'b1001111011: data <= 17'h001ef; 
        10'b1001111100: data <= 17'h001c2; 
        10'b1001111101: data <= 17'h001af; 
        10'b1001111110: data <= 17'h00176; 
        10'b1001111111: data <= 17'h0019c; 
        10'b1010000000: data <= 17'h00099; 
        10'b1010000001: data <= 17'h1ffef; 
        10'b1010000010: data <= 17'h1ffe6; 
        10'b1010000011: data <= 17'h1ffb8; 
        10'b1010000100: data <= 17'h1ffe7; 
        10'b1010000101: data <= 17'h1ffea; 
        10'b1010000110: data <= 17'h1ffd3; 
        10'b1010000111: data <= 17'h1ffcc; 
        10'b1010001000: data <= 17'h1ffc6; 
        10'b1010001001: data <= 17'h1ff8d; 
        10'b1010001010: data <= 17'h1ff73; 
        10'b1010001011: data <= 17'h1ff85; 
        10'b1010001100: data <= 17'h1ff37; 
        10'b1010001101: data <= 17'h1ff8a; 
        10'b1010001110: data <= 17'h1ffb1; 
        10'b1010001111: data <= 17'h00066; 
        10'b1010010000: data <= 17'h00009; 
        10'b1010010001: data <= 17'h1ff62; 
        10'b1010010010: data <= 17'h1ff2a; 
        10'b1010010011: data <= 17'h1fee8; 
        10'b1010010100: data <= 17'h1fed0; 
        10'b1010010101: data <= 17'h1ff62; 
        10'b1010010110: data <= 17'h0003e; 
        10'b1010010111: data <= 17'h00183; 
        10'b1010011000: data <= 17'h00153; 
        10'b1010011001: data <= 17'h0019f; 
        10'b1010011010: data <= 17'h0012a; 
        10'b1010011011: data <= 17'h00072; 
        10'b1010011100: data <= 17'h00045; 
        10'b1010011101: data <= 17'h0002c; 
        10'b1010011110: data <= 17'h1fff6; 
        10'b1010011111: data <= 17'h1ffcb; 
        10'b1010100000: data <= 17'h1ffda; 
        10'b1010100001: data <= 17'h1ffb1; 
        10'b1010100010: data <= 17'h1fffc; 
        10'b1010100011: data <= 17'h1fff3; 
        10'b1010100100: data <= 17'h1ffad; 
        10'b1010100101: data <= 17'h1ff27; 
        10'b1010100110: data <= 17'h1fe5d; 
        10'b1010100111: data <= 17'h1fec7; 
        10'b1010101000: data <= 17'h1febe; 
        10'b1010101001: data <= 17'h1fea8; 
        10'b1010101010: data <= 17'h1feab; 
        10'b1010101011: data <= 17'h1fefa; 
        10'b1010101100: data <= 17'h1fef8; 
        10'b1010101101: data <= 17'h1ff71; 
        10'b1010101110: data <= 17'h1ff45; 
        10'b1010101111: data <= 17'h1fef6; 
        10'b1010110000: data <= 17'h1ff03; 
        10'b1010110001: data <= 17'h1ff3a; 
        10'b1010110010: data <= 17'h1ff0e; 
        10'b1010110011: data <= 17'h1ff7d; 
        10'b1010110100: data <= 17'h1ff8c; 
        10'b1010110101: data <= 17'h1ff8d; 
        10'b1010110110: data <= 17'h1ffbd; 
        10'b1010110111: data <= 17'h1ffcb; 
        10'b1010111000: data <= 17'h1fff8; 
        10'b1010111001: data <= 17'h0002b; 
        10'b1010111010: data <= 17'h1ffa6; 
        10'b1010111011: data <= 17'h1ffa8; 
        10'b1010111100: data <= 17'h1fffc; 
        10'b1010111101: data <= 17'h1ff8f; 
        10'b1010111110: data <= 17'h1ffc6; 
        10'b1010111111: data <= 17'h1ffbb; 
        10'b1011000000: data <= 17'h1ffa7; 
        10'b1011000001: data <= 17'h1ff67; 
        10'b1011000010: data <= 17'h1ff35; 
        10'b1011000011: data <= 17'h1feca; 
        10'b1011000100: data <= 17'h1fea8; 
        10'b1011000101: data <= 17'h1fec1; 
        10'b1011000110: data <= 17'h1fedf; 
        10'b1011000111: data <= 17'h1fe90; 
        10'b1011001000: data <= 17'h1ff0a; 
        10'b1011001001: data <= 17'h1ff19; 
        10'b1011001010: data <= 17'h1fece; 
        10'b1011001011: data <= 17'h1ff04; 
        10'b1011001100: data <= 17'h1ff45; 
        10'b1011001101: data <= 17'h1ff50; 
        10'b1011001110: data <= 17'h1ffbd; 
        10'b1011001111: data <= 17'h1ff5f; 
        10'b1011010000: data <= 17'h1ffc6; 
        10'b1011010001: data <= 17'h1ffc2; 
        10'b1011010010: data <= 17'h1fffd; 
        10'b1011010011: data <= 17'h1ffa9; 
        10'b1011010100: data <= 17'h1ffe0; 
        10'b1011010101: data <= 17'h1ffab; 
        10'b1011010110: data <= 17'h1ff92; 
        10'b1011010111: data <= 17'h1ffad; 
        10'b1011011000: data <= 17'h1ff96; 
        10'b1011011001: data <= 17'h1ffbd; 
        10'b1011011010: data <= 17'h1ffcf; 
        10'b1011011011: data <= 17'h00005; 
        10'b1011011100: data <= 17'h1ffef; 
        10'b1011011101: data <= 17'h1ffcb; 
        10'b1011011110: data <= 17'h1ffeb; 
        10'b1011011111: data <= 17'h1fffc; 
        10'b1011100000: data <= 17'h1ffc9; 
        10'b1011100001: data <= 17'h00006; 
        10'b1011100010: data <= 17'h1fffe; 
        10'b1011100011: data <= 17'h00004; 
        10'b1011100100: data <= 17'h0000a; 
        10'b1011100101: data <= 17'h1ffe0; 
        10'b1011100110: data <= 17'h1ffb7; 
        10'b1011100111: data <= 17'h1ff88; 
        10'b1011101000: data <= 17'h1ffc1; 
        10'b1011101001: data <= 17'h1ffdf; 
        10'b1011101010: data <= 17'h1ffd8; 
        10'b1011101011: data <= 17'h1ffaa; 
        10'b1011101100: data <= 17'h0000b; 
        10'b1011101101: data <= 17'h1fffe; 
        10'b1011101110: data <= 17'h1ffab; 
        10'b1011101111: data <= 17'h1ffbd; 
        10'b1011110000: data <= 17'h1ff94; 
        10'b1011110001: data <= 17'h00005; 
        10'b1011110010: data <= 17'h00003; 
        10'b1011110011: data <= 17'h1fffa; 
        10'b1011110100: data <= 17'h1fff7; 
        10'b1011110101: data <= 17'h1ffb2; 
        10'b1011110110: data <= 17'h1ff9f; 
        10'b1011110111: data <= 17'h1ffd9; 
        10'b1011111000: data <= 17'h1ff93; 
        10'b1011111001: data <= 17'h00017; 
        10'b1011111010: data <= 17'h00014; 
        10'b1011111011: data <= 17'h1ffc1; 
        10'b1011111100: data <= 17'h1fff9; 
        10'b1011111101: data <= 17'h1ffaa; 
        10'b1011111110: data <= 17'h0000f; 
        10'b1011111111: data <= 17'h1ff90; 
        10'b1100000000: data <= 17'h1fffa; 
        10'b1100000001: data <= 17'h1ffca; 
        10'b1100000010: data <= 17'h1ffe7; 
        10'b1100000011: data <= 17'h1ffa1; 
        10'b1100000100: data <= 17'h1ffd9; 
        10'b1100000101: data <= 17'h1ffc6; 
        10'b1100000110: data <= 17'h1ffdf; 
        10'b1100000111: data <= 17'h1ffd6; 
        10'b1100001000: data <= 17'h1fff4; 
        10'b1100001001: data <= 17'h1ff8c; 
        10'b1100001010: data <= 17'h1ffce; 
        10'b1100001011: data <= 17'h00004; 
        10'b1100001100: data <= 17'h1ff8c; 
        10'b1100001101: data <= 17'h1ffd4; 
        10'b1100001110: data <= 17'h1ffef; 
        10'b1100001111: data <= 17'h1ffc2; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 12) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 18'h3ff32; 
        10'b0000000001: data <= 18'h00005; 
        10'b0000000010: data <= 18'h3ff9a; 
        10'b0000000011: data <= 18'h3ff56; 
        10'b0000000100: data <= 18'h3ff97; 
        10'b0000000101: data <= 18'h3ff62; 
        10'b0000000110: data <= 18'h3ffbb; 
        10'b0000000111: data <= 18'h3ffc6; 
        10'b0000001000: data <= 18'h3ff2c; 
        10'b0000001001: data <= 18'h3ffaa; 
        10'b0000001010: data <= 18'h3ff3c; 
        10'b0000001011: data <= 18'h3ff7e; 
        10'b0000001100: data <= 18'h00027; 
        10'b0000001101: data <= 18'h00022; 
        10'b0000001110: data <= 18'h3ff37; 
        10'b0000001111: data <= 18'h3ffb8; 
        10'b0000010000: data <= 18'h3ff46; 
        10'b0000010001: data <= 18'h3ff48; 
        10'b0000010010: data <= 18'h00035; 
        10'b0000010011: data <= 18'h0000f; 
        10'b0000010100: data <= 18'h3ff67; 
        10'b0000010101: data <= 18'h3ffbf; 
        10'b0000010110: data <= 18'h3ff78; 
        10'b0000010111: data <= 18'h3ff20; 
        10'b0000011000: data <= 18'h3ff32; 
        10'b0000011001: data <= 18'h3ffb2; 
        10'b0000011010: data <= 18'h3fff6; 
        10'b0000011011: data <= 18'h3ffc8; 
        10'b0000011100: data <= 18'h3ffa9; 
        10'b0000011101: data <= 18'h3ff9b; 
        10'b0000011110: data <= 18'h00032; 
        10'b0000011111: data <= 18'h3ffcd; 
        10'b0000100000: data <= 18'h3ff3d; 
        10'b0000100001: data <= 18'h3ff36; 
        10'b0000100010: data <= 18'h3ff2f; 
        10'b0000100011: data <= 18'h3ff61; 
        10'b0000100100: data <= 18'h3ff63; 
        10'b0000100101: data <= 18'h3ffb7; 
        10'b0000100110: data <= 18'h00002; 
        10'b0000100111: data <= 18'h3ff44; 
        10'b0000101000: data <= 18'h3ff88; 
        10'b0000101001: data <= 18'h3ff3d; 
        10'b0000101010: data <= 18'h3ffbb; 
        10'b0000101011: data <= 18'h3ff20; 
        10'b0000101100: data <= 18'h3ffc5; 
        10'b0000101101: data <= 18'h3ff44; 
        10'b0000101110: data <= 18'h3ff82; 
        10'b0000101111: data <= 18'h3ff52; 
        10'b0000110000: data <= 18'h3ffb9; 
        10'b0000110001: data <= 18'h3ff49; 
        10'b0000110010: data <= 18'h3ff2a; 
        10'b0000110011: data <= 18'h3ff16; 
        10'b0000110100: data <= 18'h0000c; 
        10'b0000110101: data <= 18'h3ffcc; 
        10'b0000110110: data <= 18'h0000f; 
        10'b0000110111: data <= 18'h3ff73; 
        10'b0000111000: data <= 18'h3ff9c; 
        10'b0000111001: data <= 18'h3ff24; 
        10'b0000111010: data <= 18'h3ff38; 
        10'b0000111011: data <= 18'h3fffe; 
        10'b0000111100: data <= 18'h3ff2b; 
        10'b0000111101: data <= 18'h3ff3d; 
        10'b0000111110: data <= 18'h3ff92; 
        10'b0000111111: data <= 18'h3ffb2; 
        10'b0001000000: data <= 18'h3ffeb; 
        10'b0001000001: data <= 18'h3ff87; 
        10'b0001000010: data <= 18'h00074; 
        10'b0001000011: data <= 18'h0005f; 
        10'b0001000100: data <= 18'h00128; 
        10'b0001000101: data <= 18'h000ec; 
        10'b0001000110: data <= 18'h000d8; 
        10'b0001000111: data <= 18'h00056; 
        10'b0001001000: data <= 18'h00122; 
        10'b0001001001: data <= 18'h00063; 
        10'b0001001010: data <= 18'h00054; 
        10'b0001001011: data <= 18'h3ff6d; 
        10'b0001001100: data <= 18'h3fffc; 
        10'b0001001101: data <= 18'h3ffbc; 
        10'b0001001110: data <= 18'h3fed4; 
        10'b0001001111: data <= 18'h3ff96; 
        10'b0001010000: data <= 18'h3ffe0; 
        10'b0001010001: data <= 18'h00048; 
        10'b0001010010: data <= 18'h3ffaa; 
        10'b0001010011: data <= 18'h3ff86; 
        10'b0001010100: data <= 18'h3ff6e; 
        10'b0001010101: data <= 18'h3ff5a; 
        10'b0001010110: data <= 18'h3ffd0; 
        10'b0001010111: data <= 18'h3ff67; 
        10'b0001011000: data <= 18'h0002a; 
        10'b0001011001: data <= 18'h3ff46; 
        10'b0001011010: data <= 18'h3ffbc; 
        10'b0001011011: data <= 18'h00000; 
        10'b0001011100: data <= 18'h00035; 
        10'b0001011101: data <= 18'h001d7; 
        10'b0001011110: data <= 18'h002e1; 
        10'b0001011111: data <= 18'h002dc; 
        10'b0001100000: data <= 18'h002bd; 
        10'b0001100001: data <= 18'h00407; 
        10'b0001100010: data <= 18'h00232; 
        10'b0001100011: data <= 18'h000fa; 
        10'b0001100100: data <= 18'h001da; 
        10'b0001100101: data <= 18'h000d9; 
        10'b0001100110: data <= 18'h3ff33; 
        10'b0001100111: data <= 18'h3ffcd; 
        10'b0001101000: data <= 18'h3ff17; 
        10'b0001101001: data <= 18'h3feef; 
        10'b0001101010: data <= 18'h3feb2; 
        10'b0001101011: data <= 18'h3ff5a; 
        10'b0001101100: data <= 18'h00018; 
        10'b0001101101: data <= 18'h0004f; 
        10'b0001101110: data <= 18'h3ff48; 
        10'b0001101111: data <= 18'h3ffdb; 
        10'b0001110000: data <= 18'h3ff5f; 
        10'b0001110001: data <= 18'h3ff90; 
        10'b0001110010: data <= 18'h00038; 
        10'b0001110011: data <= 18'h3ff0f; 
        10'b0001110100: data <= 18'h3ff2b; 
        10'b0001110101: data <= 18'h3ffbc; 
        10'b0001110110: data <= 18'h0006d; 
        10'b0001110111: data <= 18'h00069; 
        10'b0001111000: data <= 18'h00130; 
        10'b0001111001: data <= 18'h00387; 
        10'b0001111010: data <= 18'h00390; 
        10'b0001111011: data <= 18'h0047a; 
        10'b0001111100: data <= 18'h003c8; 
        10'b0001111101: data <= 18'h00300; 
        10'b0001111110: data <= 18'h002ba; 
        10'b0001111111: data <= 18'h00134; 
        10'b0010000000: data <= 18'h0019c; 
        10'b0010000001: data <= 18'h0017d; 
        10'b0010000010: data <= 18'h3ff8e; 
        10'b0010000011: data <= 18'h3ff40; 
        10'b0010000100: data <= 18'h3ff6b; 
        10'b0010000101: data <= 18'h3fe3b; 
        10'b0010000110: data <= 18'h3fddc; 
        10'b0010000111: data <= 18'h3fdf1; 
        10'b0010001000: data <= 18'h3ffbc; 
        10'b0010001001: data <= 18'h3ffbc; 
        10'b0010001010: data <= 18'h3ff24; 
        10'b0010001011: data <= 18'h3ffd6; 
        10'b0010001100: data <= 18'h00013; 
        10'b0010001101: data <= 18'h3ffb8; 
        10'b0010001110: data <= 18'h3ff52; 
        10'b0010001111: data <= 18'h3ff18; 
        10'b0010010000: data <= 18'h3ff41; 
        10'b0010010001: data <= 18'h3ff5c; 
        10'b0010010010: data <= 18'h00065; 
        10'b0010010011: data <= 18'h001b9; 
        10'b0010010100: data <= 18'h00264; 
        10'b0010010101: data <= 18'h00417; 
        10'b0010010110: data <= 18'h00488; 
        10'b0010010111: data <= 18'h004ba; 
        10'b0010011000: data <= 18'h00454; 
        10'b0010011001: data <= 18'h004da; 
        10'b0010011010: data <= 18'h0047e; 
        10'b0010011011: data <= 18'h0042b; 
        10'b0010011100: data <= 18'h00485; 
        10'b0010011101: data <= 18'h003a8; 
        10'b0010011110: data <= 18'h002a4; 
        10'b0010011111: data <= 18'h3fee2; 
        10'b0010100000: data <= 18'h3feec; 
        10'b0010100001: data <= 18'h3fe3d; 
        10'b0010100010: data <= 18'h3fe36; 
        10'b0010100011: data <= 18'h3fd3a; 
        10'b0010100100: data <= 18'h3fecd; 
        10'b0010100101: data <= 18'h3ff52; 
        10'b0010100110: data <= 18'h0001c; 
        10'b0010100111: data <= 18'h3ff78; 
        10'b0010101000: data <= 18'h3ffa4; 
        10'b0010101001: data <= 18'h3ff5a; 
        10'b0010101010: data <= 18'h00025; 
        10'b0010101011: data <= 18'h3ffa7; 
        10'b0010101100: data <= 18'h3ff8b; 
        10'b0010101101: data <= 18'h0004a; 
        10'b0010101110: data <= 18'h001af; 
        10'b0010101111: data <= 18'h00343; 
        10'b0010110000: data <= 18'h0027e; 
        10'b0010110001: data <= 18'h002d5; 
        10'b0010110010: data <= 18'h003d5; 
        10'b0010110011: data <= 18'h00265; 
        10'b0010110100: data <= 18'h0028c; 
        10'b0010110101: data <= 18'h0034a; 
        10'b0010110110: data <= 18'h002e8; 
        10'b0010110111: data <= 18'h00195; 
        10'b0010111000: data <= 18'h001c0; 
        10'b0010111001: data <= 18'h00074; 
        10'b0010111010: data <= 18'h00055; 
        10'b0010111011: data <= 18'h3fef9; 
        10'b0010111100: data <= 18'h3ff51; 
        10'b0010111101: data <= 18'h3fdc3; 
        10'b0010111110: data <= 18'h3fdc7; 
        10'b0010111111: data <= 18'h3fce6; 
        10'b0011000000: data <= 18'h3fe27; 
        10'b0011000001: data <= 18'h3fef7; 
        10'b0011000010: data <= 18'h00022; 
        10'b0011000011: data <= 18'h3ffe5; 
        10'b0011000100: data <= 18'h3ff86; 
        10'b0011000101: data <= 18'h00018; 
        10'b0011000110: data <= 18'h0001b; 
        10'b0011000111: data <= 18'h3ff90; 
        10'b0011001000: data <= 18'h0000b; 
        10'b0011001001: data <= 18'h000e8; 
        10'b0011001010: data <= 18'h0022c; 
        10'b0011001011: data <= 18'h00325; 
        10'b0011001100: data <= 18'h00292; 
        10'b0011001101: data <= 18'h00266; 
        10'b0011001110: data <= 18'h000eb; 
        10'b0011001111: data <= 18'h00115; 
        10'b0011010000: data <= 18'h0002f; 
        10'b0011010001: data <= 18'h001af; 
        10'b0011010010: data <= 18'h00213; 
        10'b0011010011: data <= 18'h0006f; 
        10'b0011010100: data <= 18'h00047; 
        10'b0011010101: data <= 18'h3fd5f; 
        10'b0011010110: data <= 18'h3ff1c; 
        10'b0011010111: data <= 18'h3ff42; 
        10'b0011011000: data <= 18'h3ff29; 
        10'b0011011001: data <= 18'h3ff04; 
        10'b0011011010: data <= 18'h3ff44; 
        10'b0011011011: data <= 18'h3fd73; 
        10'b0011011100: data <= 18'h3fe3c; 
        10'b0011011101: data <= 18'h3ff76; 
        10'b0011011110: data <= 18'h3ff52; 
        10'b0011011111: data <= 18'h3ff2c; 
        10'b0011100000: data <= 18'h3ffcf; 
        10'b0011100001: data <= 18'h00020; 
        10'b0011100010: data <= 18'h3ffa6; 
        10'b0011100011: data <= 18'h0001d; 
        10'b0011100100: data <= 18'h00079; 
        10'b0011100101: data <= 18'h00178; 
        10'b0011100110: data <= 18'h00110; 
        10'b0011100111: data <= 18'h00180; 
        10'b0011101000: data <= 18'h00185; 
        10'b0011101001: data <= 18'h001b1; 
        10'b0011101010: data <= 18'h001b3; 
        10'b0011101011: data <= 18'h001f0; 
        10'b0011101100: data <= 18'h00127; 
        10'b0011101101: data <= 18'h00160; 
        10'b0011101110: data <= 18'h003a2; 
        10'b0011101111: data <= 18'h0020b; 
        10'b0011110000: data <= 18'h3ffc0; 
        10'b0011110001: data <= 18'h3ff01; 
        10'b0011110010: data <= 18'h3fff9; 
        10'b0011110011: data <= 18'h000ce; 
        10'b0011110100: data <= 18'h00005; 
        10'b0011110101: data <= 18'h3ff72; 
        10'b0011110110: data <= 18'h3fe85; 
        10'b0011110111: data <= 18'h3fd06; 
        10'b0011111000: data <= 18'h3fdb7; 
        10'b0011111001: data <= 18'h3ff0c; 
        10'b0011111010: data <= 18'h3ff8e; 
        10'b0011111011: data <= 18'h3ff45; 
        10'b0011111100: data <= 18'h3ff5f; 
        10'b0011111101: data <= 18'h3ffd9; 
        10'b0011111110: data <= 18'h3fff7; 
        10'b0011111111: data <= 18'h00061; 
        10'b0100000000: data <= 18'h000bd; 
        10'b0100000001: data <= 18'h001a5; 
        10'b0100000010: data <= 18'h00094; 
        10'b0100000011: data <= 18'h0001c; 
        10'b0100000100: data <= 18'h3ff6e; 
        10'b0100000101: data <= 18'h000e3; 
        10'b0100000110: data <= 18'h000b0; 
        10'b0100000111: data <= 18'h000e3; 
        10'b0100001000: data <= 18'h0003b; 
        10'b0100001001: data <= 18'h3ffe8; 
        10'b0100001010: data <= 18'h0025f; 
        10'b0100001011: data <= 18'h00290; 
        10'b0100001100: data <= 18'h000e2; 
        10'b0100001101: data <= 18'h00011; 
        10'b0100001110: data <= 18'h3ffc3; 
        10'b0100001111: data <= 18'h3fffb; 
        10'b0100010000: data <= 18'h3ffe4; 
        10'b0100010001: data <= 18'h3fff1; 
        10'b0100010010: data <= 18'h3ff0f; 
        10'b0100010011: data <= 18'h3fd78; 
        10'b0100010100: data <= 18'h3fdd7; 
        10'b0100010101: data <= 18'h3ff4c; 
        10'b0100010110: data <= 18'h0001d; 
        10'b0100010111: data <= 18'h3ff2f; 
        10'b0100011000: data <= 18'h00029; 
        10'b0100011001: data <= 18'h3ffd1; 
        10'b0100011010: data <= 18'h3ffa0; 
        10'b0100011011: data <= 18'h3ff78; 
        10'b0100011100: data <= 18'h0001d; 
        10'b0100011101: data <= 18'h3ff99; 
        10'b0100011110: data <= 18'h3ff2d; 
        10'b0100011111: data <= 18'h3fc01; 
        10'b0100100000: data <= 18'h3fc6d; 
        10'b0100100001: data <= 18'h3fd4d; 
        10'b0100100010: data <= 18'h3fbdf; 
        10'b0100100011: data <= 18'h3fb6c; 
        10'b0100100100: data <= 18'h3faac; 
        10'b0100100101: data <= 18'h3fa05; 
        10'b0100100110: data <= 18'h3fd7d; 
        10'b0100100111: data <= 18'h00075; 
        10'b0100101000: data <= 18'h000a6; 
        10'b0100101001: data <= 18'h0001c; 
        10'b0100101010: data <= 18'h00055; 
        10'b0100101011: data <= 18'h3ff84; 
        10'b0100101100: data <= 18'h3ffa5; 
        10'b0100101101: data <= 18'h3ff83; 
        10'b0100101110: data <= 18'h3febf; 
        10'b0100101111: data <= 18'h3fd17; 
        10'b0100110000: data <= 18'h3fe66; 
        10'b0100110001: data <= 18'h3ffef; 
        10'b0100110010: data <= 18'h3ffed; 
        10'b0100110011: data <= 18'h3ff54; 
        10'b0100110100: data <= 18'h3ff2b; 
        10'b0100110101: data <= 18'h00035; 
        10'b0100110110: data <= 18'h3ffea; 
        10'b0100110111: data <= 18'h3ff3c; 
        10'b0100111000: data <= 18'h3fe81; 
        10'b0100111001: data <= 18'h3fcba; 
        10'b0100111010: data <= 18'h3fa62; 
        10'b0100111011: data <= 18'h3f814; 
        10'b0100111100: data <= 18'h3f864; 
        10'b0100111101: data <= 18'h3f70a; 
        10'b0100111110: data <= 18'h3f703; 
        10'b0100111111: data <= 18'h3f7cc; 
        10'b0101000000: data <= 18'h3f74b; 
        10'b0101000001: data <= 18'h3f564; 
        10'b0101000010: data <= 18'h3f7d6; 
        10'b0101000011: data <= 18'h3fc19; 
        10'b0101000100: data <= 18'h3fea6; 
        10'b0101000101: data <= 18'h3fed6; 
        10'b0101000110: data <= 18'h3fee2; 
        10'b0101000111: data <= 18'h3ffc7; 
        10'b0101001000: data <= 18'h3ff54; 
        10'b0101001001: data <= 18'h3ff4c; 
        10'b0101001010: data <= 18'h3fe25; 
        10'b0101001011: data <= 18'h3febb; 
        10'b0101001100: data <= 18'h3ffc5; 
        10'b0101001101: data <= 18'h3ff90; 
        10'b0101001110: data <= 18'h3ff4e; 
        10'b0101001111: data <= 18'h3ffcf; 
        10'b0101010000: data <= 18'h3ffb6; 
        10'b0101010001: data <= 18'h3ffc3; 
        10'b0101010010: data <= 18'h00015; 
        10'b0101010011: data <= 18'h3ffa7; 
        10'b0101010100: data <= 18'h3fe63; 
        10'b0101010101: data <= 18'h3fb20; 
        10'b0101010110: data <= 18'h3f684; 
        10'b0101010111: data <= 18'h3f466; 
        10'b0101011000: data <= 18'h3f52d; 
        10'b0101011001: data <= 18'h3f5be; 
        10'b0101011010: data <= 18'h3f6a1; 
        10'b0101011011: data <= 18'h3f73b; 
        10'b0101011100: data <= 18'h3f741; 
        10'b0101011101: data <= 18'h3f6e6; 
        10'b0101011110: data <= 18'h3f887; 
        10'b0101011111: data <= 18'h3fb04; 
        10'b0101100000: data <= 18'h3fc94; 
        10'b0101100001: data <= 18'h3fced; 
        10'b0101100010: data <= 18'h3fe74; 
        10'b0101100011: data <= 18'h00002; 
        10'b0101100100: data <= 18'h3fff8; 
        10'b0101100101: data <= 18'h3ff22; 
        10'b0101100110: data <= 18'h3fe07; 
        10'b0101100111: data <= 18'h3fd00; 
        10'b0101101000: data <= 18'h3ffa2; 
        10'b0101101001: data <= 18'h3ff81; 
        10'b0101101010: data <= 18'h00039; 
        10'b0101101011: data <= 18'h3ffc3; 
        10'b0101101100: data <= 18'h3ff66; 
        10'b0101101101: data <= 18'h3ff9b; 
        10'b0101101110: data <= 18'h00035; 
        10'b0101101111: data <= 18'h3ff60; 
        10'b0101110000: data <= 18'h3fd64; 
        10'b0101110001: data <= 18'h3f9da; 
        10'b0101110010: data <= 18'h3f63f; 
        10'b0101110011: data <= 18'h3f70c; 
        10'b0101110100: data <= 18'h3f7a4; 
        10'b0101110101: data <= 18'h3fa41; 
        10'b0101110110: data <= 18'h3fbee; 
        10'b0101110111: data <= 18'h3fe18; 
        10'b0101111000: data <= 18'h3fcfc; 
        10'b0101111001: data <= 18'h3fea1; 
        10'b0101111010: data <= 18'h3fc8e; 
        10'b0101111011: data <= 18'h3fc7c; 
        10'b0101111100: data <= 18'h3fbd5; 
        10'b0101111101: data <= 18'h3fcfe; 
        10'b0101111110: data <= 18'h3fe58; 
        10'b0101111111: data <= 18'h3ffaf; 
        10'b0110000000: data <= 18'h3ff83; 
        10'b0110000001: data <= 18'h3feef; 
        10'b0110000010: data <= 18'h3fd85; 
        10'b0110000011: data <= 18'h3fdbe; 
        10'b0110000100: data <= 18'h3fedb; 
        10'b0110000101: data <= 18'h00049; 
        10'b0110000110: data <= 18'h3ff9e; 
        10'b0110000111: data <= 18'h3fffa; 
        10'b0110001000: data <= 18'h00021; 
        10'b0110001001: data <= 18'h3ffcb; 
        10'b0110001010: data <= 18'h00006; 
        10'b0110001011: data <= 18'h3ff79; 
        10'b0110001100: data <= 18'h3ff00; 
        10'b0110001101: data <= 18'h3fbd9; 
        10'b0110001110: data <= 18'h3fabf; 
        10'b0110001111: data <= 18'h3fbb8; 
        10'b0110010000: data <= 18'h3fe48; 
        10'b0110010001: data <= 18'h3ffb4; 
        10'b0110010010: data <= 18'h00112; 
        10'b0110010011: data <= 18'h0016b; 
        10'b0110010100: data <= 18'h001ae; 
        10'b0110010101: data <= 18'h0029e; 
        10'b0110010110: data <= 18'h0002e; 
        10'b0110010111: data <= 18'h3fe53; 
        10'b0110011000: data <= 18'h3fec1; 
        10'b0110011001: data <= 18'h3fdd8; 
        10'b0110011010: data <= 18'h3ffa3; 
        10'b0110011011: data <= 18'h3fe9d; 
        10'b0110011100: data <= 18'h3ff90; 
        10'b0110011101: data <= 18'h3fe67; 
        10'b0110011110: data <= 18'h3fd21; 
        10'b0110011111: data <= 18'h3fde9; 
        10'b0110100000: data <= 18'h3ff97; 
        10'b0110100001: data <= 18'h00104; 
        10'b0110100010: data <= 18'h00127; 
        10'b0110100011: data <= 18'h3ff5c; 
        10'b0110100100: data <= 18'h3ff8d; 
        10'b0110100101: data <= 18'h3ffa5; 
        10'b0110100110: data <= 18'h3ff89; 
        10'b0110100111: data <= 18'h000f3; 
        10'b0110101000: data <= 18'h00076; 
        10'b0110101001: data <= 18'h00035; 
        10'b0110101010: data <= 18'h00120; 
        10'b0110101011: data <= 18'h00151; 
        10'b0110101100: data <= 18'h00272; 
        10'b0110101101: data <= 18'h001ba; 
        10'b0110101110: data <= 18'h00212; 
        10'b0110101111: data <= 18'h00138; 
        10'b0110110000: data <= 18'h00114; 
        10'b0110110001: data <= 18'h00287; 
        10'b0110110010: data <= 18'h00030; 
        10'b0110110011: data <= 18'h000fe; 
        10'b0110110100: data <= 18'h00024; 
        10'b0110110101: data <= 18'h3fdff; 
        10'b0110110110: data <= 18'h3fe18; 
        10'b0110110111: data <= 18'h3fed4; 
        10'b0110111000: data <= 18'h3ff26; 
        10'b0110111001: data <= 18'h3feb6; 
        10'b0110111010: data <= 18'h3fd66; 
        10'b0110111011: data <= 18'h3fea9; 
        10'b0110111100: data <= 18'h000cd; 
        10'b0110111101: data <= 18'h0015d; 
        10'b0110111110: data <= 18'h000bd; 
        10'b0110111111: data <= 18'h3ff45; 
        10'b0111000000: data <= 18'h3ff71; 
        10'b0111000001: data <= 18'h3ff23; 
        10'b0111000010: data <= 18'h3ff05; 
        10'b0111000011: data <= 18'h00102; 
        10'b0111000100: data <= 18'h0021e; 
        10'b0111000101: data <= 18'h00375; 
        10'b0111000110: data <= 18'h00385; 
        10'b0111000111: data <= 18'h00218; 
        10'b0111001000: data <= 18'h000de; 
        10'b0111001001: data <= 18'h001cf; 
        10'b0111001010: data <= 18'h001ae; 
        10'b0111001011: data <= 18'h00188; 
        10'b0111001100: data <= 18'h00329; 
        10'b0111001101: data <= 18'h002c8; 
        10'b0111001110: data <= 18'h00095; 
        10'b0111001111: data <= 18'h3ffab; 
        10'b0111010000: data <= 18'h3fffd; 
        10'b0111010001: data <= 18'h3feb3; 
        10'b0111010010: data <= 18'h3fedc; 
        10'b0111010011: data <= 18'h3fe01; 
        10'b0111010100: data <= 18'h3ff4a; 
        10'b0111010101: data <= 18'h0001c; 
        10'b0111010110: data <= 18'h00070; 
        10'b0111010111: data <= 18'h000ee; 
        10'b0111011000: data <= 18'h002f3; 
        10'b0111011001: data <= 18'h003a7; 
        10'b0111011010: data <= 18'h0009d; 
        10'b0111011011: data <= 18'h3ff6e; 
        10'b0111011100: data <= 18'h3ff87; 
        10'b0111011101: data <= 18'h0002b; 
        10'b0111011110: data <= 18'h3ffa2; 
        10'b0111011111: data <= 18'h00139; 
        10'b0111100000: data <= 18'h0039e; 
        10'b0111100001: data <= 18'h0050a; 
        10'b0111100010: data <= 18'h0049b; 
        10'b0111100011: data <= 18'h00328; 
        10'b0111100100: data <= 18'h00232; 
        10'b0111100101: data <= 18'h002a9; 
        10'b0111100110: data <= 18'h00418; 
        10'b0111100111: data <= 18'h0035b; 
        10'b0111101000: data <= 18'h003d9; 
        10'b0111101001: data <= 18'h001cd; 
        10'b0111101010: data <= 18'h000ed; 
        10'b0111101011: data <= 18'h00140; 
        10'b0111101100: data <= 18'h00143; 
        10'b0111101101: data <= 18'h3ffce; 
        10'b0111101110: data <= 18'h000d2; 
        10'b0111101111: data <= 18'h3ff7a; 
        10'b0111110000: data <= 18'h00183; 
        10'b0111110001: data <= 18'h0019d; 
        10'b0111110010: data <= 18'h00133; 
        10'b0111110011: data <= 18'h001a9; 
        10'b0111110100: data <= 18'h004ba; 
        10'b0111110101: data <= 18'h00419; 
        10'b0111110110: data <= 18'h000f0; 
        10'b0111110111: data <= 18'h00020; 
        10'b0111111000: data <= 18'h3ffe5; 
        10'b0111111001: data <= 18'h3fff1; 
        10'b0111111010: data <= 18'h3fec1; 
        10'b0111111011: data <= 18'h00054; 
        10'b0111111100: data <= 18'h003eb; 
        10'b0111111101: data <= 18'h0069f; 
        10'b0111111110: data <= 18'h0063b; 
        10'b0111111111: data <= 18'h0047c; 
        10'b1000000000: data <= 18'h002fe; 
        10'b1000000001: data <= 18'h00353; 
        10'b1000000010: data <= 18'h00515; 
        10'b1000000011: data <= 18'h00497; 
        10'b1000000100: data <= 18'h00750; 
        10'b1000000101: data <= 18'h00556; 
        10'b1000000110: data <= 18'h004a9; 
        10'b1000000111: data <= 18'h00245; 
        10'b1000001000: data <= 18'h00190; 
        10'b1000001001: data <= 18'h002de; 
        10'b1000001010: data <= 18'h001da; 
        10'b1000001011: data <= 18'h00142; 
        10'b1000001100: data <= 18'h00362; 
        10'b1000001101: data <= 18'h0037f; 
        10'b1000001110: data <= 18'h003cf; 
        10'b1000001111: data <= 18'h00508; 
        10'b1000010000: data <= 18'h0063f; 
        10'b1000010001: data <= 18'h0039a; 
        10'b1000010010: data <= 18'h3ffa8; 
        10'b1000010011: data <= 18'h3ff42; 
        10'b1000010100: data <= 18'h3ff5e; 
        10'b1000010101: data <= 18'h3ff69; 
        10'b1000010110: data <= 18'h3ff22; 
        10'b1000010111: data <= 18'h3fffc; 
        10'b1000011000: data <= 18'h00227; 
        10'b1000011001: data <= 18'h00406; 
        10'b1000011010: data <= 18'h00515; 
        10'b1000011011: data <= 18'h00468; 
        10'b1000011100: data <= 18'h00411; 
        10'b1000011101: data <= 18'h0044e; 
        10'b1000011110: data <= 18'h0041f; 
        10'b1000011111: data <= 18'h00460; 
        10'b1000100000: data <= 18'h004e6; 
        10'b1000100001: data <= 18'h003c4; 
        10'b1000100010: data <= 18'h00270; 
        10'b1000100011: data <= 18'h00128; 
        10'b1000100100: data <= 18'h001cc; 
        10'b1000100101: data <= 18'h0031f; 
        10'b1000100110: data <= 18'h00182; 
        10'b1000100111: data <= 18'h00179; 
        10'b1000101000: data <= 18'h00283; 
        10'b1000101001: data <= 18'h00323; 
        10'b1000101010: data <= 18'h00419; 
        10'b1000101011: data <= 18'h00465; 
        10'b1000101100: data <= 18'h003c9; 
        10'b1000101101: data <= 18'h001fc; 
        10'b1000101110: data <= 18'h0002b; 
        10'b1000101111: data <= 18'h0000c; 
        10'b1000110000: data <= 18'h3ff37; 
        10'b1000110001: data <= 18'h3fff0; 
        10'b1000110010: data <= 18'h3ffca; 
        10'b1000110011: data <= 18'h3feec; 
        10'b1000110100: data <= 18'h001e9; 
        10'b1000110101: data <= 18'h0025c; 
        10'b1000110110: data <= 18'h003aa; 
        10'b1000110111: data <= 18'h00518; 
        10'b1000111000: data <= 18'h004d7; 
        10'b1000111001: data <= 18'h00335; 
        10'b1000111010: data <= 18'h00315; 
        10'b1000111011: data <= 18'h00529; 
        10'b1000111100: data <= 18'h002df; 
        10'b1000111101: data <= 18'h000f3; 
        10'b1000111110: data <= 18'h000a3; 
        10'b1000111111: data <= 18'h000c8; 
        10'b1001000000: data <= 18'h00103; 
        10'b1001000001: data <= 18'h0000c; 
        10'b1001000010: data <= 18'h0023b; 
        10'b1001000011: data <= 18'h0037c; 
        10'b1001000100: data <= 18'h0025d; 
        10'b1001000101: data <= 18'h0035d; 
        10'b1001000110: data <= 18'h004af; 
        10'b1001000111: data <= 18'h00410; 
        10'b1001001000: data <= 18'h002ed; 
        10'b1001001001: data <= 18'h00163; 
        10'b1001001010: data <= 18'h3fffb; 
        10'b1001001011: data <= 18'h3ffdf; 
        10'b1001001100: data <= 18'h3ffb1; 
        10'b1001001101: data <= 18'h3ff40; 
        10'b1001001110: data <= 18'h3ffde; 
        10'b1001001111: data <= 18'h3ff92; 
        10'b1001010000: data <= 18'h00066; 
        10'b1001010001: data <= 18'h00104; 
        10'b1001010010: data <= 18'h0028b; 
        10'b1001010011: data <= 18'h002db; 
        10'b1001010100: data <= 18'h00284; 
        10'b1001010101: data <= 18'h00324; 
        10'b1001010110: data <= 18'h002c7; 
        10'b1001010111: data <= 18'h002bb; 
        10'b1001011000: data <= 18'h00112; 
        10'b1001011001: data <= 18'h00083; 
        10'b1001011010: data <= 18'h3ffb9; 
        10'b1001011011: data <= 18'h0001e; 
        10'b1001011100: data <= 18'h0015b; 
        10'b1001011101: data <= 18'h0017d; 
        10'b1001011110: data <= 18'h00342; 
        10'b1001011111: data <= 18'h0036d; 
        10'b1001100000: data <= 18'h00181; 
        10'b1001100001: data <= 18'h0035c; 
        10'b1001100010: data <= 18'h00427; 
        10'b1001100011: data <= 18'h004bb; 
        10'b1001100100: data <= 18'h00255; 
        10'b1001100101: data <= 18'h000ed; 
        10'b1001100110: data <= 18'h00037; 
        10'b1001100111: data <= 18'h3ffe5; 
        10'b1001101000: data <= 18'h3ff36; 
        10'b1001101001: data <= 18'h3ffca; 
        10'b1001101010: data <= 18'h3ff52; 
        10'b1001101011: data <= 18'h00039; 
        10'b1001101100: data <= 18'h000cd; 
        10'b1001101101: data <= 18'h0004a; 
        10'b1001101110: data <= 18'h001bb; 
        10'b1001101111: data <= 18'h00184; 
        10'b1001110000: data <= 18'h0016a; 
        10'b1001110001: data <= 18'h001fd; 
        10'b1001110010: data <= 18'h001f9; 
        10'b1001110011: data <= 18'h00257; 
        10'b1001110100: data <= 18'h00041; 
        10'b1001110101: data <= 18'h3fe27; 
        10'b1001110110: data <= 18'h3fdac; 
        10'b1001110111: data <= 18'h3feaf; 
        10'b1001111000: data <= 18'h3fec2; 
        10'b1001111001: data <= 18'h000f7; 
        10'b1001111010: data <= 18'h00307; 
        10'b1001111011: data <= 18'h003de; 
        10'b1001111100: data <= 18'h00384; 
        10'b1001111101: data <= 18'h0035d; 
        10'b1001111110: data <= 18'h002ec; 
        10'b1001111111: data <= 18'h00339; 
        10'b1010000000: data <= 18'h00132; 
        10'b1010000001: data <= 18'h3ffde; 
        10'b1010000010: data <= 18'h3ffcc; 
        10'b1010000011: data <= 18'h3ff70; 
        10'b1010000100: data <= 18'h3ffcf; 
        10'b1010000101: data <= 18'h3ffd5; 
        10'b1010000110: data <= 18'h3ffa7; 
        10'b1010000111: data <= 18'h3ff98; 
        10'b1010001000: data <= 18'h3ff8c; 
        10'b1010001001: data <= 18'h3ff1a; 
        10'b1010001010: data <= 18'h3fee5; 
        10'b1010001011: data <= 18'h3ff0a; 
        10'b1010001100: data <= 18'h3fe6d; 
        10'b1010001101: data <= 18'h3ff14; 
        10'b1010001110: data <= 18'h3ff62; 
        10'b1010001111: data <= 18'h000cc; 
        10'b1010010000: data <= 18'h00013; 
        10'b1010010001: data <= 18'h3fec3; 
        10'b1010010010: data <= 18'h3fe53; 
        10'b1010010011: data <= 18'h3fdd0; 
        10'b1010010100: data <= 18'h3fda0; 
        10'b1010010101: data <= 18'h3fec3; 
        10'b1010010110: data <= 18'h0007c; 
        10'b1010010111: data <= 18'h00307; 
        10'b1010011000: data <= 18'h002a6; 
        10'b1010011001: data <= 18'h0033f; 
        10'b1010011010: data <= 18'h00254; 
        10'b1010011011: data <= 18'h000e4; 
        10'b1010011100: data <= 18'h0008a; 
        10'b1010011101: data <= 18'h00058; 
        10'b1010011110: data <= 18'h3ffed; 
        10'b1010011111: data <= 18'h3ff95; 
        10'b1010100000: data <= 18'h3ffb4; 
        10'b1010100001: data <= 18'h3ff63; 
        10'b1010100010: data <= 18'h3fff8; 
        10'b1010100011: data <= 18'h3ffe5; 
        10'b1010100100: data <= 18'h3ff5a; 
        10'b1010100101: data <= 18'h3fe4e; 
        10'b1010100110: data <= 18'h3fcba; 
        10'b1010100111: data <= 18'h3fd8d; 
        10'b1010101000: data <= 18'h3fd7b; 
        10'b1010101001: data <= 18'h3fd50; 
        10'b1010101010: data <= 18'h3fd55; 
        10'b1010101011: data <= 18'h3fdf5; 
        10'b1010101100: data <= 18'h3fdf1; 
        10'b1010101101: data <= 18'h3fee2; 
        10'b1010101110: data <= 18'h3fe8a; 
        10'b1010101111: data <= 18'h3fdeb; 
        10'b1010110000: data <= 18'h3fe06; 
        10'b1010110001: data <= 18'h3fe74; 
        10'b1010110010: data <= 18'h3fe1b; 
        10'b1010110011: data <= 18'h3fefa; 
        10'b1010110100: data <= 18'h3ff18; 
        10'b1010110101: data <= 18'h3ff1a; 
        10'b1010110110: data <= 18'h3ff79; 
        10'b1010110111: data <= 18'h3ff96; 
        10'b1010111000: data <= 18'h3fff0; 
        10'b1010111001: data <= 18'h00056; 
        10'b1010111010: data <= 18'h3ff4b; 
        10'b1010111011: data <= 18'h3ff50; 
        10'b1010111100: data <= 18'h3fff8; 
        10'b1010111101: data <= 18'h3ff1e; 
        10'b1010111110: data <= 18'h3ff8d; 
        10'b1010111111: data <= 18'h3ff75; 
        10'b1011000000: data <= 18'h3ff4d; 
        10'b1011000001: data <= 18'h3fece; 
        10'b1011000010: data <= 18'h3fe69; 
        10'b1011000011: data <= 18'h3fd95; 
        10'b1011000100: data <= 18'h3fd51; 
        10'b1011000101: data <= 18'h3fd83; 
        10'b1011000110: data <= 18'h3fdbf; 
        10'b1011000111: data <= 18'h3fd21; 
        10'b1011001000: data <= 18'h3fe14; 
        10'b1011001001: data <= 18'h3fe32; 
        10'b1011001010: data <= 18'h3fd9b; 
        10'b1011001011: data <= 18'h3fe07; 
        10'b1011001100: data <= 18'h3fe89; 
        10'b1011001101: data <= 18'h3fea1; 
        10'b1011001110: data <= 18'h3ff7a; 
        10'b1011001111: data <= 18'h3febf; 
        10'b1011010000: data <= 18'h3ff8d; 
        10'b1011010001: data <= 18'h3ff84; 
        10'b1011010010: data <= 18'h3fffb; 
        10'b1011010011: data <= 18'h3ff53; 
        10'b1011010100: data <= 18'h3ffbf; 
        10'b1011010101: data <= 18'h3ff57; 
        10'b1011010110: data <= 18'h3ff24; 
        10'b1011010111: data <= 18'h3ff5a; 
        10'b1011011000: data <= 18'h3ff2c; 
        10'b1011011001: data <= 18'h3ff7a; 
        10'b1011011010: data <= 18'h3ff9f; 
        10'b1011011011: data <= 18'h0000a; 
        10'b1011011100: data <= 18'h3ffdd; 
        10'b1011011101: data <= 18'h3ff96; 
        10'b1011011110: data <= 18'h3ffd5; 
        10'b1011011111: data <= 18'h3fff8; 
        10'b1011100000: data <= 18'h3ff91; 
        10'b1011100001: data <= 18'h0000d; 
        10'b1011100010: data <= 18'h3fffc; 
        10'b1011100011: data <= 18'h00007; 
        10'b1011100100: data <= 18'h00014; 
        10'b1011100101: data <= 18'h3ffbf; 
        10'b1011100110: data <= 18'h3ff6d; 
        10'b1011100111: data <= 18'h3ff10; 
        10'b1011101000: data <= 18'h3ff82; 
        10'b1011101001: data <= 18'h3ffbd; 
        10'b1011101010: data <= 18'h3ffb0; 
        10'b1011101011: data <= 18'h3ff55; 
        10'b1011101100: data <= 18'h00016; 
        10'b1011101101: data <= 18'h3fffc; 
        10'b1011101110: data <= 18'h3ff56; 
        10'b1011101111: data <= 18'h3ff7a; 
        10'b1011110000: data <= 18'h3ff29; 
        10'b1011110001: data <= 18'h0000a; 
        10'b1011110010: data <= 18'h00007; 
        10'b1011110011: data <= 18'h3fff5; 
        10'b1011110100: data <= 18'h3ffee; 
        10'b1011110101: data <= 18'h3ff64; 
        10'b1011110110: data <= 18'h3ff3d; 
        10'b1011110111: data <= 18'h3ffb3; 
        10'b1011111000: data <= 18'h3ff26; 
        10'b1011111001: data <= 18'h0002d; 
        10'b1011111010: data <= 18'h00029; 
        10'b1011111011: data <= 18'h3ff81; 
        10'b1011111100: data <= 18'h3fff3; 
        10'b1011111101: data <= 18'h3ff54; 
        10'b1011111110: data <= 18'h0001e; 
        10'b1011111111: data <= 18'h3ff20; 
        10'b1100000000: data <= 18'h3fff4; 
        10'b1100000001: data <= 18'h3ff94; 
        10'b1100000010: data <= 18'h3ffce; 
        10'b1100000011: data <= 18'h3ff42; 
        10'b1100000100: data <= 18'h3ffb2; 
        10'b1100000101: data <= 18'h3ff8b; 
        10'b1100000110: data <= 18'h3ffbd; 
        10'b1100000111: data <= 18'h3ffad; 
        10'b1100001000: data <= 18'h3ffe7; 
        10'b1100001001: data <= 18'h3ff18; 
        10'b1100001010: data <= 18'h3ff9c; 
        10'b1100001011: data <= 18'h00008; 
        10'b1100001100: data <= 18'h3ff18; 
        10'b1100001101: data <= 18'h3ffa8; 
        10'b1100001110: data <= 18'h3ffdf; 
        10'b1100001111: data <= 18'h3ff84; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 13) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 19'h7fe64; 
        10'b0000000001: data <= 19'h0000a; 
        10'b0000000010: data <= 19'h7ff33; 
        10'b0000000011: data <= 19'h7feac; 
        10'b0000000100: data <= 19'h7ff2d; 
        10'b0000000101: data <= 19'h7fec3; 
        10'b0000000110: data <= 19'h7ff75; 
        10'b0000000111: data <= 19'h7ff8b; 
        10'b0000001000: data <= 19'h7fe59; 
        10'b0000001001: data <= 19'h7ff54; 
        10'b0000001010: data <= 19'h7fe77; 
        10'b0000001011: data <= 19'h7fefb; 
        10'b0000001100: data <= 19'h0004f; 
        10'b0000001101: data <= 19'h00045; 
        10'b0000001110: data <= 19'h7fe6f; 
        10'b0000001111: data <= 19'h7ff6f; 
        10'b0000010000: data <= 19'h7fe8c; 
        10'b0000010001: data <= 19'h7fe90; 
        10'b0000010010: data <= 19'h0006b; 
        10'b0000010011: data <= 19'h0001e; 
        10'b0000010100: data <= 19'h7fece; 
        10'b0000010101: data <= 19'h7ff7d; 
        10'b0000010110: data <= 19'h7fef1; 
        10'b0000010111: data <= 19'h7fe40; 
        10'b0000011000: data <= 19'h7fe64; 
        10'b0000011001: data <= 19'h7ff65; 
        10'b0000011010: data <= 19'h7ffec; 
        10'b0000011011: data <= 19'h7ff8f; 
        10'b0000011100: data <= 19'h7ff52; 
        10'b0000011101: data <= 19'h7ff36; 
        10'b0000011110: data <= 19'h00064; 
        10'b0000011111: data <= 19'h7ff9a; 
        10'b0000100000: data <= 19'h7fe79; 
        10'b0000100001: data <= 19'h7fe6d; 
        10'b0000100010: data <= 19'h7fe5d; 
        10'b0000100011: data <= 19'h7fec2; 
        10'b0000100100: data <= 19'h7fec7; 
        10'b0000100101: data <= 19'h7ff6e; 
        10'b0000100110: data <= 19'h00004; 
        10'b0000100111: data <= 19'h7fe88; 
        10'b0000101000: data <= 19'h7ff0f; 
        10'b0000101001: data <= 19'h7fe7b; 
        10'b0000101010: data <= 19'h7ff76; 
        10'b0000101011: data <= 19'h7fe40; 
        10'b0000101100: data <= 19'h7ff89; 
        10'b0000101101: data <= 19'h7fe89; 
        10'b0000101110: data <= 19'h7ff04; 
        10'b0000101111: data <= 19'h7fea5; 
        10'b0000110000: data <= 19'h7ff72; 
        10'b0000110001: data <= 19'h7fe93; 
        10'b0000110010: data <= 19'h7fe54; 
        10'b0000110011: data <= 19'h7fe2b; 
        10'b0000110100: data <= 19'h00017; 
        10'b0000110101: data <= 19'h7ff98; 
        10'b0000110110: data <= 19'h0001e; 
        10'b0000110111: data <= 19'h7fee6; 
        10'b0000111000: data <= 19'h7ff38; 
        10'b0000111001: data <= 19'h7fe47; 
        10'b0000111010: data <= 19'h7fe70; 
        10'b0000111011: data <= 19'h7fffc; 
        10'b0000111100: data <= 19'h7fe56; 
        10'b0000111101: data <= 19'h7fe7a; 
        10'b0000111110: data <= 19'h7ff23; 
        10'b0000111111: data <= 19'h7ff65; 
        10'b0001000000: data <= 19'h7ffd6; 
        10'b0001000001: data <= 19'h7ff0e; 
        10'b0001000010: data <= 19'h000e7; 
        10'b0001000011: data <= 19'h000bf; 
        10'b0001000100: data <= 19'h0024f; 
        10'b0001000101: data <= 19'h001d8; 
        10'b0001000110: data <= 19'h001af; 
        10'b0001000111: data <= 19'h000ab; 
        10'b0001001000: data <= 19'h00245; 
        10'b0001001001: data <= 19'h000c6; 
        10'b0001001010: data <= 19'h000a8; 
        10'b0001001011: data <= 19'h7feda; 
        10'b0001001100: data <= 19'h7fff8; 
        10'b0001001101: data <= 19'h7ff77; 
        10'b0001001110: data <= 19'h7fda7; 
        10'b0001001111: data <= 19'h7ff2c; 
        10'b0001010000: data <= 19'h7ffc0; 
        10'b0001010001: data <= 19'h00091; 
        10'b0001010010: data <= 19'h7ff53; 
        10'b0001010011: data <= 19'h7ff0d; 
        10'b0001010100: data <= 19'h7fedb; 
        10'b0001010101: data <= 19'h7feb3; 
        10'b0001010110: data <= 19'h7ffa1; 
        10'b0001010111: data <= 19'h7fece; 
        10'b0001011000: data <= 19'h00053; 
        10'b0001011001: data <= 19'h7fe8d; 
        10'b0001011010: data <= 19'h7ff79; 
        10'b0001011011: data <= 19'h00000; 
        10'b0001011100: data <= 19'h0006a; 
        10'b0001011101: data <= 19'h003ae; 
        10'b0001011110: data <= 19'h005c2; 
        10'b0001011111: data <= 19'h005b8; 
        10'b0001100000: data <= 19'h00579; 
        10'b0001100001: data <= 19'h0080d; 
        10'b0001100010: data <= 19'h00465; 
        10'b0001100011: data <= 19'h001f3; 
        10'b0001100100: data <= 19'h003b4; 
        10'b0001100101: data <= 19'h001b2; 
        10'b0001100110: data <= 19'h7fe66; 
        10'b0001100111: data <= 19'h7ff9b; 
        10'b0001101000: data <= 19'h7fe2e; 
        10'b0001101001: data <= 19'h7fdde; 
        10'b0001101010: data <= 19'h7fd65; 
        10'b0001101011: data <= 19'h7feb5; 
        10'b0001101100: data <= 19'h00031; 
        10'b0001101101: data <= 19'h0009d; 
        10'b0001101110: data <= 19'h7fe8f; 
        10'b0001101111: data <= 19'h7ffb6; 
        10'b0001110000: data <= 19'h7febd; 
        10'b0001110001: data <= 19'h7ff20; 
        10'b0001110010: data <= 19'h00071; 
        10'b0001110011: data <= 19'h7fe1e; 
        10'b0001110100: data <= 19'h7fe57; 
        10'b0001110101: data <= 19'h7ff79; 
        10'b0001110110: data <= 19'h000da; 
        10'b0001110111: data <= 19'h000d3; 
        10'b0001111000: data <= 19'h0025f; 
        10'b0001111001: data <= 19'h0070d; 
        10'b0001111010: data <= 19'h00720; 
        10'b0001111011: data <= 19'h008f3; 
        10'b0001111100: data <= 19'h00790; 
        10'b0001111101: data <= 19'h00600; 
        10'b0001111110: data <= 19'h00574; 
        10'b0001111111: data <= 19'h00269; 
        10'b0010000000: data <= 19'h00339; 
        10'b0010000001: data <= 19'h002fb; 
        10'b0010000010: data <= 19'h7ff1b; 
        10'b0010000011: data <= 19'h7fe7f; 
        10'b0010000100: data <= 19'h7fed7; 
        10'b0010000101: data <= 19'h7fc76; 
        10'b0010000110: data <= 19'h7fbb7; 
        10'b0010000111: data <= 19'h7fbe2; 
        10'b0010001000: data <= 19'h7ff79; 
        10'b0010001001: data <= 19'h7ff79; 
        10'b0010001010: data <= 19'h7fe47; 
        10'b0010001011: data <= 19'h7ffad; 
        10'b0010001100: data <= 19'h00026; 
        10'b0010001101: data <= 19'h7ff71; 
        10'b0010001110: data <= 19'h7fea4; 
        10'b0010001111: data <= 19'h7fe2f; 
        10'b0010010000: data <= 19'h7fe82; 
        10'b0010010001: data <= 19'h7feb8; 
        10'b0010010010: data <= 19'h000ca; 
        10'b0010010011: data <= 19'h00372; 
        10'b0010010100: data <= 19'h004c7; 
        10'b0010010101: data <= 19'h0082e; 
        10'b0010010110: data <= 19'h00910; 
        10'b0010010111: data <= 19'h00973; 
        10'b0010011000: data <= 19'h008a8; 
        10'b0010011001: data <= 19'h009b5; 
        10'b0010011010: data <= 19'h008fc; 
        10'b0010011011: data <= 19'h00856; 
        10'b0010011100: data <= 19'h0090a; 
        10'b0010011101: data <= 19'h00750; 
        10'b0010011110: data <= 19'h00549; 
        10'b0010011111: data <= 19'h7fdc5; 
        10'b0010100000: data <= 19'h7fdd8; 
        10'b0010100001: data <= 19'h7fc7b; 
        10'b0010100010: data <= 19'h7fc6c; 
        10'b0010100011: data <= 19'h7fa73; 
        10'b0010100100: data <= 19'h7fd9b; 
        10'b0010100101: data <= 19'h7fea3; 
        10'b0010100110: data <= 19'h00038; 
        10'b0010100111: data <= 19'h7fef1; 
        10'b0010101000: data <= 19'h7ff47; 
        10'b0010101001: data <= 19'h7feb5; 
        10'b0010101010: data <= 19'h0004b; 
        10'b0010101011: data <= 19'h7ff4e; 
        10'b0010101100: data <= 19'h7ff17; 
        10'b0010101101: data <= 19'h00094; 
        10'b0010101110: data <= 19'h0035f; 
        10'b0010101111: data <= 19'h00686; 
        10'b0010110000: data <= 19'h004fc; 
        10'b0010110001: data <= 19'h005a9; 
        10'b0010110010: data <= 19'h007aa; 
        10'b0010110011: data <= 19'h004cb; 
        10'b0010110100: data <= 19'h00518; 
        10'b0010110101: data <= 19'h00694; 
        10'b0010110110: data <= 19'h005cf; 
        10'b0010110111: data <= 19'h00329; 
        10'b0010111000: data <= 19'h0037f; 
        10'b0010111001: data <= 19'h000e7; 
        10'b0010111010: data <= 19'h000ab; 
        10'b0010111011: data <= 19'h7fdf2; 
        10'b0010111100: data <= 19'h7fea2; 
        10'b0010111101: data <= 19'h7fb86; 
        10'b0010111110: data <= 19'h7fb8e; 
        10'b0010111111: data <= 19'h7f9cd; 
        10'b0011000000: data <= 19'h7fc4f; 
        10'b0011000001: data <= 19'h7fdee; 
        10'b0011000010: data <= 19'h00043; 
        10'b0011000011: data <= 19'h7ffca; 
        10'b0011000100: data <= 19'h7ff0b; 
        10'b0011000101: data <= 19'h00031; 
        10'b0011000110: data <= 19'h00035; 
        10'b0011000111: data <= 19'h7ff20; 
        10'b0011001000: data <= 19'h00016; 
        10'b0011001001: data <= 19'h001d0; 
        10'b0011001010: data <= 19'h00458; 
        10'b0011001011: data <= 19'h00649; 
        10'b0011001100: data <= 19'h00525; 
        10'b0011001101: data <= 19'h004cd; 
        10'b0011001110: data <= 19'h001d5; 
        10'b0011001111: data <= 19'h0022b; 
        10'b0011010000: data <= 19'h0005f; 
        10'b0011010001: data <= 19'h0035e; 
        10'b0011010010: data <= 19'h00426; 
        10'b0011010011: data <= 19'h000df; 
        10'b0011010100: data <= 19'h0008f; 
        10'b0011010101: data <= 19'h7fabe; 
        10'b0011010110: data <= 19'h7fe38; 
        10'b0011010111: data <= 19'h7fe84; 
        10'b0011011000: data <= 19'h7fe51; 
        10'b0011011001: data <= 19'h7fe08; 
        10'b0011011010: data <= 19'h7fe88; 
        10'b0011011011: data <= 19'h7fae6; 
        10'b0011011100: data <= 19'h7fc77; 
        10'b0011011101: data <= 19'h7feec; 
        10'b0011011110: data <= 19'h7fea4; 
        10'b0011011111: data <= 19'h7fe58; 
        10'b0011100000: data <= 19'h7ff9f; 
        10'b0011100001: data <= 19'h00040; 
        10'b0011100010: data <= 19'h7ff4b; 
        10'b0011100011: data <= 19'h0003b; 
        10'b0011100100: data <= 19'h000f3; 
        10'b0011100101: data <= 19'h002f0; 
        10'b0011100110: data <= 19'h00220; 
        10'b0011100111: data <= 19'h00300; 
        10'b0011101000: data <= 19'h0030a; 
        10'b0011101001: data <= 19'h00362; 
        10'b0011101010: data <= 19'h00366; 
        10'b0011101011: data <= 19'h003e1; 
        10'b0011101100: data <= 19'h0024e; 
        10'b0011101101: data <= 19'h002c1; 
        10'b0011101110: data <= 19'h00744; 
        10'b0011101111: data <= 19'h00416; 
        10'b0011110000: data <= 19'h7ff7f; 
        10'b0011110001: data <= 19'h7fe02; 
        10'b0011110010: data <= 19'h7fff3; 
        10'b0011110011: data <= 19'h0019d; 
        10'b0011110100: data <= 19'h0000a; 
        10'b0011110101: data <= 19'h7fee3; 
        10'b0011110110: data <= 19'h7fd0a; 
        10'b0011110111: data <= 19'h7fa0c; 
        10'b0011111000: data <= 19'h7fb6f; 
        10'b0011111001: data <= 19'h7fe19; 
        10'b0011111010: data <= 19'h7ff1c; 
        10'b0011111011: data <= 19'h7fe8a; 
        10'b0011111100: data <= 19'h7febe; 
        10'b0011111101: data <= 19'h7ffb1; 
        10'b0011111110: data <= 19'h7ffef; 
        10'b0011111111: data <= 19'h000c3; 
        10'b0100000000: data <= 19'h0017a; 
        10'b0100000001: data <= 19'h0034b; 
        10'b0100000010: data <= 19'h00127; 
        10'b0100000011: data <= 19'h00039; 
        10'b0100000100: data <= 19'h7fedd; 
        10'b0100000101: data <= 19'h001c5; 
        10'b0100000110: data <= 19'h00160; 
        10'b0100000111: data <= 19'h001c7; 
        10'b0100001000: data <= 19'h00076; 
        10'b0100001001: data <= 19'h7ffd1; 
        10'b0100001010: data <= 19'h004bd; 
        10'b0100001011: data <= 19'h00520; 
        10'b0100001100: data <= 19'h001c5; 
        10'b0100001101: data <= 19'h00022; 
        10'b0100001110: data <= 19'h7ff86; 
        10'b0100001111: data <= 19'h7fff5; 
        10'b0100010000: data <= 19'h7ffc9; 
        10'b0100010001: data <= 19'h7ffe3; 
        10'b0100010010: data <= 19'h7fe1e; 
        10'b0100010011: data <= 19'h7faf0; 
        10'b0100010100: data <= 19'h7fbae; 
        10'b0100010101: data <= 19'h7fe98; 
        10'b0100010110: data <= 19'h00039; 
        10'b0100010111: data <= 19'h7fe5e; 
        10'b0100011000: data <= 19'h00051; 
        10'b0100011001: data <= 19'h7ffa1; 
        10'b0100011010: data <= 19'h7ff40; 
        10'b0100011011: data <= 19'h7fef0; 
        10'b0100011100: data <= 19'h0003a; 
        10'b0100011101: data <= 19'h7ff32; 
        10'b0100011110: data <= 19'h7fe5b; 
        10'b0100011111: data <= 19'h7f802; 
        10'b0100100000: data <= 19'h7f8da; 
        10'b0100100001: data <= 19'h7fa99; 
        10'b0100100010: data <= 19'h7f7be; 
        10'b0100100011: data <= 19'h7f6d8; 
        10'b0100100100: data <= 19'h7f559; 
        10'b0100100101: data <= 19'h7f409; 
        10'b0100100110: data <= 19'h7fafa; 
        10'b0100100111: data <= 19'h000e9; 
        10'b0100101000: data <= 19'h0014b; 
        10'b0100101001: data <= 19'h00038; 
        10'b0100101010: data <= 19'h000aa; 
        10'b0100101011: data <= 19'h7ff07; 
        10'b0100101100: data <= 19'h7ff4b; 
        10'b0100101101: data <= 19'h7ff06; 
        10'b0100101110: data <= 19'h7fd7e; 
        10'b0100101111: data <= 19'h7fa2d; 
        10'b0100110000: data <= 19'h7fccd; 
        10'b0100110001: data <= 19'h7ffdd; 
        10'b0100110010: data <= 19'h7ffda; 
        10'b0100110011: data <= 19'h7fea8; 
        10'b0100110100: data <= 19'h7fe56; 
        10'b0100110101: data <= 19'h00069; 
        10'b0100110110: data <= 19'h7ffd5; 
        10'b0100110111: data <= 19'h7fe78; 
        10'b0100111000: data <= 19'h7fd01; 
        10'b0100111001: data <= 19'h7f974; 
        10'b0100111010: data <= 19'h7f4c3; 
        10'b0100111011: data <= 19'h7f028; 
        10'b0100111100: data <= 19'h7f0c8; 
        10'b0100111101: data <= 19'h7ee13; 
        10'b0100111110: data <= 19'h7ee06; 
        10'b0100111111: data <= 19'h7ef98; 
        10'b0101000000: data <= 19'h7ee95; 
        10'b0101000001: data <= 19'h7eac7; 
        10'b0101000010: data <= 19'h7efad; 
        10'b0101000011: data <= 19'h7f831; 
        10'b0101000100: data <= 19'h7fd4b; 
        10'b0101000101: data <= 19'h7fdac; 
        10'b0101000110: data <= 19'h7fdc3; 
        10'b0101000111: data <= 19'h7ff8d; 
        10'b0101001000: data <= 19'h7fea8; 
        10'b0101001001: data <= 19'h7fe99; 
        10'b0101001010: data <= 19'h7fc4a; 
        10'b0101001011: data <= 19'h7fd76; 
        10'b0101001100: data <= 19'h7ff8a; 
        10'b0101001101: data <= 19'h7ff1f; 
        10'b0101001110: data <= 19'h7fe9d; 
        10'b0101001111: data <= 19'h7ff9d; 
        10'b0101010000: data <= 19'h7ff6c; 
        10'b0101010001: data <= 19'h7ff86; 
        10'b0101010010: data <= 19'h0002b; 
        10'b0101010011: data <= 19'h7ff4d; 
        10'b0101010100: data <= 19'h7fcc6; 
        10'b0101010101: data <= 19'h7f640; 
        10'b0101010110: data <= 19'h7ed09; 
        10'b0101010111: data <= 19'h7e8cb; 
        10'b0101011000: data <= 19'h7ea5b; 
        10'b0101011001: data <= 19'h7eb7d; 
        10'b0101011010: data <= 19'h7ed41; 
        10'b0101011011: data <= 19'h7ee75; 
        10'b0101011100: data <= 19'h7ee82; 
        10'b0101011101: data <= 19'h7edcd; 
        10'b0101011110: data <= 19'h7f10d; 
        10'b0101011111: data <= 19'h7f608; 
        10'b0101100000: data <= 19'h7f929; 
        10'b0101100001: data <= 19'h7f9db; 
        10'b0101100010: data <= 19'h7fce7; 
        10'b0101100011: data <= 19'h00003; 
        10'b0101100100: data <= 19'h7fff1; 
        10'b0101100101: data <= 19'h7fe43; 
        10'b0101100110: data <= 19'h7fc0d; 
        10'b0101100111: data <= 19'h7f9ff; 
        10'b0101101000: data <= 19'h7ff45; 
        10'b0101101001: data <= 19'h7ff01; 
        10'b0101101010: data <= 19'h00072; 
        10'b0101101011: data <= 19'h7ff86; 
        10'b0101101100: data <= 19'h7fecb; 
        10'b0101101101: data <= 19'h7ff36; 
        10'b0101101110: data <= 19'h0006a; 
        10'b0101101111: data <= 19'h7fec1; 
        10'b0101110000: data <= 19'h7fac7; 
        10'b0101110001: data <= 19'h7f3b5; 
        10'b0101110010: data <= 19'h7ec7d; 
        10'b0101110011: data <= 19'h7ee17; 
        10'b0101110100: data <= 19'h7ef49; 
        10'b0101110101: data <= 19'h7f483; 
        10'b0101110110: data <= 19'h7f7dc; 
        10'b0101110111: data <= 19'h7fc30; 
        10'b0101111000: data <= 19'h7f9f8; 
        10'b0101111001: data <= 19'h7fd42; 
        10'b0101111010: data <= 19'h7f91d; 
        10'b0101111011: data <= 19'h7f8f9; 
        10'b0101111100: data <= 19'h7f7aa; 
        10'b0101111101: data <= 19'h7f9fb; 
        10'b0101111110: data <= 19'h7fcaf; 
        10'b0101111111: data <= 19'h7ff5d; 
        10'b0110000000: data <= 19'h7ff07; 
        10'b0110000001: data <= 19'h7fddd; 
        10'b0110000010: data <= 19'h7fb09; 
        10'b0110000011: data <= 19'h7fb7b; 
        10'b0110000100: data <= 19'h7fdb7; 
        10'b0110000101: data <= 19'h00093; 
        10'b0110000110: data <= 19'h7ff3d; 
        10'b0110000111: data <= 19'h7fff3; 
        10'b0110001000: data <= 19'h00043; 
        10'b0110001001: data <= 19'h7ff96; 
        10'b0110001010: data <= 19'h0000b; 
        10'b0110001011: data <= 19'h7fef3; 
        10'b0110001100: data <= 19'h7fe00; 
        10'b0110001101: data <= 19'h7f7b2; 
        10'b0110001110: data <= 19'h7f57f; 
        10'b0110001111: data <= 19'h7f76f; 
        10'b0110010000: data <= 19'h7fc91; 
        10'b0110010001: data <= 19'h7ff68; 
        10'b0110010010: data <= 19'h00224; 
        10'b0110010011: data <= 19'h002d6; 
        10'b0110010100: data <= 19'h0035d; 
        10'b0110010101: data <= 19'h0053b; 
        10'b0110010110: data <= 19'h0005b; 
        10'b0110010111: data <= 19'h7fca6; 
        10'b0110011000: data <= 19'h7fd83; 
        10'b0110011001: data <= 19'h7fbb0; 
        10'b0110011010: data <= 19'h7ff46; 
        10'b0110011011: data <= 19'h7fd3a; 
        10'b0110011100: data <= 19'h7ff1f; 
        10'b0110011101: data <= 19'h7fcce; 
        10'b0110011110: data <= 19'h7fa41; 
        10'b0110011111: data <= 19'h7fbd3; 
        10'b0110100000: data <= 19'h7ff2f; 
        10'b0110100001: data <= 19'h00209; 
        10'b0110100010: data <= 19'h0024f; 
        10'b0110100011: data <= 19'h7feb8; 
        10'b0110100100: data <= 19'h7ff1a; 
        10'b0110100101: data <= 19'h7ff4a; 
        10'b0110100110: data <= 19'h7ff13; 
        10'b0110100111: data <= 19'h001e6; 
        10'b0110101000: data <= 19'h000eb; 
        10'b0110101001: data <= 19'h0006a; 
        10'b0110101010: data <= 19'h0023f; 
        10'b0110101011: data <= 19'h002a2; 
        10'b0110101100: data <= 19'h004e4; 
        10'b0110101101: data <= 19'h00374; 
        10'b0110101110: data <= 19'h00425; 
        10'b0110101111: data <= 19'h0026f; 
        10'b0110110000: data <= 19'h00228; 
        10'b0110110001: data <= 19'h0050e; 
        10'b0110110010: data <= 19'h00060; 
        10'b0110110011: data <= 19'h001fc; 
        10'b0110110100: data <= 19'h00049; 
        10'b0110110101: data <= 19'h7fbfe; 
        10'b0110110110: data <= 19'h7fc2f; 
        10'b0110110111: data <= 19'h7fda9; 
        10'b0110111000: data <= 19'h7fe4b; 
        10'b0110111001: data <= 19'h7fd6c; 
        10'b0110111010: data <= 19'h7facc; 
        10'b0110111011: data <= 19'h7fd52; 
        10'b0110111100: data <= 19'h0019a; 
        10'b0110111101: data <= 19'h002ba; 
        10'b0110111110: data <= 19'h00179; 
        10'b0110111111: data <= 19'h7fe8b; 
        10'b0111000000: data <= 19'h7fee3; 
        10'b0111000001: data <= 19'h7fe45; 
        10'b0111000010: data <= 19'h7fe0a; 
        10'b0111000011: data <= 19'h00205; 
        10'b0111000100: data <= 19'h0043c; 
        10'b0111000101: data <= 19'h006ea; 
        10'b0111000110: data <= 19'h0070b; 
        10'b0111000111: data <= 19'h00431; 
        10'b0111001000: data <= 19'h001bd; 
        10'b0111001001: data <= 19'h0039d; 
        10'b0111001010: data <= 19'h0035c; 
        10'b0111001011: data <= 19'h00311; 
        10'b0111001100: data <= 19'h00651; 
        10'b0111001101: data <= 19'h00590; 
        10'b0111001110: data <= 19'h0012b; 
        10'b0111001111: data <= 19'h7ff56; 
        10'b0111010000: data <= 19'h7fffa; 
        10'b0111010001: data <= 19'h7fd65; 
        10'b0111010010: data <= 19'h7fdb9; 
        10'b0111010011: data <= 19'h7fc01; 
        10'b0111010100: data <= 19'h7fe94; 
        10'b0111010101: data <= 19'h00037; 
        10'b0111010110: data <= 19'h000e1; 
        10'b0111010111: data <= 19'h001db; 
        10'b0111011000: data <= 19'h005e6; 
        10'b0111011001: data <= 19'h0074f; 
        10'b0111011010: data <= 19'h00139; 
        10'b0111011011: data <= 19'h7fedb; 
        10'b0111011100: data <= 19'h7ff0e; 
        10'b0111011101: data <= 19'h00055; 
        10'b0111011110: data <= 19'h7ff44; 
        10'b0111011111: data <= 19'h00273; 
        10'b0111100000: data <= 19'h0073b; 
        10'b0111100001: data <= 19'h00a13; 
        10'b0111100010: data <= 19'h00935; 
        10'b0111100011: data <= 19'h0064f; 
        10'b0111100100: data <= 19'h00464; 
        10'b0111100101: data <= 19'h00553; 
        10'b0111100110: data <= 19'h00830; 
        10'b0111100111: data <= 19'h006b6; 
        10'b0111101000: data <= 19'h007b2; 
        10'b0111101001: data <= 19'h0039a; 
        10'b0111101010: data <= 19'h001db; 
        10'b0111101011: data <= 19'h00280; 
        10'b0111101100: data <= 19'h00287; 
        10'b0111101101: data <= 19'h7ff9c; 
        10'b0111101110: data <= 19'h001a3; 
        10'b0111101111: data <= 19'h7fef4; 
        10'b0111110000: data <= 19'h00306; 
        10'b0111110001: data <= 19'h00339; 
        10'b0111110010: data <= 19'h00265; 
        10'b0111110011: data <= 19'h00352; 
        10'b0111110100: data <= 19'h00974; 
        10'b0111110101: data <= 19'h00833; 
        10'b0111110110: data <= 19'h001df; 
        10'b0111110111: data <= 19'h00040; 
        10'b0111111000: data <= 19'h7ffc9; 
        10'b0111111001: data <= 19'h7ffe2; 
        10'b0111111010: data <= 19'h7fd83; 
        10'b0111111011: data <= 19'h000a9; 
        10'b0111111100: data <= 19'h007d6; 
        10'b0111111101: data <= 19'h00d3f; 
        10'b0111111110: data <= 19'h00c75; 
        10'b0111111111: data <= 19'h008f8; 
        10'b1000000000: data <= 19'h005fb; 
        10'b1000000001: data <= 19'h006a6; 
        10'b1000000010: data <= 19'h00a2a; 
        10'b1000000011: data <= 19'h0092f; 
        10'b1000000100: data <= 19'h00ea0; 
        10'b1000000101: data <= 19'h00aad; 
        10'b1000000110: data <= 19'h00953; 
        10'b1000000111: data <= 19'h00489; 
        10'b1000001000: data <= 19'h0031f; 
        10'b1000001001: data <= 19'h005bc; 
        10'b1000001010: data <= 19'h003b3; 
        10'b1000001011: data <= 19'h00285; 
        10'b1000001100: data <= 19'h006c4; 
        10'b1000001101: data <= 19'h006fd; 
        10'b1000001110: data <= 19'h0079e; 
        10'b1000001111: data <= 19'h00a11; 
        10'b1000010000: data <= 19'h00c7e; 
        10'b1000010001: data <= 19'h00734; 
        10'b1000010010: data <= 19'h7ff4f; 
        10'b1000010011: data <= 19'h7fe84; 
        10'b1000010100: data <= 19'h7febc; 
        10'b1000010101: data <= 19'h7fed2; 
        10'b1000010110: data <= 19'h7fe43; 
        10'b1000010111: data <= 19'h7fff9; 
        10'b1000011000: data <= 19'h0044e; 
        10'b1000011001: data <= 19'h0080c; 
        10'b1000011010: data <= 19'h00a29; 
        10'b1000011011: data <= 19'h008cf; 
        10'b1000011100: data <= 19'h00822; 
        10'b1000011101: data <= 19'h0089c; 
        10'b1000011110: data <= 19'h0083d; 
        10'b1000011111: data <= 19'h008c0; 
        10'b1000100000: data <= 19'h009cb; 
        10'b1000100001: data <= 19'h00788; 
        10'b1000100010: data <= 19'h004e1; 
        10'b1000100011: data <= 19'h00250; 
        10'b1000100100: data <= 19'h00398; 
        10'b1000100101: data <= 19'h0063d; 
        10'b1000100110: data <= 19'h00304; 
        10'b1000100111: data <= 19'h002f2; 
        10'b1000101000: data <= 19'h00507; 
        10'b1000101001: data <= 19'h00646; 
        10'b1000101010: data <= 19'h00831; 
        10'b1000101011: data <= 19'h008c9; 
        10'b1000101100: data <= 19'h00793; 
        10'b1000101101: data <= 19'h003f7; 
        10'b1000101110: data <= 19'h00056; 
        10'b1000101111: data <= 19'h00017; 
        10'b1000110000: data <= 19'h7fe6e; 
        10'b1000110001: data <= 19'h7ffe1; 
        10'b1000110010: data <= 19'h7ff95; 
        10'b1000110011: data <= 19'h7fdd8; 
        10'b1000110100: data <= 19'h003d2; 
        10'b1000110101: data <= 19'h004b8; 
        10'b1000110110: data <= 19'h00754; 
        10'b1000110111: data <= 19'h00a31; 
        10'b1000111000: data <= 19'h009ae; 
        10'b1000111001: data <= 19'h0066a; 
        10'b1000111010: data <= 19'h0062b; 
        10'b1000111011: data <= 19'h00a52; 
        10'b1000111100: data <= 19'h005bd; 
        10'b1000111101: data <= 19'h001e6; 
        10'b1000111110: data <= 19'h00146; 
        10'b1000111111: data <= 19'h00190; 
        10'b1001000000: data <= 19'h00206; 
        10'b1001000001: data <= 19'h00017; 
        10'b1001000010: data <= 19'h00476; 
        10'b1001000011: data <= 19'h006f8; 
        10'b1001000100: data <= 19'h004ba; 
        10'b1001000101: data <= 19'h006ba; 
        10'b1001000110: data <= 19'h0095e; 
        10'b1001000111: data <= 19'h00820; 
        10'b1001001000: data <= 19'h005d9; 
        10'b1001001001: data <= 19'h002c6; 
        10'b1001001010: data <= 19'h7fff7; 
        10'b1001001011: data <= 19'h7ffbe; 
        10'b1001001100: data <= 19'h7ff63; 
        10'b1001001101: data <= 19'h7fe81; 
        10'b1001001110: data <= 19'h7ffbb; 
        10'b1001001111: data <= 19'h7ff23; 
        10'b1001010000: data <= 19'h000cd; 
        10'b1001010001: data <= 19'h00208; 
        10'b1001010010: data <= 19'h00515; 
        10'b1001010011: data <= 19'h005b6; 
        10'b1001010100: data <= 19'h00509; 
        10'b1001010101: data <= 19'h00648; 
        10'b1001010110: data <= 19'h0058f; 
        10'b1001010111: data <= 19'h00575; 
        10'b1001011000: data <= 19'h00225; 
        10'b1001011001: data <= 19'h00105; 
        10'b1001011010: data <= 19'h7ff72; 
        10'b1001011011: data <= 19'h0003d; 
        10'b1001011100: data <= 19'h002b7; 
        10'b1001011101: data <= 19'h002f9; 
        10'b1001011110: data <= 19'h00684; 
        10'b1001011111: data <= 19'h006db; 
        10'b1001100000: data <= 19'h00302; 
        10'b1001100001: data <= 19'h006b9; 
        10'b1001100010: data <= 19'h0084e; 
        10'b1001100011: data <= 19'h00976; 
        10'b1001100100: data <= 19'h004a9; 
        10'b1001100101: data <= 19'h001d9; 
        10'b1001100110: data <= 19'h0006d; 
        10'b1001100111: data <= 19'h7ffcb; 
        10'b1001101000: data <= 19'h7fe6b; 
        10'b1001101001: data <= 19'h7ff94; 
        10'b1001101010: data <= 19'h7fea3; 
        10'b1001101011: data <= 19'h00073; 
        10'b1001101100: data <= 19'h00199; 
        10'b1001101101: data <= 19'h00094; 
        10'b1001101110: data <= 19'h00376; 
        10'b1001101111: data <= 19'h00309; 
        10'b1001110000: data <= 19'h002d4; 
        10'b1001110001: data <= 19'h003f9; 
        10'b1001110010: data <= 19'h003f2; 
        10'b1001110011: data <= 19'h004ae; 
        10'b1001110100: data <= 19'h00082; 
        10'b1001110101: data <= 19'h7fc4e; 
        10'b1001110110: data <= 19'h7fb59; 
        10'b1001110111: data <= 19'h7fd5e; 
        10'b1001111000: data <= 19'h7fd85; 
        10'b1001111001: data <= 19'h001ee; 
        10'b1001111010: data <= 19'h0060f; 
        10'b1001111011: data <= 19'h007bc; 
        10'b1001111100: data <= 19'h00708; 
        10'b1001111101: data <= 19'h006ba; 
        10'b1001111110: data <= 19'h005d7; 
        10'b1001111111: data <= 19'h00671; 
        10'b1010000000: data <= 19'h00265; 
        10'b1010000001: data <= 19'h7ffbc; 
        10'b1010000010: data <= 19'h7ff97; 
        10'b1010000011: data <= 19'h7fee1; 
        10'b1010000100: data <= 19'h7ff9e; 
        10'b1010000101: data <= 19'h7ffaa; 
        10'b1010000110: data <= 19'h7ff4d; 
        10'b1010000111: data <= 19'h7ff30; 
        10'b1010001000: data <= 19'h7ff18; 
        10'b1010001001: data <= 19'h7fe33; 
        10'b1010001010: data <= 19'h7fdca; 
        10'b1010001011: data <= 19'h7fe15; 
        10'b1010001100: data <= 19'h7fcda; 
        10'b1010001101: data <= 19'h7fe28; 
        10'b1010001110: data <= 19'h7fec4; 
        10'b1010001111: data <= 19'h00197; 
        10'b1010010000: data <= 19'h00025; 
        10'b1010010001: data <= 19'h7fd86; 
        10'b1010010010: data <= 19'h7fca6; 
        10'b1010010011: data <= 19'h7fba0; 
        10'b1010010100: data <= 19'h7fb40; 
        10'b1010010101: data <= 19'h7fd86; 
        10'b1010010110: data <= 19'h000f8; 
        10'b1010010111: data <= 19'h0060e; 
        10'b1010011000: data <= 19'h0054c; 
        10'b1010011001: data <= 19'h0067d; 
        10'b1010011010: data <= 19'h004a8; 
        10'b1010011011: data <= 19'h001c7; 
        10'b1010011100: data <= 19'h00113; 
        10'b1010011101: data <= 19'h000b0; 
        10'b1010011110: data <= 19'h7ffd9; 
        10'b1010011111: data <= 19'h7ff2b; 
        10'b1010100000: data <= 19'h7ff68; 
        10'b1010100001: data <= 19'h7fec6; 
        10'b1010100010: data <= 19'h7fff1; 
        10'b1010100011: data <= 19'h7ffca; 
        10'b1010100100: data <= 19'h7feb3; 
        10'b1010100101: data <= 19'h7fc9d; 
        10'b1010100110: data <= 19'h7f974; 
        10'b1010100111: data <= 19'h7fb1b; 
        10'b1010101000: data <= 19'h7faf6; 
        10'b1010101001: data <= 19'h7faa0; 
        10'b1010101010: data <= 19'h7faaa; 
        10'b1010101011: data <= 19'h7fbea; 
        10'b1010101100: data <= 19'h7fbe2; 
        10'b1010101101: data <= 19'h7fdc3; 
        10'b1010101110: data <= 19'h7fd15; 
        10'b1010101111: data <= 19'h7fbd7; 
        10'b1010110000: data <= 19'h7fc0d; 
        10'b1010110001: data <= 19'h7fce7; 
        10'b1010110010: data <= 19'h7fc37; 
        10'b1010110011: data <= 19'h7fdf5; 
        10'b1010110100: data <= 19'h7fe31; 
        10'b1010110101: data <= 19'h7fe34; 
        10'b1010110110: data <= 19'h7fef3; 
        10'b1010110111: data <= 19'h7ff2b; 
        10'b1010111000: data <= 19'h7ffe0; 
        10'b1010111001: data <= 19'h000ad; 
        10'b1010111010: data <= 19'h7fe96; 
        10'b1010111011: data <= 19'h7fea0; 
        10'b1010111100: data <= 19'h7fff1; 
        10'b1010111101: data <= 19'h7fe3b; 
        10'b1010111110: data <= 19'h7ff1a; 
        10'b1010111111: data <= 19'h7feeb; 
        10'b1011000000: data <= 19'h7fe9a; 
        10'b1011000001: data <= 19'h7fd9d; 
        10'b1011000010: data <= 19'h7fcd2; 
        10'b1011000011: data <= 19'h7fb2a; 
        10'b1011000100: data <= 19'h7faa1; 
        10'b1011000101: data <= 19'h7fb05; 
        10'b1011000110: data <= 19'h7fb7e; 
        10'b1011000111: data <= 19'h7fa42; 
        10'b1011001000: data <= 19'h7fc27; 
        10'b1011001001: data <= 19'h7fc65; 
        10'b1011001010: data <= 19'h7fb37; 
        10'b1011001011: data <= 19'h7fc0e; 
        10'b1011001100: data <= 19'h7fd13; 
        10'b1011001101: data <= 19'h7fd41; 
        10'b1011001110: data <= 19'h7fef3; 
        10'b1011001111: data <= 19'h7fd7e; 
        10'b1011010000: data <= 19'h7ff19; 
        10'b1011010001: data <= 19'h7ff08; 
        10'b1011010010: data <= 19'h7fff5; 
        10'b1011010011: data <= 19'h7fea6; 
        10'b1011010100: data <= 19'h7ff7e; 
        10'b1011010101: data <= 19'h7fead; 
        10'b1011010110: data <= 19'h7fe48; 
        10'b1011010111: data <= 19'h7feb3; 
        10'b1011011000: data <= 19'h7fe58; 
        10'b1011011001: data <= 19'h7fef4; 
        10'b1011011010: data <= 19'h7ff3d; 
        10'b1011011011: data <= 19'h00014; 
        10'b1011011100: data <= 19'h7ffbb; 
        10'b1011011101: data <= 19'h7ff2c; 
        10'b1011011110: data <= 19'h7ffab; 
        10'b1011011111: data <= 19'h7fff1; 
        10'b1011100000: data <= 19'h7ff23; 
        10'b1011100001: data <= 19'h0001a; 
        10'b1011100010: data <= 19'h7fff8; 
        10'b1011100011: data <= 19'h0000f; 
        10'b1011100100: data <= 19'h00029; 
        10'b1011100101: data <= 19'h7ff7e; 
        10'b1011100110: data <= 19'h7feda; 
        10'b1011100111: data <= 19'h7fe1f; 
        10'b1011101000: data <= 19'h7ff03; 
        10'b1011101001: data <= 19'h7ff7a; 
        10'b1011101010: data <= 19'h7ff60; 
        10'b1011101011: data <= 19'h7fea9; 
        10'b1011101100: data <= 19'h0002c; 
        10'b1011101101: data <= 19'h7fff8; 
        10'b1011101110: data <= 19'h7fead; 
        10'b1011101111: data <= 19'h7fef4; 
        10'b1011110000: data <= 19'h7fe52; 
        10'b1011110001: data <= 19'h00013; 
        10'b1011110010: data <= 19'h0000e; 
        10'b1011110011: data <= 19'h7ffe9; 
        10'b1011110100: data <= 19'h7ffdc; 
        10'b1011110101: data <= 19'h7fec7; 
        10'b1011110110: data <= 19'h7fe7a; 
        10'b1011110111: data <= 19'h7ff65; 
        10'b1011111000: data <= 19'h7fe4c; 
        10'b1011111001: data <= 19'h0005a; 
        10'b1011111010: data <= 19'h00052; 
        10'b1011111011: data <= 19'h7ff02; 
        10'b1011111100: data <= 19'h7ffe5; 
        10'b1011111101: data <= 19'h7fea9; 
        10'b1011111110: data <= 19'h0003c; 
        10'b1011111111: data <= 19'h7fe41; 
        10'b1100000000: data <= 19'h7ffe8; 
        10'b1100000001: data <= 19'h7ff28; 
        10'b1100000010: data <= 19'h7ff9b; 
        10'b1100000011: data <= 19'h7fe84; 
        10'b1100000100: data <= 19'h7ff63; 
        10'b1100000101: data <= 19'h7ff17; 
        10'b1100000110: data <= 19'h7ff7a; 
        10'b1100000111: data <= 19'h7ff59; 
        10'b1100001000: data <= 19'h7ffce; 
        10'b1100001001: data <= 19'h7fe30; 
        10'b1100001010: data <= 19'h7ff38; 
        10'b1100001011: data <= 19'h0000f; 
        10'b1100001100: data <= 19'h7fe2f; 
        10'b1100001101: data <= 19'h7ff50; 
        10'b1100001110: data <= 19'h7ffbe; 
        10'b1100001111: data <= 19'h7ff07; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 14) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 20'hffcc9; 
        10'b0000000001: data <= 20'h00013; 
        10'b0000000010: data <= 20'hffe66; 
        10'b0000000011: data <= 20'hffd59; 
        10'b0000000100: data <= 20'hffe5b; 
        10'b0000000101: data <= 20'hffd87; 
        10'b0000000110: data <= 20'hffeeb; 
        10'b0000000111: data <= 20'hfff16; 
        10'b0000001000: data <= 20'hffcb2; 
        10'b0000001001: data <= 20'hffea8; 
        10'b0000001010: data <= 20'hffcef; 
        10'b0000001011: data <= 20'hffdf6; 
        10'b0000001100: data <= 20'h0009e; 
        10'b0000001101: data <= 20'h0008a; 
        10'b0000001110: data <= 20'hffcde; 
        10'b0000001111: data <= 20'hffedf; 
        10'b0000010000: data <= 20'hffd17; 
        10'b0000010001: data <= 20'hffd21; 
        10'b0000010010: data <= 20'h000d5; 
        10'b0000010011: data <= 20'h0003d; 
        10'b0000010100: data <= 20'hffd9d; 
        10'b0000010101: data <= 20'hffefa; 
        10'b0000010110: data <= 20'hffde2; 
        10'b0000010111: data <= 20'hffc80; 
        10'b0000011000: data <= 20'hffcc9; 
        10'b0000011001: data <= 20'hffec9; 
        10'b0000011010: data <= 20'hfffd8; 
        10'b0000011011: data <= 20'hfff1e; 
        10'b0000011100: data <= 20'hffea3; 
        10'b0000011101: data <= 20'hffe6b; 
        10'b0000011110: data <= 20'h000c7; 
        10'b0000011111: data <= 20'hfff33; 
        10'b0000100000: data <= 20'hffcf3; 
        10'b0000100001: data <= 20'hffcd9; 
        10'b0000100010: data <= 20'hffcba; 
        10'b0000100011: data <= 20'hffd85; 
        10'b0000100100: data <= 20'hffd8e; 
        10'b0000100101: data <= 20'hffedb; 
        10'b0000100110: data <= 20'h00008; 
        10'b0000100111: data <= 20'hffd10; 
        10'b0000101000: data <= 20'hffe1f; 
        10'b0000101001: data <= 20'hffcf5; 
        10'b0000101010: data <= 20'hffeeb; 
        10'b0000101011: data <= 20'hffc80; 
        10'b0000101100: data <= 20'hfff12; 
        10'b0000101101: data <= 20'hffd12; 
        10'b0000101110: data <= 20'hffe07; 
        10'b0000101111: data <= 20'hffd49; 
        10'b0000110000: data <= 20'hffee4; 
        10'b0000110001: data <= 20'hffd25; 
        10'b0000110010: data <= 20'hffca8; 
        10'b0000110011: data <= 20'hffc57; 
        10'b0000110100: data <= 20'h0002e; 
        10'b0000110101: data <= 20'hfff31; 
        10'b0000110110: data <= 20'h0003c; 
        10'b0000110111: data <= 20'hffdcc; 
        10'b0000111000: data <= 20'hffe70; 
        10'b0000111001: data <= 20'hffc8e; 
        10'b0000111010: data <= 20'hffce0; 
        10'b0000111011: data <= 20'hffff9; 
        10'b0000111100: data <= 20'hffcad; 
        10'b0000111101: data <= 20'hffcf5; 
        10'b0000111110: data <= 20'hffe46; 
        10'b0000111111: data <= 20'hffec9; 
        10'b0001000000: data <= 20'hfffad; 
        10'b0001000001: data <= 20'hffe1c; 
        10'b0001000010: data <= 20'h001cf; 
        10'b0001000011: data <= 20'h0017e; 
        10'b0001000100: data <= 20'h0049f; 
        10'b0001000101: data <= 20'h003af; 
        10'b0001000110: data <= 20'h0035f; 
        10'b0001000111: data <= 20'h00157; 
        10'b0001001000: data <= 20'h00489; 
        10'b0001001001: data <= 20'h0018c; 
        10'b0001001010: data <= 20'h00150; 
        10'b0001001011: data <= 20'hffdb3; 
        10'b0001001100: data <= 20'hffff0; 
        10'b0001001101: data <= 20'hffeef; 
        10'b0001001110: data <= 20'hffb4e; 
        10'b0001001111: data <= 20'hffe59; 
        10'b0001010000: data <= 20'hfff80; 
        10'b0001010001: data <= 20'h00122; 
        10'b0001010010: data <= 20'hffea7; 
        10'b0001010011: data <= 20'hffe19; 
        10'b0001010100: data <= 20'hffdb6; 
        10'b0001010101: data <= 20'hffd66; 
        10'b0001010110: data <= 20'hfff42; 
        10'b0001010111: data <= 20'hffd9d; 
        10'b0001011000: data <= 20'h000a6; 
        10'b0001011001: data <= 20'hffd1a; 
        10'b0001011010: data <= 20'hffef1; 
        10'b0001011011: data <= 20'h00001; 
        10'b0001011100: data <= 20'h000d3; 
        10'b0001011101: data <= 20'h0075c; 
        10'b0001011110: data <= 20'h00b85; 
        10'b0001011111: data <= 20'h00b71; 
        10'b0001100000: data <= 20'h00af3; 
        10'b0001100001: data <= 20'h0101b; 
        10'b0001100010: data <= 20'h008ca; 
        10'b0001100011: data <= 20'h003e6; 
        10'b0001100100: data <= 20'h00768; 
        10'b0001100101: data <= 20'h00365; 
        10'b0001100110: data <= 20'hffccc; 
        10'b0001100111: data <= 20'hfff35; 
        10'b0001101000: data <= 20'hffc5c; 
        10'b0001101001: data <= 20'hffbbc; 
        10'b0001101010: data <= 20'hffac9; 
        10'b0001101011: data <= 20'hffd6a; 
        10'b0001101100: data <= 20'h00062; 
        10'b0001101101: data <= 20'h0013a; 
        10'b0001101110: data <= 20'hffd1e; 
        10'b0001101111: data <= 20'hfff6b; 
        10'b0001110000: data <= 20'hffd7a; 
        10'b0001110001: data <= 20'hffe3f; 
        10'b0001110010: data <= 20'h000e2; 
        10'b0001110011: data <= 20'hffc3c; 
        10'b0001110100: data <= 20'hffcae; 
        10'b0001110101: data <= 20'hffef1; 
        10'b0001110110: data <= 20'h001b5; 
        10'b0001110111: data <= 20'h001a5; 
        10'b0001111000: data <= 20'h004be; 
        10'b0001111001: data <= 20'h00e1a; 
        10'b0001111010: data <= 20'h00e3f; 
        10'b0001111011: data <= 20'h011e7; 
        10'b0001111100: data <= 20'h00f21; 
        10'b0001111101: data <= 20'h00c00; 
        10'b0001111110: data <= 20'h00ae7; 
        10'b0001111111: data <= 20'h004d1; 
        10'b0010000000: data <= 20'h00672; 
        10'b0010000001: data <= 20'h005f5; 
        10'b0010000010: data <= 20'hffe37; 
        10'b0010000011: data <= 20'hffcfe; 
        10'b0010000100: data <= 20'hffdae; 
        10'b0010000101: data <= 20'hff8ec; 
        10'b0010000110: data <= 20'hff76e; 
        10'b0010000111: data <= 20'hff7c4; 
        10'b0010001000: data <= 20'hffef2; 
        10'b0010001001: data <= 20'hffef1; 
        10'b0010001010: data <= 20'hffc8e; 
        10'b0010001011: data <= 20'hfff5a; 
        10'b0010001100: data <= 20'h0004c; 
        10'b0010001101: data <= 20'hffee2; 
        10'b0010001110: data <= 20'hffd49; 
        10'b0010001111: data <= 20'hffc5f; 
        10'b0010010000: data <= 20'hffd05; 
        10'b0010010001: data <= 20'hffd70; 
        10'b0010010010: data <= 20'h00194; 
        10'b0010010011: data <= 20'h006e4; 
        10'b0010010100: data <= 20'h0098e; 
        10'b0010010101: data <= 20'h0105c; 
        10'b0010010110: data <= 20'h0121f; 
        10'b0010010111: data <= 20'h012e7; 
        10'b0010011000: data <= 20'h01150; 
        10'b0010011001: data <= 20'h0136a; 
        10'b0010011010: data <= 20'h011f8; 
        10'b0010011011: data <= 20'h010ac; 
        10'b0010011100: data <= 20'h01215; 
        10'b0010011101: data <= 20'h00ea0; 
        10'b0010011110: data <= 20'h00a91; 
        10'b0010011111: data <= 20'hffb89; 
        10'b0010100000: data <= 20'hffbb1; 
        10'b0010100001: data <= 20'hff8f6; 
        10'b0010100010: data <= 20'hff8d8; 
        10'b0010100011: data <= 20'hff4e7; 
        10'b0010100100: data <= 20'hffb36; 
        10'b0010100101: data <= 20'hffd47; 
        10'b0010100110: data <= 20'h00071; 
        10'b0010100111: data <= 20'hffde2; 
        10'b0010101000: data <= 20'hffe8e; 
        10'b0010101001: data <= 20'hffd6a; 
        10'b0010101010: data <= 20'h00095; 
        10'b0010101011: data <= 20'hffe9c; 
        10'b0010101100: data <= 20'hffe2e; 
        10'b0010101101: data <= 20'h00127; 
        10'b0010101110: data <= 20'h006bd; 
        10'b0010101111: data <= 20'h00d0c; 
        10'b0010110000: data <= 20'h009f9; 
        10'b0010110001: data <= 20'h00b52; 
        10'b0010110010: data <= 20'h00f53; 
        10'b0010110011: data <= 20'h00996; 
        10'b0010110100: data <= 20'h00a2f; 
        10'b0010110101: data <= 20'h00d27; 
        10'b0010110110: data <= 20'h00b9e; 
        10'b0010110111: data <= 20'h00652; 
        10'b0010111000: data <= 20'h006ff; 
        10'b0010111001: data <= 20'h001cf; 
        10'b0010111010: data <= 20'h00156; 
        10'b0010111011: data <= 20'hffbe5; 
        10'b0010111100: data <= 20'hffd45; 
        10'b0010111101: data <= 20'hff70b; 
        10'b0010111110: data <= 20'hff71c; 
        10'b0010111111: data <= 20'hff399; 
        10'b0011000000: data <= 20'hff89d; 
        10'b0011000001: data <= 20'hffbdc; 
        10'b0011000010: data <= 20'h00086; 
        10'b0011000011: data <= 20'hfff94; 
        10'b0011000100: data <= 20'hffe16; 
        10'b0011000101: data <= 20'h00062; 
        10'b0011000110: data <= 20'h0006b; 
        10'b0011000111: data <= 20'hffe41; 
        10'b0011001000: data <= 20'h0002d; 
        10'b0011001001: data <= 20'h0039f; 
        10'b0011001010: data <= 20'h008af; 
        10'b0011001011: data <= 20'h00c92; 
        10'b0011001100: data <= 20'h00a49; 
        10'b0011001101: data <= 20'h00999; 
        10'b0011001110: data <= 20'h003ab; 
        10'b0011001111: data <= 20'h00455; 
        10'b0011010000: data <= 20'h000bd; 
        10'b0011010001: data <= 20'h006bd; 
        10'b0011010010: data <= 20'h0084d; 
        10'b0011010011: data <= 20'h001bd; 
        10'b0011010100: data <= 20'h0011d; 
        10'b0011010101: data <= 20'hff57c; 
        10'b0011010110: data <= 20'hffc6f; 
        10'b0011010111: data <= 20'hffd08; 
        10'b0011011000: data <= 20'hffca2; 
        10'b0011011001: data <= 20'hffc0f; 
        10'b0011011010: data <= 20'hffd10; 
        10'b0011011011: data <= 20'hff5cc; 
        10'b0011011100: data <= 20'hff8ef; 
        10'b0011011101: data <= 20'hffdd8; 
        10'b0011011110: data <= 20'hffd48; 
        10'b0011011111: data <= 20'hffcaf; 
        10'b0011100000: data <= 20'hfff3e; 
        10'b0011100001: data <= 20'h0007f; 
        10'b0011100010: data <= 20'hffe96; 
        10'b0011100011: data <= 20'h00075; 
        10'b0011100100: data <= 20'h001e5; 
        10'b0011100101: data <= 20'h005e1; 
        10'b0011100110: data <= 20'h00440; 
        10'b0011100111: data <= 20'h00601; 
        10'b0011101000: data <= 20'h00614; 
        10'b0011101001: data <= 20'h006c3; 
        10'b0011101010: data <= 20'h006cb; 
        10'b0011101011: data <= 20'h007c1; 
        10'b0011101100: data <= 20'h0049c; 
        10'b0011101101: data <= 20'h00582; 
        10'b0011101110: data <= 20'h00e87; 
        10'b0011101111: data <= 20'h0082b; 
        10'b0011110000: data <= 20'hffefe; 
        10'b0011110001: data <= 20'hffc03; 
        10'b0011110010: data <= 20'hfffe6; 
        10'b0011110011: data <= 20'h00339; 
        10'b0011110100: data <= 20'h00013; 
        10'b0011110101: data <= 20'hffdc6; 
        10'b0011110110: data <= 20'hffa14; 
        10'b0011110111: data <= 20'hff418; 
        10'b0011111000: data <= 20'hff6dd; 
        10'b0011111001: data <= 20'hffc31; 
        10'b0011111010: data <= 20'hffe38; 
        10'b0011111011: data <= 20'hffd13; 
        10'b0011111100: data <= 20'hffd7d; 
        10'b0011111101: data <= 20'hfff63; 
        10'b0011111110: data <= 20'hfffdd; 
        10'b0011111111: data <= 20'h00186; 
        10'b0100000000: data <= 20'h002f5; 
        10'b0100000001: data <= 20'h00696; 
        10'b0100000010: data <= 20'h0024e; 
        10'b0100000011: data <= 20'h00072; 
        10'b0100000100: data <= 20'hffdba; 
        10'b0100000101: data <= 20'h0038b; 
        10'b0100000110: data <= 20'h002c0; 
        10'b0100000111: data <= 20'h0038e; 
        10'b0100001000: data <= 20'h000ec; 
        10'b0100001001: data <= 20'hfffa2; 
        10'b0100001010: data <= 20'h0097b; 
        10'b0100001011: data <= 20'h00a40; 
        10'b0100001100: data <= 20'h00389; 
        10'b0100001101: data <= 20'h00045; 
        10'b0100001110: data <= 20'hfff0c; 
        10'b0100001111: data <= 20'hfffea; 
        10'b0100010000: data <= 20'hfff92; 
        10'b0100010001: data <= 20'hfffc5; 
        10'b0100010010: data <= 20'hffc3d; 
        10'b0100010011: data <= 20'hff5e0; 
        10'b0100010100: data <= 20'hff75c; 
        10'b0100010101: data <= 20'hffd30; 
        10'b0100010110: data <= 20'h00072; 
        10'b0100010111: data <= 20'hffcbc; 
        10'b0100011000: data <= 20'h000a3; 
        10'b0100011001: data <= 20'hfff42; 
        10'b0100011010: data <= 20'hffe80; 
        10'b0100011011: data <= 20'hffde0; 
        10'b0100011100: data <= 20'h00073; 
        10'b0100011101: data <= 20'hffe64; 
        10'b0100011110: data <= 20'hffcb5; 
        10'b0100011111: data <= 20'hff005; 
        10'b0100100000: data <= 20'hff1b3; 
        10'b0100100001: data <= 20'hff532; 
        10'b0100100010: data <= 20'hfef7d; 
        10'b0100100011: data <= 20'hfedb0; 
        10'b0100100100: data <= 20'hfeab1; 
        10'b0100100101: data <= 20'hfe813; 
        10'b0100100110: data <= 20'hff5f4; 
        10'b0100100111: data <= 20'h001d3; 
        10'b0100101000: data <= 20'h00296; 
        10'b0100101001: data <= 20'h0006f; 
        10'b0100101010: data <= 20'h00154; 
        10'b0100101011: data <= 20'hffe0e; 
        10'b0100101100: data <= 20'hffe96; 
        10'b0100101101: data <= 20'hffe0d; 
        10'b0100101110: data <= 20'hffafc; 
        10'b0100101111: data <= 20'hff45a; 
        10'b0100110000: data <= 20'hff99a; 
        10'b0100110001: data <= 20'hfffba; 
        10'b0100110010: data <= 20'hfffb5; 
        10'b0100110011: data <= 20'hffd4f; 
        10'b0100110100: data <= 20'hffcac; 
        10'b0100110101: data <= 20'h000d2; 
        10'b0100110110: data <= 20'hfffa9; 
        10'b0100110111: data <= 20'hffcf1; 
        10'b0100111000: data <= 20'hffa02; 
        10'b0100111001: data <= 20'hff2e8; 
        10'b0100111010: data <= 20'hfe987; 
        10'b0100111011: data <= 20'hfe050; 
        10'b0100111100: data <= 20'hfe190; 
        10'b0100111101: data <= 20'hfdc27; 
        10'b0100111110: data <= 20'hfdc0c; 
        10'b0100111111: data <= 20'hfdf2f; 
        10'b0101000000: data <= 20'hfdd2b; 
        10'b0101000001: data <= 20'hfd58e; 
        10'b0101000010: data <= 20'hfdf59; 
        10'b0101000011: data <= 20'hff062; 
        10'b0101000100: data <= 20'hffa96; 
        10'b0101000101: data <= 20'hffb58; 
        10'b0101000110: data <= 20'hffb86; 
        10'b0101000111: data <= 20'hfff1b; 
        10'b0101001000: data <= 20'hffd50; 
        10'b0101001001: data <= 20'hffd32; 
        10'b0101001010: data <= 20'hff895; 
        10'b0101001011: data <= 20'hffaec; 
        10'b0101001100: data <= 20'hfff14; 
        10'b0101001101: data <= 20'hffe3f; 
        10'b0101001110: data <= 20'hffd39; 
        10'b0101001111: data <= 20'hfff3b; 
        10'b0101010000: data <= 20'hffed9; 
        10'b0101010001: data <= 20'hfff0c; 
        10'b0101010010: data <= 20'h00055; 
        10'b0101010011: data <= 20'hffe9a; 
        10'b0101010100: data <= 20'hff98d; 
        10'b0101010101: data <= 20'hfec80; 
        10'b0101010110: data <= 20'hfda11; 
        10'b0101010111: data <= 20'hfd196; 
        10'b0101011000: data <= 20'hfd4b6; 
        10'b0101011001: data <= 20'hfd6f9; 
        10'b0101011010: data <= 20'hfda82; 
        10'b0101011011: data <= 20'hfdceb; 
        10'b0101011100: data <= 20'hfdd05; 
        10'b0101011101: data <= 20'hfdb9a; 
        10'b0101011110: data <= 20'hfe21a; 
        10'b0101011111: data <= 20'hfec10; 
        10'b0101100000: data <= 20'hff251; 
        10'b0101100001: data <= 20'hff3b6; 
        10'b0101100010: data <= 20'hff9cf; 
        10'b0101100011: data <= 20'h00007; 
        10'b0101100100: data <= 20'hfffe1; 
        10'b0101100101: data <= 20'hffc87; 
        10'b0101100110: data <= 20'hff81b; 
        10'b0101100111: data <= 20'hff3fe; 
        10'b0101101000: data <= 20'hffe8a; 
        10'b0101101001: data <= 20'hffe03; 
        10'b0101101010: data <= 20'h000e4; 
        10'b0101101011: data <= 20'hfff0c; 
        10'b0101101100: data <= 20'hffd96; 
        10'b0101101101: data <= 20'hffe6b; 
        10'b0101101110: data <= 20'h000d5; 
        10'b0101101111: data <= 20'hffd81; 
        10'b0101110000: data <= 20'hff58f; 
        10'b0101110001: data <= 20'hfe769; 
        10'b0101110010: data <= 20'hfd8fb; 
        10'b0101110011: data <= 20'hfdc2f; 
        10'b0101110100: data <= 20'hfde92; 
        10'b0101110101: data <= 20'hfe906; 
        10'b0101110110: data <= 20'hfefb7; 
        10'b0101110111: data <= 20'hff860; 
        10'b0101111000: data <= 20'hff3f0; 
        10'b0101111001: data <= 20'hffa84; 
        10'b0101111010: data <= 20'hff23a; 
        10'b0101111011: data <= 20'hff1f2; 
        10'b0101111100: data <= 20'hfef54; 
        10'b0101111101: data <= 20'hff3f7; 
        10'b0101111110: data <= 20'hff95f; 
        10'b0101111111: data <= 20'hffebb; 
        10'b0110000000: data <= 20'hffe0e; 
        10'b0110000001: data <= 20'hffbba; 
        10'b0110000010: data <= 20'hff613; 
        10'b0110000011: data <= 20'hff6f7; 
        10'b0110000100: data <= 20'hffb6e; 
        10'b0110000101: data <= 20'h00125; 
        10'b0110000110: data <= 20'hffe79; 
        10'b0110000111: data <= 20'hfffe6; 
        10'b0110001000: data <= 20'h00085; 
        10'b0110001001: data <= 20'hfff2c; 
        10'b0110001010: data <= 20'h00016; 
        10'b0110001011: data <= 20'hffde6; 
        10'b0110001100: data <= 20'hffc00; 
        10'b0110001101: data <= 20'hfef64; 
        10'b0110001110: data <= 20'hfeafd; 
        10'b0110001111: data <= 20'hfeedf; 
        10'b0110010000: data <= 20'hff921; 
        10'b0110010001: data <= 20'hffed1; 
        10'b0110010010: data <= 20'h00449; 
        10'b0110010011: data <= 20'h005ab; 
        10'b0110010100: data <= 20'h006ba; 
        10'b0110010101: data <= 20'h00a77; 
        10'b0110010110: data <= 20'h000b7; 
        10'b0110010111: data <= 20'hff94d; 
        10'b0110011000: data <= 20'hffb05; 
        10'b0110011001: data <= 20'hff760; 
        10'b0110011010: data <= 20'hffe8c; 
        10'b0110011011: data <= 20'hffa74; 
        10'b0110011100: data <= 20'hffe3f; 
        10'b0110011101: data <= 20'hff99c; 
        10'b0110011110: data <= 20'hff483; 
        10'b0110011111: data <= 20'hff7a5; 
        10'b0110100000: data <= 20'hffe5e; 
        10'b0110100001: data <= 20'h00411; 
        10'b0110100010: data <= 20'h0049d; 
        10'b0110100011: data <= 20'hffd6f; 
        10'b0110100100: data <= 20'hffe34; 
        10'b0110100101: data <= 20'hffe95; 
        10'b0110100110: data <= 20'hffe26; 
        10'b0110100111: data <= 20'h003cc; 
        10'b0110101000: data <= 20'h001d6; 
        10'b0110101001: data <= 20'h000d4; 
        10'b0110101010: data <= 20'h0047e; 
        10'b0110101011: data <= 20'h00543; 
        10'b0110101100: data <= 20'h009c7; 
        10'b0110101101: data <= 20'h006e9; 
        10'b0110101110: data <= 20'h00849; 
        10'b0110101111: data <= 20'h004df; 
        10'b0110110000: data <= 20'h00450; 
        10'b0110110001: data <= 20'h00a1c; 
        10'b0110110010: data <= 20'h000c0; 
        10'b0110110011: data <= 20'h003f8; 
        10'b0110110100: data <= 20'h00091; 
        10'b0110110101: data <= 20'hff7fb; 
        10'b0110110110: data <= 20'hff85f; 
        10'b0110110111: data <= 20'hffb52; 
        10'b0110111000: data <= 20'hffc97; 
        10'b0110111001: data <= 20'hffad7; 
        10'b0110111010: data <= 20'hff597; 
        10'b0110111011: data <= 20'hffaa5; 
        10'b0110111100: data <= 20'h00333; 
        10'b0110111101: data <= 20'h00574; 
        10'b0110111110: data <= 20'h002f2; 
        10'b0110111111: data <= 20'hffd15; 
        10'b0111000000: data <= 20'hffdc6; 
        10'b0111000001: data <= 20'hffc8a; 
        10'b0111000010: data <= 20'hffc14; 
        10'b0111000011: data <= 20'h0040a; 
        10'b0111000100: data <= 20'h00878; 
        10'b0111000101: data <= 20'h00dd4; 
        10'b0111000110: data <= 20'h00e16; 
        10'b0111000111: data <= 20'h00862; 
        10'b0111001000: data <= 20'h0037a; 
        10'b0111001001: data <= 20'h0073b; 
        10'b0111001010: data <= 20'h006b7; 
        10'b0111001011: data <= 20'h00622; 
        10'b0111001100: data <= 20'h00ca3; 
        10'b0111001101: data <= 20'h00b20; 
        10'b0111001110: data <= 20'h00256; 
        10'b0111001111: data <= 20'hffeac; 
        10'b0111010000: data <= 20'hffff3; 
        10'b0111010001: data <= 20'hffacb; 
        10'b0111010010: data <= 20'hffb72; 
        10'b0111010011: data <= 20'hff803; 
        10'b0111010100: data <= 20'hffd29; 
        10'b0111010101: data <= 20'h0006f; 
        10'b0111010110: data <= 20'h001c2; 
        10'b0111010111: data <= 20'h003b6; 
        10'b0111011000: data <= 20'h00bcc; 
        10'b0111011001: data <= 20'h00e9d; 
        10'b0111011010: data <= 20'h00272; 
        10'b0111011011: data <= 20'hffdb7; 
        10'b0111011100: data <= 20'hffe1c; 
        10'b0111011101: data <= 20'h000ab; 
        10'b0111011110: data <= 20'hffe87; 
        10'b0111011111: data <= 20'h004e5; 
        10'b0111100000: data <= 20'h00e77; 
        10'b0111100001: data <= 20'h01427; 
        10'b0111100010: data <= 20'h0126b; 
        10'b0111100011: data <= 20'h00c9e; 
        10'b0111100100: data <= 20'h008c8; 
        10'b0111100101: data <= 20'h00aa6; 
        10'b0111100110: data <= 20'h01060; 
        10'b0111100111: data <= 20'h00d6b; 
        10'b0111101000: data <= 20'h00f64; 
        10'b0111101001: data <= 20'h00733; 
        10'b0111101010: data <= 20'h003b6; 
        10'b0111101011: data <= 20'h00501; 
        10'b0111101100: data <= 20'h0050e; 
        10'b0111101101: data <= 20'hfff38; 
        10'b0111101110: data <= 20'h00347; 
        10'b0111101111: data <= 20'hffde9; 
        10'b0111110000: data <= 20'h0060c; 
        10'b0111110001: data <= 20'h00673; 
        10'b0111110010: data <= 20'h004cb; 
        10'b0111110011: data <= 20'h006a4; 
        10'b0111110100: data <= 20'h012e7; 
        10'b0111110101: data <= 20'h01066; 
        10'b0111110110: data <= 20'h003be; 
        10'b0111110111: data <= 20'h0007f; 
        10'b0111111000: data <= 20'hfff93; 
        10'b0111111001: data <= 20'hfffc5; 
        10'b0111111010: data <= 20'hffb05; 
        10'b0111111011: data <= 20'h00151; 
        10'b0111111100: data <= 20'h00fad; 
        10'b0111111101: data <= 20'h01a7d; 
        10'b0111111110: data <= 20'h018ea; 
        10'b0111111111: data <= 20'h011ef; 
        10'b1000000000: data <= 20'h00bf7; 
        10'b1000000001: data <= 20'h00d4d; 
        10'b1000000010: data <= 20'h01453; 
        10'b1000000011: data <= 20'h0125d; 
        10'b1000000100: data <= 20'h01d41; 
        10'b1000000101: data <= 20'h0155a; 
        10'b1000000110: data <= 20'h012a5; 
        10'b1000000111: data <= 20'h00913; 
        10'b1000001000: data <= 20'h0063f; 
        10'b1000001001: data <= 20'h00b78; 
        10'b1000001010: data <= 20'h00767; 
        10'b1000001011: data <= 20'h0050a; 
        10'b1000001100: data <= 20'h00d88; 
        10'b1000001101: data <= 20'h00dfb; 
        10'b1000001110: data <= 20'h00f3c; 
        10'b1000001111: data <= 20'h01422; 
        10'b1000010000: data <= 20'h018fc; 
        10'b1000010001: data <= 20'h00e68; 
        10'b1000010010: data <= 20'hffe9e; 
        10'b1000010011: data <= 20'hffd08; 
        10'b1000010100: data <= 20'hffd78; 
        10'b1000010101: data <= 20'hffda3; 
        10'b1000010110: data <= 20'hffc86; 
        10'b1000010111: data <= 20'hffff1; 
        10'b1000011000: data <= 20'h0089d; 
        10'b1000011001: data <= 20'h01017; 
        10'b1000011010: data <= 20'h01452; 
        10'b1000011011: data <= 20'h0119f; 
        10'b1000011100: data <= 20'h01044; 
        10'b1000011101: data <= 20'h01138; 
        10'b1000011110: data <= 20'h0107a; 
        10'b1000011111: data <= 20'h01180; 
        10'b1000100000: data <= 20'h01396; 
        10'b1000100001: data <= 20'h00f11; 
        10'b1000100010: data <= 20'h009c2; 
        10'b1000100011: data <= 20'h004a0; 
        10'b1000100100: data <= 20'h00730; 
        10'b1000100101: data <= 20'h00c7b; 
        10'b1000100110: data <= 20'h00607; 
        10'b1000100111: data <= 20'h005e4; 
        10'b1000101000: data <= 20'h00a0e; 
        10'b1000101001: data <= 20'h00c8c; 
        10'b1000101010: data <= 20'h01062; 
        10'b1000101011: data <= 20'h01192; 
        10'b1000101100: data <= 20'h00f25; 
        10'b1000101101: data <= 20'h007ef; 
        10'b1000101110: data <= 20'h000ac; 
        10'b1000101111: data <= 20'h0002f; 
        10'b1000110000: data <= 20'hffcdd; 
        10'b1000110001: data <= 20'hfffc1; 
        10'b1000110010: data <= 20'hfff2a; 
        10'b1000110011: data <= 20'hffbb0; 
        10'b1000110100: data <= 20'h007a5; 
        10'b1000110101: data <= 20'h00971; 
        10'b1000110110: data <= 20'h00ea8; 
        10'b1000110111: data <= 20'h01462; 
        10'b1000111000: data <= 20'h0135c; 
        10'b1000111001: data <= 20'h00cd4; 
        10'b1000111010: data <= 20'h00c55; 
        10'b1000111011: data <= 20'h014a5; 
        10'b1000111100: data <= 20'h00b7a; 
        10'b1000111101: data <= 20'h003cd; 
        10'b1000111110: data <= 20'h0028c; 
        10'b1000111111: data <= 20'h00320; 
        10'b1001000000: data <= 20'h0040c; 
        10'b1001000001: data <= 20'h0002f; 
        10'b1001000010: data <= 20'h008ed; 
        10'b1001000011: data <= 20'h00df0; 
        10'b1001000100: data <= 20'h00975; 
        10'b1001000101: data <= 20'h00d73; 
        10'b1001000110: data <= 20'h012bc; 
        10'b1001000111: data <= 20'h01040; 
        10'b1001001000: data <= 20'h00bb2; 
        10'b1001001001: data <= 20'h0058c; 
        10'b1001001010: data <= 20'hfffee; 
        10'b1001001011: data <= 20'hfff7c; 
        10'b1001001100: data <= 20'hffec5; 
        10'b1001001101: data <= 20'hffd01; 
        10'b1001001110: data <= 20'hfff76; 
        10'b1001001111: data <= 20'hffe46; 
        10'b1001010000: data <= 20'h00199; 
        10'b1001010001: data <= 20'h0040f; 
        10'b1001010010: data <= 20'h00a2b; 
        10'b1001010011: data <= 20'h00b6c; 
        10'b1001010100: data <= 20'h00a11; 
        10'b1001010101: data <= 20'h00c91; 
        10'b1001010110: data <= 20'h00b1e; 
        10'b1001010111: data <= 20'h00aea; 
        10'b1001011000: data <= 20'h00449; 
        10'b1001011001: data <= 20'h0020a; 
        10'b1001011010: data <= 20'hffee5; 
        10'b1001011011: data <= 20'h00079; 
        10'b1001011100: data <= 20'h0056e; 
        10'b1001011101: data <= 20'h005f3; 
        10'b1001011110: data <= 20'h00d08; 
        10'b1001011111: data <= 20'h00db6; 
        10'b1001100000: data <= 20'h00604; 
        10'b1001100001: data <= 20'h00d72; 
        10'b1001100010: data <= 20'h0109c; 
        10'b1001100011: data <= 20'h012eb; 
        10'b1001100100: data <= 20'h00953; 
        10'b1001100101: data <= 20'h003b2; 
        10'b1001100110: data <= 20'h000db; 
        10'b1001100111: data <= 20'hfff96; 
        10'b1001101000: data <= 20'hffcd7; 
        10'b1001101001: data <= 20'hfff27; 
        10'b1001101010: data <= 20'hffd46; 
        10'b1001101011: data <= 20'h000e6; 
        10'b1001101100: data <= 20'h00333; 
        10'b1001101101: data <= 20'h00128; 
        10'b1001101110: data <= 20'h006ec; 
        10'b1001101111: data <= 20'h00612; 
        10'b1001110000: data <= 20'h005a9; 
        10'b1001110001: data <= 20'h007f3; 
        10'b1001110010: data <= 20'h007e4; 
        10'b1001110011: data <= 20'h0095b; 
        10'b1001110100: data <= 20'h00103; 
        10'b1001110101: data <= 20'hff89c; 
        10'b1001110110: data <= 20'hff6b2; 
        10'b1001110111: data <= 20'hffabb; 
        10'b1001111000: data <= 20'hffb0a; 
        10'b1001111001: data <= 20'h003db; 
        10'b1001111010: data <= 20'h00c1e; 
        10'b1001111011: data <= 20'h00f77; 
        10'b1001111100: data <= 20'h00e10; 
        10'b1001111101: data <= 20'h00d74; 
        10'b1001111110: data <= 20'h00baf; 
        10'b1001111111: data <= 20'h00ce3; 
        10'b1010000000: data <= 20'h004ca; 
        10'b1010000001: data <= 20'hfff78; 
        10'b1010000010: data <= 20'hfff2f; 
        10'b1010000011: data <= 20'hffdc2; 
        10'b1010000100: data <= 20'hfff3c; 
        10'b1010000101: data <= 20'hfff54; 
        10'b1010000110: data <= 20'hffe9b; 
        10'b1010000111: data <= 20'hffe60; 
        10'b1010001000: data <= 20'hffe30; 
        10'b1010001001: data <= 20'hffc67; 
        10'b1010001010: data <= 20'hffb95; 
        10'b1010001011: data <= 20'hffc2a; 
        10'b1010001100: data <= 20'hff9b5; 
        10'b1010001101: data <= 20'hffc4f; 
        10'b1010001110: data <= 20'hffd88; 
        10'b1010001111: data <= 20'h0032e; 
        10'b1010010000: data <= 20'h0004b; 
        10'b1010010001: data <= 20'hffb0c; 
        10'b1010010010: data <= 20'hff94c; 
        10'b1010010011: data <= 20'hff740; 
        10'b1010010100: data <= 20'hff680; 
        10'b1010010101: data <= 20'hffb0d; 
        10'b1010010110: data <= 20'h001f1; 
        10'b1010010111: data <= 20'h00c1c; 
        10'b1010011000: data <= 20'h00a99; 
        10'b1010011001: data <= 20'h00cfa; 
        10'b1010011010: data <= 20'h00950; 
        10'b1010011011: data <= 20'h0038f; 
        10'b1010011100: data <= 20'h00227; 
        10'b1010011101: data <= 20'h0015f; 
        10'b1010011110: data <= 20'hfffb2; 
        10'b1010011111: data <= 20'hffe55; 
        10'b1010100000: data <= 20'hffed0; 
        10'b1010100001: data <= 20'hffd8b; 
        10'b1010100010: data <= 20'hfffe1; 
        10'b1010100011: data <= 20'hfff95; 
        10'b1010100100: data <= 20'hffd66; 
        10'b1010100101: data <= 20'hff939; 
        10'b1010100110: data <= 20'hff2e8; 
        10'b1010100111: data <= 20'hff636; 
        10'b1010101000: data <= 20'hff5ed; 
        10'b1010101001: data <= 20'hff53f; 
        10'b1010101010: data <= 20'hff554; 
        10'b1010101011: data <= 20'hff7d4; 
        10'b1010101100: data <= 20'hff7c3; 
        10'b1010101101: data <= 20'hffb87; 
        10'b1010101110: data <= 20'hffa29; 
        10'b1010101111: data <= 20'hff7ae; 
        10'b1010110000: data <= 20'hff81a; 
        10'b1010110001: data <= 20'hff9cf; 
        10'b1010110010: data <= 20'hff86e; 
        10'b1010110011: data <= 20'hffbe9; 
        10'b1010110100: data <= 20'hffc62; 
        10'b1010110101: data <= 20'hffc68; 
        10'b1010110110: data <= 20'hffde6; 
        10'b1010110111: data <= 20'hffe56; 
        10'b1010111000: data <= 20'hfffc0; 
        10'b1010111001: data <= 20'h0015a; 
        10'b1010111010: data <= 20'hffd2c; 
        10'b1010111011: data <= 20'hffd41; 
        10'b1010111100: data <= 20'hfffe2; 
        10'b1010111101: data <= 20'hffc76; 
        10'b1010111110: data <= 20'hffe33; 
        10'b1010111111: data <= 20'hffdd6; 
        10'b1011000000: data <= 20'hffd35; 
        10'b1011000001: data <= 20'hffb3a; 
        10'b1011000010: data <= 20'hff9a5; 
        10'b1011000011: data <= 20'hff653; 
        10'b1011000100: data <= 20'hff542; 
        10'b1011000101: data <= 20'hff60a; 
        10'b1011000110: data <= 20'hff6fb; 
        10'b1011000111: data <= 20'hff484; 
        10'b1011001000: data <= 20'hff84f; 
        10'b1011001001: data <= 20'hff8c9; 
        10'b1011001010: data <= 20'hff66e; 
        10'b1011001011: data <= 20'hff81d; 
        10'b1011001100: data <= 20'hffa25; 
        10'b1011001101: data <= 20'hffa83; 
        10'b1011001110: data <= 20'hffde7; 
        10'b1011001111: data <= 20'hffafb; 
        10'b1011010000: data <= 20'hffe32; 
        10'b1011010001: data <= 20'hffe10; 
        10'b1011010010: data <= 20'hfffeb; 
        10'b1011010011: data <= 20'hffd4b; 
        10'b1011010100: data <= 20'hffefc; 
        10'b1011010101: data <= 20'hffd5b; 
        10'b1011010110: data <= 20'hffc90; 
        10'b1011010111: data <= 20'hffd67; 
        10'b1011011000: data <= 20'hffcb0; 
        10'b1011011001: data <= 20'hffde8; 
        10'b1011011010: data <= 20'hffe7b; 
        10'b1011011011: data <= 20'h00028; 
        10'b1011011100: data <= 20'hfff75; 
        10'b1011011101: data <= 20'hffe57; 
        10'b1011011110: data <= 20'hfff55; 
        10'b1011011111: data <= 20'hfffe2; 
        10'b1011100000: data <= 20'hffe45; 
        10'b1011100001: data <= 20'h00033; 
        10'b1011100010: data <= 20'hffff0; 
        10'b1011100011: data <= 20'h0001d; 
        10'b1011100100: data <= 20'h00052; 
        10'b1011100101: data <= 20'hffefc; 
        10'b1011100110: data <= 20'hffdb4; 
        10'b1011100111: data <= 20'hffc3e; 
        10'b1011101000: data <= 20'hffe07; 
        10'b1011101001: data <= 20'hffef4; 
        10'b1011101010: data <= 20'hffec0; 
        10'b1011101011: data <= 20'hffd53; 
        10'b1011101100: data <= 20'h00059; 
        10'b1011101101: data <= 20'hfffef; 
        10'b1011101110: data <= 20'hffd5a; 
        10'b1011101111: data <= 20'hffde9; 
        10'b1011110000: data <= 20'hffca3; 
        10'b1011110001: data <= 20'h00027; 
        10'b1011110010: data <= 20'h0001c; 
        10'b1011110011: data <= 20'hfffd2; 
        10'b1011110100: data <= 20'hfffb8; 
        10'b1011110101: data <= 20'hffd8e; 
        10'b1011110110: data <= 20'hffcf5; 
        10'b1011110111: data <= 20'hffecb; 
        10'b1011111000: data <= 20'hffc98; 
        10'b1011111001: data <= 20'h000b5; 
        10'b1011111010: data <= 20'h000a3; 
        10'b1011111011: data <= 20'hffe05; 
        10'b1011111100: data <= 20'hfffcb; 
        10'b1011111101: data <= 20'hffd51; 
        10'b1011111110: data <= 20'h00077; 
        10'b1011111111: data <= 20'hffc82; 
        10'b1100000000: data <= 20'hfffd1; 
        10'b1100000001: data <= 20'hffe50; 
        10'b1100000010: data <= 20'hfff37; 
        10'b1100000011: data <= 20'hffd08; 
        10'b1100000100: data <= 20'hffec6; 
        10'b1100000101: data <= 20'hffe2d; 
        10'b1100000110: data <= 20'hffef5; 
        10'b1100000111: data <= 20'hffeb3; 
        10'b1100001000: data <= 20'hfff9d; 
        10'b1100001001: data <= 20'hffc5f; 
        10'b1100001010: data <= 20'hffe70; 
        10'b1100001011: data <= 20'h0001f; 
        10'b1100001100: data <= 20'hffc5f; 
        10'b1100001101: data <= 20'hffea0; 
        10'b1100001110: data <= 20'hfff7b; 
        10'b1100001111: data <= 20'hffe0f; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 15) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 21'h1ff991; 
        10'b0000000001: data <= 21'h000027; 
        10'b0000000010: data <= 21'h1ffccc; 
        10'b0000000011: data <= 21'h1ffab1; 
        10'b0000000100: data <= 21'h1ffcb5; 
        10'b0000000101: data <= 21'h1ffb0d; 
        10'b0000000110: data <= 21'h1ffdd5; 
        10'b0000000111: data <= 21'h1ffe2c; 
        10'b0000001000: data <= 21'h1ff964; 
        10'b0000001001: data <= 21'h1ffd50; 
        10'b0000001010: data <= 21'h1ff9dd; 
        10'b0000001011: data <= 21'h1ffbec; 
        10'b0000001100: data <= 21'h00013b; 
        10'b0000001101: data <= 21'h000114; 
        10'b0000001110: data <= 21'h1ff9bc; 
        10'b0000001111: data <= 21'h1ffdbd; 
        10'b0000010000: data <= 21'h1ffa2e; 
        10'b0000010001: data <= 21'h1ffa41; 
        10'b0000010010: data <= 21'h0001ab; 
        10'b0000010011: data <= 21'h00007a; 
        10'b0000010100: data <= 21'h1ffb3a; 
        10'b0000010101: data <= 21'h1ffdf4; 
        10'b0000010110: data <= 21'h1ffbc4; 
        10'b0000010111: data <= 21'h1ff8ff; 
        10'b0000011000: data <= 21'h1ff992; 
        10'b0000011001: data <= 21'h1ffd93; 
        10'b0000011010: data <= 21'h1fffaf; 
        10'b0000011011: data <= 21'h1ffe3c; 
        10'b0000011100: data <= 21'h1ffd46; 
        10'b0000011101: data <= 21'h1ffcd6; 
        10'b0000011110: data <= 21'h00018e; 
        10'b0000011111: data <= 21'h1ffe67; 
        10'b0000100000: data <= 21'h1ff9e6; 
        10'b0000100001: data <= 21'h1ff9b3; 
        10'b0000100010: data <= 21'h1ff974; 
        10'b0000100011: data <= 21'h1ffb0a; 
        10'b0000100100: data <= 21'h1ffb1c; 
        10'b0000100101: data <= 21'h1ffdb7; 
        10'b0000100110: data <= 21'h000011; 
        10'b0000100111: data <= 21'h1ffa21; 
        10'b0000101000: data <= 21'h1ffc3e; 
        10'b0000101001: data <= 21'h1ff9eb; 
        10'b0000101010: data <= 21'h1ffdd7; 
        10'b0000101011: data <= 21'h1ff900; 
        10'b0000101100: data <= 21'h1ffe25; 
        10'b0000101101: data <= 21'h1ffa24; 
        10'b0000101110: data <= 21'h1ffc0f; 
        10'b0000101111: data <= 21'h1ffa93; 
        10'b0000110000: data <= 21'h1ffdc8; 
        10'b0000110001: data <= 21'h1ffa4a; 
        10'b0000110010: data <= 21'h1ff950; 
        10'b0000110011: data <= 21'h1ff8ad; 
        10'b0000110100: data <= 21'h00005c; 
        10'b0000110101: data <= 21'h1ffe61; 
        10'b0000110110: data <= 21'h000078; 
        10'b0000110111: data <= 21'h1ffb97; 
        10'b0000111000: data <= 21'h1ffce0; 
        10'b0000111001: data <= 21'h1ff91c; 
        10'b0000111010: data <= 21'h1ff9c1; 
        10'b0000111011: data <= 21'h1ffff2; 
        10'b0000111100: data <= 21'h1ff95a; 
        10'b0000111101: data <= 21'h1ff9e9; 
        10'b0000111110: data <= 21'h1ffc8c; 
        10'b0000111111: data <= 21'h1ffd93; 
        10'b0001000000: data <= 21'h1fff5a; 
        10'b0001000001: data <= 21'h1ffc39; 
        10'b0001000010: data <= 21'h00039e; 
        10'b0001000011: data <= 21'h0002fc; 
        10'b0001000100: data <= 21'h00093e; 
        10'b0001000101: data <= 21'h00075f; 
        10'b0001000110: data <= 21'h0006bd; 
        10'b0001000111: data <= 21'h0002ad; 
        10'b0001001000: data <= 21'h000913; 
        10'b0001001001: data <= 21'h000318; 
        10'b0001001010: data <= 21'h0002a0; 
        10'b0001001011: data <= 21'h1ffb66; 
        10'b0001001100: data <= 21'h1fffdf; 
        10'b0001001101: data <= 21'h1ffddd; 
        10'b0001001110: data <= 21'h1ff69c; 
        10'b0001001111: data <= 21'h1ffcb1; 
        10'b0001010000: data <= 21'h1fff01; 
        10'b0001010001: data <= 21'h000243; 
        10'b0001010010: data <= 21'h1ffd4e; 
        10'b0001010011: data <= 21'h1ffc32; 
        10'b0001010100: data <= 21'h1ffb6c; 
        10'b0001010101: data <= 21'h1ffacd; 
        10'b0001010110: data <= 21'h1ffe83; 
        10'b0001010111: data <= 21'h1ffb3a; 
        10'b0001011000: data <= 21'h00014d; 
        10'b0001011001: data <= 21'h1ffa34; 
        10'b0001011010: data <= 21'h1ffde3; 
        10'b0001011011: data <= 21'h000001; 
        10'b0001011100: data <= 21'h0001a7; 
        10'b0001011101: data <= 21'h000eb8; 
        10'b0001011110: data <= 21'h001709; 
        10'b0001011111: data <= 21'h0016e1; 
        10'b0001100000: data <= 21'h0015e5; 
        10'b0001100001: data <= 21'h002036; 
        10'b0001100010: data <= 21'h001193; 
        10'b0001100011: data <= 21'h0007cc; 
        10'b0001100100: data <= 21'h000ecf; 
        10'b0001100101: data <= 21'h0006ca; 
        10'b0001100110: data <= 21'h1ff998; 
        10'b0001100111: data <= 21'h1ffe6a; 
        10'b0001101000: data <= 21'h1ff8b8; 
        10'b0001101001: data <= 21'h1ff779; 
        10'b0001101010: data <= 21'h1ff593; 
        10'b0001101011: data <= 21'h1ffad4; 
        10'b0001101100: data <= 21'h0000c3; 
        10'b0001101101: data <= 21'h000274; 
        10'b0001101110: data <= 21'h1ffa3d; 
        10'b0001101111: data <= 21'h1ffed7; 
        10'b0001110000: data <= 21'h1ffaf5; 
        10'b0001110001: data <= 21'h1ffc7f; 
        10'b0001110010: data <= 21'h0001c3; 
        10'b0001110011: data <= 21'h1ff879; 
        10'b0001110100: data <= 21'h1ff95c; 
        10'b0001110101: data <= 21'h1ffde3; 
        10'b0001110110: data <= 21'h000369; 
        10'b0001110111: data <= 21'h00034b; 
        10'b0001111000: data <= 21'h00097c; 
        10'b0001111001: data <= 21'h001c35; 
        10'b0001111010: data <= 21'h001c7e; 
        10'b0001111011: data <= 21'h0023ce; 
        10'b0001111100: data <= 21'h001e41; 
        10'b0001111101: data <= 21'h001800; 
        10'b0001111110: data <= 21'h0015ce; 
        10'b0001111111: data <= 21'h0009a2; 
        10'b0010000000: data <= 21'h000ce4; 
        10'b0010000001: data <= 21'h000bea; 
        10'b0010000010: data <= 21'h1ffc6e; 
        10'b0010000011: data <= 21'h1ff9fc; 
        10'b0010000100: data <= 21'h1ffb5b; 
        10'b0010000101: data <= 21'h1ff1d7; 
        10'b0010000110: data <= 21'h1feedc; 
        10'b0010000111: data <= 21'h1fef88; 
        10'b0010001000: data <= 21'h1ffde3; 
        10'b0010001001: data <= 21'h1ffde2; 
        10'b0010001010: data <= 21'h1ff91c; 
        10'b0010001011: data <= 21'h1ffeb3; 
        10'b0010001100: data <= 21'h000098; 
        10'b0010001101: data <= 21'h1ffdc4; 
        10'b0010001110: data <= 21'h1ffa91; 
        10'b0010001111: data <= 21'h1ff8bd; 
        10'b0010010000: data <= 21'h1ffa0a; 
        10'b0010010001: data <= 21'h1ffae0; 
        10'b0010010010: data <= 21'h000328; 
        10'b0010010011: data <= 21'h000dc9; 
        10'b0010010100: data <= 21'h00131d; 
        10'b0010010101: data <= 21'h0020b8; 
        10'b0010010110: data <= 21'h00243e; 
        10'b0010010111: data <= 21'h0025cd; 
        10'b0010011000: data <= 21'h0022a0; 
        10'b0010011001: data <= 21'h0026d3; 
        10'b0010011010: data <= 21'h0023f0; 
        10'b0010011011: data <= 21'h002157; 
        10'b0010011100: data <= 21'h002429; 
        10'b0010011101: data <= 21'h001d41; 
        10'b0010011110: data <= 21'h001522; 
        10'b0010011111: data <= 21'h1ff713; 
        10'b0010100000: data <= 21'h1ff761; 
        10'b0010100001: data <= 21'h1ff1eb; 
        10'b0010100010: data <= 21'h1ff1b0; 
        10'b0010100011: data <= 21'h1fe9ce; 
        10'b0010100100: data <= 21'h1ff66c; 
        10'b0010100101: data <= 21'h1ffa8e; 
        10'b0010100110: data <= 21'h0000e2; 
        10'b0010100111: data <= 21'h1ffbc3; 
        10'b0010101000: data <= 21'h1ffd1d; 
        10'b0010101001: data <= 21'h1ffad4; 
        10'b0010101010: data <= 21'h00012b; 
        10'b0010101011: data <= 21'h1ffd38; 
        10'b0010101100: data <= 21'h1ffc5b; 
        10'b0010101101: data <= 21'h00024f; 
        10'b0010101110: data <= 21'h000d7a; 
        10'b0010101111: data <= 21'h001a18; 
        10'b0010110000: data <= 21'h0013f2; 
        10'b0010110001: data <= 21'h0016a4; 
        10'b0010110010: data <= 21'h001ea7; 
        10'b0010110011: data <= 21'h00132b; 
        10'b0010110100: data <= 21'h00145f; 
        10'b0010110101: data <= 21'h001a4e; 
        10'b0010110110: data <= 21'h00173d; 
        10'b0010110111: data <= 21'h000ca4; 
        10'b0010111000: data <= 21'h000dfe; 
        10'b0010111001: data <= 21'h00039e; 
        10'b0010111010: data <= 21'h0002ab; 
        10'b0010111011: data <= 21'h1ff7c9; 
        10'b0010111100: data <= 21'h1ffa8a; 
        10'b0010111101: data <= 21'h1fee16; 
        10'b0010111110: data <= 21'h1fee39; 
        10'b0010111111: data <= 21'h1fe733; 
        10'b0011000000: data <= 21'h1ff13a; 
        10'b0011000001: data <= 21'h1ff7b9; 
        10'b0011000010: data <= 21'h00010d; 
        10'b0011000011: data <= 21'h1fff29; 
        10'b0011000100: data <= 21'h1ffc2c; 
        10'b0011000101: data <= 21'h0000c3; 
        10'b0011000110: data <= 21'h0000d6; 
        10'b0011000111: data <= 21'h1ffc82; 
        10'b0011001000: data <= 21'h00005a; 
        10'b0011001001: data <= 21'h00073f; 
        10'b0011001010: data <= 21'h00115e; 
        10'b0011001011: data <= 21'h001924; 
        10'b0011001100: data <= 21'h001492; 
        10'b0011001101: data <= 21'h001332; 
        10'b0011001110: data <= 21'h000756; 
        10'b0011001111: data <= 21'h0008ab; 
        10'b0011010000: data <= 21'h00017b; 
        10'b0011010001: data <= 21'h000d79; 
        10'b0011010010: data <= 21'h00109a; 
        10'b0011010011: data <= 21'h00037a; 
        10'b0011010100: data <= 21'h00023a; 
        10'b0011010101: data <= 21'h1feaf8; 
        10'b0011010110: data <= 21'h1ff8df; 
        10'b0011010111: data <= 21'h1ffa11; 
        10'b0011011000: data <= 21'h1ff944; 
        10'b0011011001: data <= 21'h1ff81f; 
        10'b0011011010: data <= 21'h1ffa20; 
        10'b0011011011: data <= 21'h1feb98; 
        10'b0011011100: data <= 21'h1ff1dd; 
        10'b0011011101: data <= 21'h1ffbaf; 
        10'b0011011110: data <= 21'h1ffa8f; 
        10'b0011011111: data <= 21'h1ff95e; 
        10'b0011100000: data <= 21'h1ffe7b; 
        10'b0011100001: data <= 21'h0000ff; 
        10'b0011100010: data <= 21'h1ffd2d; 
        10'b0011100011: data <= 21'h0000ea; 
        10'b0011100100: data <= 21'h0003cb; 
        10'b0011100101: data <= 21'h000bc2; 
        10'b0011100110: data <= 21'h000881; 
        10'b0011100111: data <= 21'h000c01; 
        10'b0011101000: data <= 21'h000c28; 
        10'b0011101001: data <= 21'h000d86; 
        10'b0011101010: data <= 21'h000d97; 
        10'b0011101011: data <= 21'h000f82; 
        10'b0011101100: data <= 21'h000938; 
        10'b0011101101: data <= 21'h000b04; 
        10'b0011101110: data <= 21'h001d0f; 
        10'b0011101111: data <= 21'h001056; 
        10'b0011110000: data <= 21'h1ffdfc; 
        10'b0011110001: data <= 21'h1ff806; 
        10'b0011110010: data <= 21'h1fffcb; 
        10'b0011110011: data <= 21'h000673; 
        10'b0011110100: data <= 21'h000027; 
        10'b0011110101: data <= 21'h1ffb8c; 
        10'b0011110110: data <= 21'h1ff428; 
        10'b0011110111: data <= 21'h1fe82f; 
        10'b0011111000: data <= 21'h1fedba; 
        10'b0011111001: data <= 21'h1ff863; 
        10'b0011111010: data <= 21'h1ffc70; 
        10'b0011111011: data <= 21'h1ffa27; 
        10'b0011111100: data <= 21'h1ffafa; 
        10'b0011111101: data <= 21'h1ffec5; 
        10'b0011111110: data <= 21'h1fffba; 
        10'b0011111111: data <= 21'h00030c; 
        10'b0100000000: data <= 21'h0005e9; 
        10'b0100000001: data <= 21'h000d2b; 
        10'b0100000010: data <= 21'h00049d; 
        10'b0100000011: data <= 21'h0000e4; 
        10'b0100000100: data <= 21'h1ffb73; 
        10'b0100000101: data <= 21'h000716; 
        10'b0100000110: data <= 21'h000581; 
        10'b0100000111: data <= 21'h00071b; 
        10'b0100001000: data <= 21'h0001d8; 
        10'b0100001001: data <= 21'h1fff43; 
        10'b0100001010: data <= 21'h0012f6; 
        10'b0100001011: data <= 21'h001481; 
        10'b0100001100: data <= 21'h000712; 
        10'b0100001101: data <= 21'h00008a; 
        10'b0100001110: data <= 21'h1ffe19; 
        10'b0100001111: data <= 21'h1fffd4; 
        10'b0100010000: data <= 21'h1fff24; 
        10'b0100010001: data <= 21'h1fff8b; 
        10'b0100010010: data <= 21'h1ff87a; 
        10'b0100010011: data <= 21'h1febbf; 
        10'b0100010100: data <= 21'h1feeb7; 
        10'b0100010101: data <= 21'h1ffa60; 
        10'b0100010110: data <= 21'h0000e5; 
        10'b0100010111: data <= 21'h1ff979; 
        10'b0100011000: data <= 21'h000146; 
        10'b0100011001: data <= 21'h1ffe85; 
        10'b0100011010: data <= 21'h1ffd01; 
        10'b0100011011: data <= 21'h1ffbc0; 
        10'b0100011100: data <= 21'h0000e6; 
        10'b0100011101: data <= 21'h1ffcc9; 
        10'b0100011110: data <= 21'h1ff96b; 
        10'b0100011111: data <= 21'h1fe009; 
        10'b0100100000: data <= 21'h1fe367; 
        10'b0100100001: data <= 21'h1fea65; 
        10'b0100100010: data <= 21'h1fdef9; 
        10'b0100100011: data <= 21'h1fdb60; 
        10'b0100100100: data <= 21'h1fd563; 
        10'b0100100101: data <= 21'h1fd025; 
        10'b0100100110: data <= 21'h1febe8; 
        10'b0100100111: data <= 21'h0003a5; 
        10'b0100101000: data <= 21'h00052c; 
        10'b0100101001: data <= 21'h0000de; 
        10'b0100101010: data <= 21'h0002a9; 
        10'b0100101011: data <= 21'h1ffc1d; 
        10'b0100101100: data <= 21'h1ffd2b; 
        10'b0100101101: data <= 21'h1ffc19; 
        10'b0100101110: data <= 21'h1ff5f8; 
        10'b0100101111: data <= 21'h1fe8b5; 
        10'b0100110000: data <= 21'h1ff334; 
        10'b0100110001: data <= 21'h1fff75; 
        10'b0100110010: data <= 21'h1fff6a; 
        10'b0100110011: data <= 21'h1ffa9e; 
        10'b0100110100: data <= 21'h1ff957; 
        10'b0100110101: data <= 21'h0001a4; 
        10'b0100110110: data <= 21'h1fff52; 
        10'b0100110111: data <= 21'h1ff9e2; 
        10'b0100111000: data <= 21'h1ff404; 
        10'b0100111001: data <= 21'h1fe5cf; 
        10'b0100111010: data <= 21'h1fd30e; 
        10'b0100111011: data <= 21'h1fc0a1; 
        10'b0100111100: data <= 21'h1fc31f; 
        10'b0100111101: data <= 21'h1fb84e; 
        10'b0100111110: data <= 21'h1fb819; 
        10'b0100111111: data <= 21'h1fbe5e; 
        10'b0101000000: data <= 21'h1fba55; 
        10'b0101000001: data <= 21'h1fab1c; 
        10'b0101000010: data <= 21'h1fbeb3; 
        10'b0101000011: data <= 21'h1fe0c4; 
        10'b0101000100: data <= 21'h1ff52c; 
        10'b0101000101: data <= 21'h1ff6b0; 
        10'b0101000110: data <= 21'h1ff70d; 
        10'b0101000111: data <= 21'h1ffe36; 
        10'b0101001000: data <= 21'h1ffa9f; 
        10'b0101001001: data <= 21'h1ffa64; 
        10'b0101001010: data <= 21'h1ff12a; 
        10'b0101001011: data <= 21'h1ff5d9; 
        10'b0101001100: data <= 21'h1ffe28; 
        10'b0101001101: data <= 21'h1ffc7e; 
        10'b0101001110: data <= 21'h1ffa72; 
        10'b0101001111: data <= 21'h1ffe75; 
        10'b0101010000: data <= 21'h1ffdb2; 
        10'b0101010001: data <= 21'h1ffe18; 
        10'b0101010010: data <= 21'h0000aa; 
        10'b0101010011: data <= 21'h1ffd35; 
        10'b0101010100: data <= 21'h1ff319; 
        10'b0101010101: data <= 21'h1fd901; 
        10'b0101010110: data <= 21'h1fb423; 
        10'b0101010111: data <= 21'h1fa32d; 
        10'b0101011000: data <= 21'h1fa96c; 
        10'b0101011001: data <= 21'h1fadf2; 
        10'b0101011010: data <= 21'h1fb505; 
        10'b0101011011: data <= 21'h1fb9d6; 
        10'b0101011100: data <= 21'h1fba09; 
        10'b0101011101: data <= 21'h1fb734; 
        10'b0101011110: data <= 21'h1fc435; 
        10'b0101011111: data <= 21'h1fd81f; 
        10'b0101100000: data <= 21'h1fe4a3; 
        10'b0101100001: data <= 21'h1fe76c; 
        10'b0101100010: data <= 21'h1ff39d; 
        10'b0101100011: data <= 21'h00000e; 
        10'b0101100100: data <= 21'h1fffc3; 
        10'b0101100101: data <= 21'h1ff90e; 
        10'b0101100110: data <= 21'h1ff036; 
        10'b0101100111: data <= 21'h1fe7fc; 
        10'b0101101000: data <= 21'h1ffd13; 
        10'b0101101001: data <= 21'h1ffc06; 
        10'b0101101010: data <= 21'h0001c9; 
        10'b0101101011: data <= 21'h1ffe18; 
        10'b0101101100: data <= 21'h1ffb2c; 
        10'b0101101101: data <= 21'h1ffcd6; 
        10'b0101101110: data <= 21'h0001aa; 
        10'b0101101111: data <= 21'h1ffb02; 
        10'b0101110000: data <= 21'h1feb1e; 
        10'b0101110001: data <= 21'h1fced3; 
        10'b0101110010: data <= 21'h1fb1f5; 
        10'b0101110011: data <= 21'h1fb85d; 
        10'b0101110100: data <= 21'h1fbd23; 
        10'b0101110101: data <= 21'h1fd20b; 
        10'b0101110110: data <= 21'h1fdf6e; 
        10'b0101110111: data <= 21'h1ff0c0; 
        10'b0101111000: data <= 21'h1fe7e0; 
        10'b0101111001: data <= 21'h1ff507; 
        10'b0101111010: data <= 21'h1fe473; 
        10'b0101111011: data <= 21'h1fe3e3; 
        10'b0101111100: data <= 21'h1fdea8; 
        10'b0101111101: data <= 21'h1fe7ee; 
        10'b0101111110: data <= 21'h1ff2bd; 
        10'b0101111111: data <= 21'h1ffd76; 
        10'b0110000000: data <= 21'h1ffc1c; 
        10'b0110000001: data <= 21'h1ff774; 
        10'b0110000010: data <= 21'h1fec26; 
        10'b0110000011: data <= 21'h1fedee; 
        10'b0110000100: data <= 21'h1ff6dc; 
        10'b0110000101: data <= 21'h00024b; 
        10'b0110000110: data <= 21'h1ffcf2; 
        10'b0110000111: data <= 21'h1fffcc; 
        10'b0110001000: data <= 21'h00010b; 
        10'b0110001001: data <= 21'h1ffe57; 
        10'b0110001010: data <= 21'h00002c; 
        10'b0110001011: data <= 21'h1ffbcc; 
        10'b0110001100: data <= 21'h1ff801; 
        10'b0110001101: data <= 21'h1fdec9; 
        10'b0110001110: data <= 21'h1fd5fa; 
        10'b0110001111: data <= 21'h1fddbe; 
        10'b0110010000: data <= 21'h1ff242; 
        10'b0110010001: data <= 21'h1ffda1; 
        10'b0110010010: data <= 21'h000891; 
        10'b0110010011: data <= 21'h000b56; 
        10'b0110010100: data <= 21'h000d73; 
        10'b0110010101: data <= 21'h0014ee; 
        10'b0110010110: data <= 21'h00016d; 
        10'b0110010111: data <= 21'h1ff299; 
        10'b0110011000: data <= 21'h1ff60b; 
        10'b0110011001: data <= 21'h1feebf; 
        10'b0110011010: data <= 21'h1ffd19; 
        10'b0110011011: data <= 21'h1ff4e7; 
        10'b0110011100: data <= 21'h1ffc7e; 
        10'b0110011101: data <= 21'h1ff337; 
        10'b0110011110: data <= 21'h1fe905; 
        10'b0110011111: data <= 21'h1fef4b; 
        10'b0110100000: data <= 21'h1ffcbb; 
        10'b0110100001: data <= 21'h000822; 
        10'b0110100010: data <= 21'h00093b; 
        10'b0110100011: data <= 21'h1ffadf; 
        10'b0110100100: data <= 21'h1ffc68; 
        10'b0110100101: data <= 21'h1ffd29; 
        10'b0110100110: data <= 21'h1ffc4b; 
        10'b0110100111: data <= 21'h000797; 
        10'b0110101000: data <= 21'h0003ad; 
        10'b0110101001: data <= 21'h0001a9; 
        10'b0110101010: data <= 21'h0008fc; 
        10'b0110101011: data <= 21'h000a86; 
        10'b0110101100: data <= 21'h00138e; 
        10'b0110101101: data <= 21'h000dd2; 
        10'b0110101110: data <= 21'h001092; 
        10'b0110101111: data <= 21'h0009be; 
        10'b0110110000: data <= 21'h0008a0; 
        10'b0110110001: data <= 21'h001439; 
        10'b0110110010: data <= 21'h000181; 
        10'b0110110011: data <= 21'h0007f0; 
        10'b0110110100: data <= 21'h000122; 
        10'b0110110101: data <= 21'h1feff6; 
        10'b0110110110: data <= 21'h1ff0be; 
        10'b0110110111: data <= 21'h1ff6a4; 
        10'b0110111000: data <= 21'h1ff92d; 
        10'b0110111001: data <= 21'h1ff5ae; 
        10'b0110111010: data <= 21'h1feb2e; 
        10'b0110111011: data <= 21'h1ff54a; 
        10'b0110111100: data <= 21'h000667; 
        10'b0110111101: data <= 21'h000ae9; 
        10'b0110111110: data <= 21'h0005e5; 
        10'b0110111111: data <= 21'h1ffa2a; 
        10'b0111000000: data <= 21'h1ffb8c; 
        10'b0111000001: data <= 21'h1ff915; 
        10'b0111000010: data <= 21'h1ff828; 
        10'b0111000011: data <= 21'h000813; 
        10'b0111000100: data <= 21'h0010f1; 
        10'b0111000101: data <= 21'h001ba7; 
        10'b0111000110: data <= 21'h001c2c; 
        10'b0111000111: data <= 21'h0010c4; 
        10'b0111001000: data <= 21'h0006f4; 
        10'b0111001001: data <= 21'h000e76; 
        10'b0111001010: data <= 21'h000d6e; 
        10'b0111001011: data <= 21'h000c44; 
        10'b0111001100: data <= 21'h001945; 
        10'b0111001101: data <= 21'h001641; 
        10'b0111001110: data <= 21'h0004ab; 
        10'b0111001111: data <= 21'h1ffd57; 
        10'b0111010000: data <= 21'h1fffe6; 
        10'b0111010001: data <= 21'h1ff596; 
        10'b0111010010: data <= 21'h1ff6e4; 
        10'b0111010011: data <= 21'h1ff006; 
        10'b0111010100: data <= 21'h1ffa52; 
        10'b0111010101: data <= 21'h0000dd; 
        10'b0111010110: data <= 21'h000384; 
        10'b0111010111: data <= 21'h00076c; 
        10'b0111011000: data <= 21'h001799; 
        10'b0111011001: data <= 21'h001d3a; 
        10'b0111011010: data <= 21'h0004e5; 
        10'b0111011011: data <= 21'h1ffb6e; 
        10'b0111011100: data <= 21'h1ffc39; 
        10'b0111011101: data <= 21'h000155; 
        10'b0111011110: data <= 21'h1ffd0e; 
        10'b0111011111: data <= 21'h0009ca; 
        10'b0111100000: data <= 21'h001ced; 
        10'b0111100001: data <= 21'h00284e; 
        10'b0111100010: data <= 21'h0024d5; 
        10'b0111100011: data <= 21'h00193d; 
        10'b0111100100: data <= 21'h001190; 
        10'b0111100101: data <= 21'h00154c; 
        10'b0111100110: data <= 21'h0020bf; 
        10'b0111100111: data <= 21'h001ad7; 
        10'b0111101000: data <= 21'h001ec8; 
        10'b0111101001: data <= 21'h000e67; 
        10'b0111101010: data <= 21'h00076b; 
        10'b0111101011: data <= 21'h000a01; 
        10'b0111101100: data <= 21'h000a1b; 
        10'b0111101101: data <= 21'h1ffe70; 
        10'b0111101110: data <= 21'h00068e; 
        10'b0111101111: data <= 21'h1ffbd2; 
        10'b0111110000: data <= 21'h000c17; 
        10'b0111110001: data <= 21'h000ce6; 
        10'b0111110010: data <= 21'h000995; 
        10'b0111110011: data <= 21'h000d49; 
        10'b0111110100: data <= 21'h0025cf; 
        10'b0111110101: data <= 21'h0020cb; 
        10'b0111110110: data <= 21'h00077c; 
        10'b0111110111: data <= 21'h0000fe; 
        10'b0111111000: data <= 21'h1fff26; 
        10'b0111111001: data <= 21'h1fff8a; 
        10'b0111111010: data <= 21'h1ff60b; 
        10'b0111111011: data <= 21'h0002a2; 
        10'b0111111100: data <= 21'h001f5a; 
        10'b0111111101: data <= 21'h0034fa; 
        10'b0111111110: data <= 21'h0031d5; 
        10'b0111111111: data <= 21'h0023df; 
        10'b1000000000: data <= 21'h0017ed; 
        10'b1000000001: data <= 21'h001a99; 
        10'b1000000010: data <= 21'h0028a6; 
        10'b1000000011: data <= 21'h0024ba; 
        10'b1000000100: data <= 21'h003a81; 
        10'b1000000101: data <= 21'h002ab4; 
        10'b1000000110: data <= 21'h00254b; 
        10'b1000000111: data <= 21'h001226; 
        10'b1000001000: data <= 21'h000c7d; 
        10'b1000001001: data <= 21'h0016f1; 
        10'b1000001010: data <= 21'h000ecd; 
        10'b1000001011: data <= 21'h000a14; 
        10'b1000001100: data <= 21'h001b11; 
        10'b1000001101: data <= 21'h001bf5; 
        10'b1000001110: data <= 21'h001e79; 
        10'b1000001111: data <= 21'h002843; 
        10'b1000010000: data <= 21'h0031f7; 
        10'b1000010001: data <= 21'h001cd0; 
        10'b1000010010: data <= 21'h1ffd3c; 
        10'b1000010011: data <= 21'h1ffa10; 
        10'b1000010100: data <= 21'h1ffaf1; 
        10'b1000010101: data <= 21'h1ffb46; 
        10'b1000010110: data <= 21'h1ff90c; 
        10'b1000010111: data <= 21'h1fffe2; 
        10'b1000011000: data <= 21'h00113a; 
        10'b1000011001: data <= 21'h00202e; 
        10'b1000011010: data <= 21'h0028a4; 
        10'b1000011011: data <= 21'h00233d; 
        10'b1000011100: data <= 21'h002088; 
        10'b1000011101: data <= 21'h00226f; 
        10'b1000011110: data <= 21'h0020f5; 
        10'b1000011111: data <= 21'h002300; 
        10'b1000100000: data <= 21'h00272c; 
        10'b1000100001: data <= 21'h001e22; 
        10'b1000100010: data <= 21'h001384; 
        10'b1000100011: data <= 21'h000941; 
        10'b1000100100: data <= 21'h000e5f; 
        10'b1000100101: data <= 21'h0018f6; 
        10'b1000100110: data <= 21'h000c0f; 
        10'b1000100111: data <= 21'h000bc8; 
        10'b1000101000: data <= 21'h00141c; 
        10'b1000101001: data <= 21'h001917; 
        10'b1000101010: data <= 21'h0020c4; 
        10'b1000101011: data <= 21'h002325; 
        10'b1000101100: data <= 21'h001e4a; 
        10'b1000101101: data <= 21'h000fdd; 
        10'b1000101110: data <= 21'h000157; 
        10'b1000101111: data <= 21'h00005e; 
        10'b1000110000: data <= 21'h1ff9b9; 
        10'b1000110001: data <= 21'h1fff82; 
        10'b1000110010: data <= 21'h1ffe53; 
        10'b1000110011: data <= 21'h1ff760; 
        10'b1000110100: data <= 21'h000f4a; 
        10'b1000110101: data <= 21'h0012e2; 
        10'b1000110110: data <= 21'h001d50; 
        10'b1000110111: data <= 21'h0028c4; 
        10'b1000111000: data <= 21'h0026b9; 
        10'b1000111001: data <= 21'h0019a7; 
        10'b1000111010: data <= 21'h0018ab; 
        10'b1000111011: data <= 21'h002949; 
        10'b1000111100: data <= 21'h0016f5; 
        10'b1000111101: data <= 21'h000799; 
        10'b1000111110: data <= 21'h000518; 
        10'b1000111111: data <= 21'h000641; 
        10'b1001000000: data <= 21'h000818; 
        10'b1001000001: data <= 21'h00005e; 
        10'b1001000010: data <= 21'h0011da; 
        10'b1001000011: data <= 21'h001be0; 
        10'b1001000100: data <= 21'h0012ea; 
        10'b1001000101: data <= 21'h001ae7; 
        10'b1001000110: data <= 21'h002577; 
        10'b1001000111: data <= 21'h002081; 
        10'b1001001000: data <= 21'h001765; 
        10'b1001001001: data <= 21'h000b18; 
        10'b1001001010: data <= 21'h1fffdc; 
        10'b1001001011: data <= 21'h1ffef8; 
        10'b1001001100: data <= 21'h1ffd8a; 
        10'b1001001101: data <= 21'h1ffa02; 
        10'b1001001110: data <= 21'h1ffeed; 
        10'b1001001111: data <= 21'h1ffc8d; 
        10'b1001010000: data <= 21'h000332; 
        10'b1001010001: data <= 21'h00081f; 
        10'b1001010010: data <= 21'h001455; 
        10'b1001010011: data <= 21'h0016d8; 
        10'b1001010100: data <= 21'h001423; 
        10'b1001010101: data <= 21'h001922; 
        10'b1001010110: data <= 21'h00163c; 
        10'b1001010111: data <= 21'h0015d5; 
        10'b1001011000: data <= 21'h000892; 
        10'b1001011001: data <= 21'h000415; 
        10'b1001011010: data <= 21'h1ffdc9; 
        10'b1001011011: data <= 21'h0000f2; 
        10'b1001011100: data <= 21'h000adc; 
        10'b1001011101: data <= 21'h000be6; 
        10'b1001011110: data <= 21'h001a11; 
        10'b1001011111: data <= 21'h001b6c; 
        10'b1001100000: data <= 21'h000c07; 
        10'b1001100001: data <= 21'h001ae3; 
        10'b1001100010: data <= 21'h002137; 
        10'b1001100011: data <= 21'h0025d6; 
        10'b1001100100: data <= 21'h0012a5; 
        10'b1001100101: data <= 21'h000765; 
        10'b1001100110: data <= 21'h0001b5; 
        10'b1001100111: data <= 21'h1fff2b; 
        10'b1001101000: data <= 21'h1ff9ad; 
        10'b1001101001: data <= 21'h1ffe4e; 
        10'b1001101010: data <= 21'h1ffa8d; 
        10'b1001101011: data <= 21'h0001cb; 
        10'b1001101100: data <= 21'h000665; 
        10'b1001101101: data <= 21'h00024f; 
        10'b1001101110: data <= 21'h000dd7; 
        10'b1001101111: data <= 21'h000c24; 
        10'b1001110000: data <= 21'h000b51; 
        10'b1001110001: data <= 21'h000fe5; 
        10'b1001110010: data <= 21'h000fc9; 
        10'b1001110011: data <= 21'h0012b6; 
        10'b1001110100: data <= 21'h000207; 
        10'b1001110101: data <= 21'h1ff138; 
        10'b1001110110: data <= 21'h1fed64; 
        10'b1001110111: data <= 21'h1ff576; 
        10'b1001111000: data <= 21'h1ff613; 
        10'b1001111001: data <= 21'h0007b6; 
        10'b1001111010: data <= 21'h00183b; 
        10'b1001111011: data <= 21'h001eef; 
        10'b1001111100: data <= 21'h001c20; 
        10'b1001111101: data <= 21'h001ae9; 
        10'b1001111110: data <= 21'h00175e; 
        10'b1001111111: data <= 21'h0019c5; 
        10'b1010000000: data <= 21'h000993; 
        10'b1010000001: data <= 21'h1ffef1; 
        10'b1010000010: data <= 21'h1ffe5d; 
        10'b1010000011: data <= 21'h1ffb83; 
        10'b1010000100: data <= 21'h1ffe77; 
        10'b1010000101: data <= 21'h1ffea8; 
        10'b1010000110: data <= 21'h1ffd36; 
        10'b1010000111: data <= 21'h1ffcc0; 
        10'b1010001000: data <= 21'h1ffc60; 
        10'b1010001001: data <= 21'h1ff8cd; 
        10'b1010001010: data <= 21'h1ff72a; 
        10'b1010001011: data <= 21'h1ff854; 
        10'b1010001100: data <= 21'h1ff36a; 
        10'b1010001101: data <= 21'h1ff89e; 
        10'b1010001110: data <= 21'h1ffb11; 
        10'b1010001111: data <= 21'h00065d; 
        10'b1010010000: data <= 21'h000096; 
        10'b1010010001: data <= 21'h1ff618; 
        10'b1010010010: data <= 21'h1ff298; 
        10'b1010010011: data <= 21'h1fee80; 
        10'b1010010100: data <= 21'h1fed00; 
        10'b1010010101: data <= 21'h1ff61a; 
        10'b1010010110: data <= 21'h0003e1; 
        10'b1010010111: data <= 21'h001837; 
        10'b1010011000: data <= 21'h001532; 
        10'b1010011001: data <= 21'h0019f5; 
        10'b1010011010: data <= 21'h0012a0; 
        10'b1010011011: data <= 21'h00071e; 
        10'b1010011100: data <= 21'h00044e; 
        10'b1010011101: data <= 21'h0002bf; 
        10'b1010011110: data <= 21'h1fff65; 
        10'b1010011111: data <= 21'h1ffcab; 
        10'b1010100000: data <= 21'h1ffd9f; 
        10'b1010100001: data <= 21'h1ffb17; 
        10'b1010100010: data <= 21'h1fffc2; 
        10'b1010100011: data <= 21'h1fff2a; 
        10'b1010100100: data <= 21'h1ffacd; 
        10'b1010100101: data <= 21'h1ff272; 
        10'b1010100110: data <= 21'h1fe5d0; 
        10'b1010100111: data <= 21'h1fec6c; 
        10'b1010101000: data <= 21'h1febd9; 
        10'b1010101001: data <= 21'h1fea7e; 
        10'b1010101010: data <= 21'h1feaa9; 
        10'b1010101011: data <= 21'h1fefa8; 
        10'b1010101100: data <= 21'h1fef87; 
        10'b1010101101: data <= 21'h1ff70e; 
        10'b1010101110: data <= 21'h1ff453; 
        10'b1010101111: data <= 21'h1fef5c; 
        10'b1010110000: data <= 21'h1ff034; 
        10'b1010110001: data <= 21'h1ff39d; 
        10'b1010110010: data <= 21'h1ff0db; 
        10'b1010110011: data <= 21'h1ff7d2; 
        10'b1010110100: data <= 21'h1ff8c4; 
        10'b1010110101: data <= 21'h1ff8cf; 
        10'b1010110110: data <= 21'h1ffbcb; 
        10'b1010110111: data <= 21'h1ffcac; 
        10'b1010111000: data <= 21'h1fff80; 
        10'b1010111001: data <= 21'h0002b3; 
        10'b1010111010: data <= 21'h1ffa59; 
        10'b1010111011: data <= 21'h1ffa82; 
        10'b1010111100: data <= 21'h1fffc4; 
        10'b1010111101: data <= 21'h1ff8ec; 
        10'b1010111110: data <= 21'h1ffc66; 
        10'b1010111111: data <= 21'h1ffbac; 
        10'b1011000000: data <= 21'h1ffa6a; 
        10'b1011000001: data <= 21'h1ff673; 
        10'b1011000010: data <= 21'h1ff34a; 
        10'b1011000011: data <= 21'h1feca6; 
        10'b1011000100: data <= 21'h1fea85; 
        10'b1011000101: data <= 21'h1fec14; 
        10'b1011000110: data <= 21'h1fedf6; 
        10'b1011000111: data <= 21'h1fe908; 
        10'b1011001000: data <= 21'h1ff09d; 
        10'b1011001001: data <= 21'h1ff192; 
        10'b1011001010: data <= 21'h1fecdb; 
        10'b1011001011: data <= 21'h1ff03a; 
        10'b1011001100: data <= 21'h1ff44b; 
        10'b1011001101: data <= 21'h1ff506; 
        10'b1011001110: data <= 21'h1ffbce; 
        10'b1011001111: data <= 21'h1ff5f6; 
        10'b1011010000: data <= 21'h1ffc65; 
        10'b1011010001: data <= 21'h1ffc1f; 
        10'b1011010010: data <= 21'h1fffd5; 
        10'b1011010011: data <= 21'h1ffa96; 
        10'b1011010100: data <= 21'h1ffdf8; 
        10'b1011010101: data <= 21'h1ffab5; 
        10'b1011010110: data <= 21'h1ff920; 
        10'b1011010111: data <= 21'h1ffacd; 
        10'b1011011000: data <= 21'h1ff95f; 
        10'b1011011001: data <= 21'h1ffbd0; 
        10'b1011011010: data <= 21'h1ffcf5; 
        10'b1011011011: data <= 21'h000050; 
        10'b1011011100: data <= 21'h1ffeea; 
        10'b1011011101: data <= 21'h1ffcae; 
        10'b1011011110: data <= 21'h1ffeab; 
        10'b1011011111: data <= 21'h1fffc4; 
        10'b1011100000: data <= 21'h1ffc8a; 
        10'b1011100001: data <= 21'h000066; 
        10'b1011100010: data <= 21'h1fffe0; 
        10'b1011100011: data <= 21'h00003a; 
        10'b1011100100: data <= 21'h0000a3; 
        10'b1011100101: data <= 21'h1ffdf8; 
        10'b1011100110: data <= 21'h1ffb69; 
        10'b1011100111: data <= 21'h1ff87d; 
        10'b1011101000: data <= 21'h1ffc0d; 
        10'b1011101001: data <= 21'h1ffde8; 
        10'b1011101010: data <= 21'h1ffd80; 
        10'b1011101011: data <= 21'h1ffaa5; 
        10'b1011101100: data <= 21'h0000b2; 
        10'b1011101101: data <= 21'h1fffdf; 
        10'b1011101110: data <= 21'h1ffab3; 
        10'b1011101111: data <= 21'h1ffbd2; 
        10'b1011110000: data <= 21'h1ff947; 
        10'b1011110001: data <= 21'h00004e; 
        10'b1011110010: data <= 21'h000037; 
        10'b1011110011: data <= 21'h1fffa4; 
        10'b1011110100: data <= 21'h1fff6f; 
        10'b1011110101: data <= 21'h1ffb1d; 
        10'b1011110110: data <= 21'h1ff9e9; 
        10'b1011110111: data <= 21'h1ffd96; 
        10'b1011111000: data <= 21'h1ff930; 
        10'b1011111001: data <= 21'h000169; 
        10'b1011111010: data <= 21'h000146; 
        10'b1011111011: data <= 21'h1ffc09; 
        10'b1011111100: data <= 21'h1fff95; 
        10'b1011111101: data <= 21'h1ffaa3; 
        10'b1011111110: data <= 21'h0000ef; 
        10'b1011111111: data <= 21'h1ff904; 
        10'b1100000000: data <= 21'h1fffa1; 
        10'b1100000001: data <= 21'h1ffc9f; 
        10'b1100000010: data <= 21'h1ffe6e; 
        10'b1100000011: data <= 21'h1ffa10; 
        10'b1100000100: data <= 21'h1ffd8d; 
        10'b1100000101: data <= 21'h1ffc5a; 
        10'b1100000110: data <= 21'h1ffdea; 
        10'b1100000111: data <= 21'h1ffd65; 
        10'b1100001000: data <= 21'h1fff39; 
        10'b1100001001: data <= 21'h1ff8bf; 
        10'b1100001010: data <= 21'h1ffce1; 
        10'b1100001011: data <= 21'h00003d; 
        10'b1100001100: data <= 21'h1ff8bd; 
        10'b1100001101: data <= 21'h1ffd40; 
        10'b1100001110: data <= 21'h1ffef6; 
        10'b1100001111: data <= 21'h1ffc1d; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 16) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 22'h3ff323; 
        10'b0000000001: data <= 22'h00004d; 
        10'b0000000010: data <= 22'h3ff999; 
        10'b0000000011: data <= 22'h3ff562; 
        10'b0000000100: data <= 22'h3ff96b; 
        10'b0000000101: data <= 22'h3ff61a; 
        10'b0000000110: data <= 22'h3ffbaa; 
        10'b0000000111: data <= 22'h3ffc59; 
        10'b0000001000: data <= 22'h3ff2c8; 
        10'b0000001001: data <= 22'h3ffaa0; 
        10'b0000001010: data <= 22'h3ff3bb; 
        10'b0000001011: data <= 22'h3ff7d9; 
        10'b0000001100: data <= 22'h000277; 
        10'b0000001101: data <= 22'h000228; 
        10'b0000001110: data <= 22'h3ff378; 
        10'b0000001111: data <= 22'h3ffb7b; 
        10'b0000010000: data <= 22'h3ff45d; 
        10'b0000010001: data <= 22'h3ff483; 
        10'b0000010010: data <= 22'h000355; 
        10'b0000010011: data <= 22'h0000f3; 
        10'b0000010100: data <= 22'h3ff673; 
        10'b0000010101: data <= 22'h3ffbe8; 
        10'b0000010110: data <= 22'h3ff787; 
        10'b0000010111: data <= 22'h3ff1ff; 
        10'b0000011000: data <= 22'h3ff323; 
        10'b0000011001: data <= 22'h3ffb26; 
        10'b0000011010: data <= 22'h3fff5e; 
        10'b0000011011: data <= 22'h3ffc79; 
        10'b0000011100: data <= 22'h3ffa8c; 
        10'b0000011101: data <= 22'h3ff9ad; 
        10'b0000011110: data <= 22'h00031c; 
        10'b0000011111: data <= 22'h3ffccd; 
        10'b0000100000: data <= 22'h3ff3cc; 
        10'b0000100001: data <= 22'h3ff365; 
        10'b0000100010: data <= 22'h3ff2e8; 
        10'b0000100011: data <= 22'h3ff613; 
        10'b0000100100: data <= 22'h3ff637; 
        10'b0000100101: data <= 22'h3ffb6e; 
        10'b0000100110: data <= 22'h000021; 
        10'b0000100111: data <= 22'h3ff442; 
        10'b0000101000: data <= 22'h3ff87c; 
        10'b0000101001: data <= 22'h3ff3d5; 
        10'b0000101010: data <= 22'h3ffbae; 
        10'b0000101011: data <= 22'h3ff201; 
        10'b0000101100: data <= 22'h3ffc4a; 
        10'b0000101101: data <= 22'h3ff448; 
        10'b0000101110: data <= 22'h3ff81d; 
        10'b0000101111: data <= 22'h3ff525; 
        10'b0000110000: data <= 22'h3ffb91; 
        10'b0000110001: data <= 22'h3ff495; 
        10'b0000110010: data <= 22'h3ff29f; 
        10'b0000110011: data <= 22'h3ff15b; 
        10'b0000110100: data <= 22'h0000b9; 
        10'b0000110101: data <= 22'h3ffcc2; 
        10'b0000110110: data <= 22'h0000f0; 
        10'b0000110111: data <= 22'h3ff72f; 
        10'b0000111000: data <= 22'h3ff9c0; 
        10'b0000111001: data <= 22'h3ff238; 
        10'b0000111010: data <= 22'h3ff382; 
        10'b0000111011: data <= 22'h3fffe4; 
        10'b0000111100: data <= 22'h3ff2b3; 
        10'b0000111101: data <= 22'h3ff3d2; 
        10'b0000111110: data <= 22'h3ff919; 
        10'b0000111111: data <= 22'h3ffb25; 
        10'b0001000000: data <= 22'h3ffeb4; 
        10'b0001000001: data <= 22'h3ff871; 
        10'b0001000010: data <= 22'h00073c; 
        10'b0001000011: data <= 22'h0005f8; 
        10'b0001000100: data <= 22'h00127c; 
        10'b0001000101: data <= 22'h000ebd; 
        10'b0001000110: data <= 22'h000d7a; 
        10'b0001000111: data <= 22'h00055a; 
        10'b0001001000: data <= 22'h001226; 
        10'b0001001001: data <= 22'h000631; 
        10'b0001001010: data <= 22'h000541; 
        10'b0001001011: data <= 22'h3ff6cd; 
        10'b0001001100: data <= 22'h3fffbe; 
        10'b0001001101: data <= 22'h3ffbba; 
        10'b0001001110: data <= 22'h3fed38; 
        10'b0001001111: data <= 22'h3ff963; 
        10'b0001010000: data <= 22'h3ffe02; 
        10'b0001010001: data <= 22'h000487; 
        10'b0001010010: data <= 22'h3ffa9b; 
        10'b0001010011: data <= 22'h3ff865; 
        10'b0001010100: data <= 22'h3ff6d8; 
        10'b0001010101: data <= 22'h3ff59a; 
        10'b0001010110: data <= 22'h3ffd07; 
        10'b0001010111: data <= 22'h3ff673; 
        10'b0001011000: data <= 22'h000299; 
        10'b0001011001: data <= 22'h3ff467; 
        10'b0001011010: data <= 22'h3ffbc5; 
        10'b0001011011: data <= 22'h000002; 
        10'b0001011100: data <= 22'h00034d; 
        10'b0001011101: data <= 22'h001d70; 
        10'b0001011110: data <= 22'h002e12; 
        10'b0001011111: data <= 22'h002dc3; 
        10'b0001100000: data <= 22'h002bcb; 
        10'b0001100001: data <= 22'h00406c; 
        10'b0001100010: data <= 22'h002326; 
        10'b0001100011: data <= 22'h000f98; 
        10'b0001100100: data <= 22'h001d9e; 
        10'b0001100101: data <= 22'h000d93; 
        10'b0001100110: data <= 22'h3ff330; 
        10'b0001100111: data <= 22'h3ffcd4; 
        10'b0001101000: data <= 22'h3ff171; 
        10'b0001101001: data <= 22'h3feef2; 
        10'b0001101010: data <= 22'h3feb26; 
        10'b0001101011: data <= 22'h3ff5a7; 
        10'b0001101100: data <= 22'h000187; 
        10'b0001101101: data <= 22'h0004e8; 
        10'b0001101110: data <= 22'h3ff479; 
        10'b0001101111: data <= 22'h3ffdad; 
        10'b0001110000: data <= 22'h3ff5e9; 
        10'b0001110001: data <= 22'h3ff8fe; 
        10'b0001110010: data <= 22'h000387; 
        10'b0001110011: data <= 22'h3ff0f2; 
        10'b0001110100: data <= 22'h3ff2b8; 
        10'b0001110101: data <= 22'h3ffbc5; 
        10'b0001110110: data <= 22'h0006d3; 
        10'b0001110111: data <= 22'h000696; 
        10'b0001111000: data <= 22'h0012f9; 
        10'b0001111001: data <= 22'h003869; 
        10'b0001111010: data <= 22'h0038fc; 
        10'b0001111011: data <= 22'h00479b; 
        10'b0001111100: data <= 22'h003c83; 
        10'b0001111101: data <= 22'h002fff; 
        10'b0001111110: data <= 22'h002b9c; 
        10'b0001111111: data <= 22'h001345; 
        10'b0010000000: data <= 22'h0019c7; 
        10'b0010000001: data <= 22'h0017d5; 
        10'b0010000010: data <= 22'h3ff8db; 
        10'b0010000011: data <= 22'h3ff3f8; 
        10'b0010000100: data <= 22'h3ff6b6; 
        10'b0010000101: data <= 22'h3fe3af; 
        10'b0010000110: data <= 22'h3fddb9; 
        10'b0010000111: data <= 22'h3fdf10; 
        10'b0010001000: data <= 22'h3ffbc7; 
        10'b0010001001: data <= 22'h3ffbc5; 
        10'b0010001010: data <= 22'h3ff238; 
        10'b0010001011: data <= 22'h3ffd66; 
        10'b0010001100: data <= 22'h00012f; 
        10'b0010001101: data <= 22'h3ffb87; 
        10'b0010001110: data <= 22'h3ff523; 
        10'b0010001111: data <= 22'h3ff17b; 
        10'b0010010000: data <= 22'h3ff414; 
        10'b0010010001: data <= 22'h3ff5c0; 
        10'b0010010010: data <= 22'h000650; 
        10'b0010010011: data <= 22'h001b92; 
        10'b0010010100: data <= 22'h002639; 
        10'b0010010101: data <= 22'h004170; 
        10'b0010010110: data <= 22'h00487d; 
        10'b0010010111: data <= 22'h004b9a; 
        10'b0010011000: data <= 22'h004540; 
        10'b0010011001: data <= 22'h004da6; 
        10'b0010011010: data <= 22'h0047df; 
        10'b0010011011: data <= 22'h0042af; 
        10'b0010011100: data <= 22'h004853; 
        10'b0010011101: data <= 22'h003a81; 
        10'b0010011110: data <= 22'h002a45; 
        10'b0010011111: data <= 22'h3fee25; 
        10'b0010100000: data <= 22'h3feec2; 
        10'b0010100001: data <= 22'h3fe3d7; 
        10'b0010100010: data <= 22'h3fe360; 
        10'b0010100011: data <= 22'h3fd39b; 
        10'b0010100100: data <= 22'h3fecd8; 
        10'b0010100101: data <= 22'h3ff51c; 
        10'b0010100110: data <= 22'h0001c4; 
        10'b0010100111: data <= 22'h3ff786; 
        10'b0010101000: data <= 22'h3ffa39; 
        10'b0010101001: data <= 22'h3ff5a7; 
        10'b0010101010: data <= 22'h000256; 
        10'b0010101011: data <= 22'h3ffa70; 
        10'b0010101100: data <= 22'h3ff8b6; 
        10'b0010101101: data <= 22'h00049e; 
        10'b0010101110: data <= 22'h001af5; 
        10'b0010101111: data <= 22'h003430; 
        10'b0010110000: data <= 22'h0027e3; 
        10'b0010110001: data <= 22'h002d49; 
        10'b0010110010: data <= 22'h003d4e; 
        10'b0010110011: data <= 22'h002657; 
        10'b0010110100: data <= 22'h0028be; 
        10'b0010110101: data <= 22'h00349d; 
        10'b0010110110: data <= 22'h002e79; 
        10'b0010110111: data <= 22'h001948; 
        10'b0010111000: data <= 22'h001bfb; 
        10'b0010111001: data <= 22'h00073b; 
        10'b0010111010: data <= 22'h000557; 
        10'b0010111011: data <= 22'h3fef92; 
        10'b0010111100: data <= 22'h3ff514; 
        10'b0010111101: data <= 22'h3fdc2c; 
        10'b0010111110: data <= 22'h3fdc72; 
        10'b0010111111: data <= 22'h3fce65; 
        10'b0011000000: data <= 22'h3fe275; 
        10'b0011000001: data <= 22'h3fef72; 
        10'b0011000010: data <= 22'h00021a; 
        10'b0011000011: data <= 22'h3ffe52; 
        10'b0011000100: data <= 22'h3ff859; 
        10'b0011000101: data <= 22'h000186; 
        10'b0011000110: data <= 22'h0001ab; 
        10'b0011000111: data <= 22'h3ff903; 
        10'b0011001000: data <= 22'h0000b4; 
        10'b0011001001: data <= 22'h000e7e; 
        10'b0011001010: data <= 22'h0022bd; 
        10'b0011001011: data <= 22'h003249; 
        10'b0011001100: data <= 22'h002924; 
        10'b0011001101: data <= 22'h002664; 
        10'b0011001110: data <= 22'h000eac; 
        10'b0011001111: data <= 22'h001155; 
        10'b0011010000: data <= 22'h0002f6; 
        10'b0011010001: data <= 22'h001af3; 
        10'b0011010010: data <= 22'h002134; 
        10'b0011010011: data <= 22'h0006f5; 
        10'b0011010100: data <= 22'h000475; 
        10'b0011010101: data <= 22'h3fd5f0; 
        10'b0011010110: data <= 22'h3ff1be; 
        10'b0011010111: data <= 22'h3ff422; 
        10'b0011011000: data <= 22'h3ff289; 
        10'b0011011001: data <= 22'h3ff03d; 
        10'b0011011010: data <= 22'h3ff440; 
        10'b0011011011: data <= 22'h3fd72f; 
        10'b0011011100: data <= 22'h3fe3bb; 
        10'b0011011101: data <= 22'h3ff75f; 
        10'b0011011110: data <= 22'h3ff51f; 
        10'b0011011111: data <= 22'h3ff2bd; 
        10'b0011100000: data <= 22'h3ffcf7; 
        10'b0011100001: data <= 22'h0001fd; 
        10'b0011100010: data <= 22'h3ffa5a; 
        10'b0011100011: data <= 22'h0001d5; 
        10'b0011100100: data <= 22'h000795; 
        10'b0011100101: data <= 22'h001783; 
        10'b0011100110: data <= 22'h001101; 
        10'b0011100111: data <= 22'h001802; 
        10'b0011101000: data <= 22'h001850; 
        10'b0011101001: data <= 22'h001b0d; 
        10'b0011101010: data <= 22'h001b2d; 
        10'b0011101011: data <= 22'h001f05; 
        10'b0011101100: data <= 22'h001270; 
        10'b0011101101: data <= 22'h001607; 
        10'b0011101110: data <= 22'h003a1e; 
        10'b0011101111: data <= 22'h0020ad; 
        10'b0011110000: data <= 22'h3ffbf9; 
        10'b0011110001: data <= 22'h3ff00c; 
        10'b0011110010: data <= 22'h3fff97; 
        10'b0011110011: data <= 22'h000ce6; 
        10'b0011110100: data <= 22'h00004d; 
        10'b0011110101: data <= 22'h3ff719; 
        10'b0011110110: data <= 22'h3fe850; 
        10'b0011110111: data <= 22'h3fd05e; 
        10'b0011111000: data <= 22'h3fdb74; 
        10'b0011111001: data <= 22'h3ff0c6; 
        10'b0011111010: data <= 22'h3ff8e0; 
        10'b0011111011: data <= 22'h3ff44d; 
        10'b0011111100: data <= 22'h3ff5f3; 
        10'b0011111101: data <= 22'h3ffd8b; 
        10'b0011111110: data <= 22'h3fff75; 
        10'b0011111111: data <= 22'h000618; 
        10'b0100000000: data <= 22'h000bd2; 
        10'b0100000001: data <= 22'h001a57; 
        10'b0100000010: data <= 22'h00093a; 
        10'b0100000011: data <= 22'h0001c8; 
        10'b0100000100: data <= 22'h3ff6e6; 
        10'b0100000101: data <= 22'h000e2c; 
        10'b0100000110: data <= 22'h000b01; 
        10'b0100000111: data <= 22'h000e37; 
        10'b0100001000: data <= 22'h0003b0; 
        10'b0100001001: data <= 22'h3ffe86; 
        10'b0100001010: data <= 22'h0025eb; 
        10'b0100001011: data <= 22'h002901; 
        10'b0100001100: data <= 22'h000e25; 
        10'b0100001101: data <= 22'h000114; 
        10'b0100001110: data <= 22'h3ffc31; 
        10'b0100001111: data <= 22'h3fffa8; 
        10'b0100010000: data <= 22'h3ffe48; 
        10'b0100010001: data <= 22'h3fff16; 
        10'b0100010010: data <= 22'h3ff0f4; 
        10'b0100010011: data <= 22'h3fd77f; 
        10'b0100010100: data <= 22'h3fdd6f; 
        10'b0100010101: data <= 22'h3ff4bf; 
        10'b0100010110: data <= 22'h0001ca; 
        10'b0100010111: data <= 22'h3ff2f1; 
        10'b0100011000: data <= 22'h00028b; 
        10'b0100011001: data <= 22'h3ffd0a; 
        10'b0100011010: data <= 22'h3ffa01; 
        10'b0100011011: data <= 22'h3ff77f; 
        10'b0100011100: data <= 22'h0001cd; 
        10'b0100011101: data <= 22'h3ff992; 
        10'b0100011110: data <= 22'h3ff2d5; 
        10'b0100011111: data <= 22'h3fc013; 
        10'b0100100000: data <= 22'h3fc6ce; 
        10'b0100100001: data <= 22'h3fd4ca; 
        10'b0100100010: data <= 22'h3fbdf3; 
        10'b0100100011: data <= 22'h3fb6bf; 
        10'b0100100100: data <= 22'h3faac6; 
        10'b0100100101: data <= 22'h3fa04b; 
        10'b0100100110: data <= 22'h3fd7d0; 
        10'b0100100111: data <= 22'h00074b; 
        10'b0100101000: data <= 22'h000a58; 
        10'b0100101001: data <= 22'h0001bc; 
        10'b0100101010: data <= 22'h000552; 
        10'b0100101011: data <= 22'h3ff839; 
        10'b0100101100: data <= 22'h3ffa57; 
        10'b0100101101: data <= 22'h3ff833; 
        10'b0100101110: data <= 22'h3febf0; 
        10'b0100101111: data <= 22'h3fd16a; 
        10'b0100110000: data <= 22'h3fe668; 
        10'b0100110001: data <= 22'h3ffeea; 
        10'b0100110010: data <= 22'h3ffed4; 
        10'b0100110011: data <= 22'h3ff53c; 
        10'b0100110100: data <= 22'h3ff2af; 
        10'b0100110101: data <= 22'h000348; 
        10'b0100110110: data <= 22'h3ffea5; 
        10'b0100110111: data <= 22'h3ff3c3; 
        10'b0100111000: data <= 22'h3fe808; 
        10'b0100111001: data <= 22'h3fcb9f; 
        10'b0100111010: data <= 22'h3fa61c; 
        10'b0100111011: data <= 22'h3f8142; 
        10'b0100111100: data <= 22'h3f863f; 
        10'b0100111101: data <= 22'h3f709b; 
        10'b0100111110: data <= 22'h3f7031; 
        10'b0100111111: data <= 22'h3f7cbd; 
        10'b0101000000: data <= 22'h3f74aa; 
        10'b0101000001: data <= 22'h3f5639; 
        10'b0101000010: data <= 22'h3f7d66; 
        10'b0101000011: data <= 22'h3fc188; 
        10'b0101000100: data <= 22'h3fea58; 
        10'b0101000101: data <= 22'h3fed60; 
        10'b0101000110: data <= 22'h3fee19; 
        10'b0101000111: data <= 22'h3ffc6c; 
        10'b0101001000: data <= 22'h3ff53f; 
        10'b0101001001: data <= 22'h3ff4c8; 
        10'b0101001010: data <= 22'h3fe253; 
        10'b0101001011: data <= 22'h3febb2; 
        10'b0101001100: data <= 22'h3ffc51; 
        10'b0101001101: data <= 22'h3ff8fc; 
        10'b0101001110: data <= 22'h3ff4e4; 
        10'b0101001111: data <= 22'h3ffcea; 
        10'b0101010000: data <= 22'h3ffb63; 
        10'b0101010001: data <= 22'h3ffc31; 
        10'b0101010010: data <= 22'h000155; 
        10'b0101010011: data <= 22'h3ffa69; 
        10'b0101010100: data <= 22'h3fe632; 
        10'b0101010101: data <= 22'h3fb201; 
        10'b0101010110: data <= 22'h3f6845; 
        10'b0101010111: data <= 22'h3f4659; 
        10'b0101011000: data <= 22'h3f52d7; 
        10'b0101011001: data <= 22'h3f5be4; 
        10'b0101011010: data <= 22'h3f6a09; 
        10'b0101011011: data <= 22'h3f73ac; 
        10'b0101011100: data <= 22'h3f7412; 
        10'b0101011101: data <= 22'h3f6e68; 
        10'b0101011110: data <= 22'h3f8869; 
        10'b0101011111: data <= 22'h3fb03f; 
        10'b0101100000: data <= 22'h3fc945; 
        10'b0101100001: data <= 22'h3fced8; 
        10'b0101100010: data <= 22'h3fe73a; 
        10'b0101100011: data <= 22'h00001b; 
        10'b0101100100: data <= 22'h3fff85; 
        10'b0101100101: data <= 22'h3ff21b; 
        10'b0101100110: data <= 22'h3fe06c; 
        10'b0101100111: data <= 22'h3fcff9; 
        10'b0101101000: data <= 22'h3ffa27; 
        10'b0101101001: data <= 22'h3ff80b; 
        10'b0101101010: data <= 22'h000391; 
        10'b0101101011: data <= 22'h3ffc30; 
        10'b0101101100: data <= 22'h3ff659; 
        10'b0101101101: data <= 22'h3ff9ac; 
        10'b0101101110: data <= 22'h000354; 
        10'b0101101111: data <= 22'h3ff604; 
        10'b0101110000: data <= 22'h3fd63b; 
        10'b0101110001: data <= 22'h3f9da6; 
        10'b0101110010: data <= 22'h3f63eb; 
        10'b0101110011: data <= 22'h3f70ba; 
        10'b0101110100: data <= 22'h3f7a47; 
        10'b0101110101: data <= 22'h3fa416; 
        10'b0101110110: data <= 22'h3fbedd; 
        10'b0101110111: data <= 22'h3fe180; 
        10'b0101111000: data <= 22'h3fcfc1; 
        10'b0101111001: data <= 22'h3fea0e; 
        10'b0101111010: data <= 22'h3fc8e6; 
        10'b0101111011: data <= 22'h3fc7c7; 
        10'b0101111100: data <= 22'h3fbd50; 
        10'b0101111101: data <= 22'h3fcfdc; 
        10'b0101111110: data <= 22'h3fe57b; 
        10'b0101111111: data <= 22'h3ffaeb; 
        10'b0110000000: data <= 22'h3ff838; 
        10'b0110000001: data <= 22'h3feee9; 
        10'b0110000010: data <= 22'h3fd84b; 
        10'b0110000011: data <= 22'h3fdbdb; 
        10'b0110000100: data <= 22'h3fedb7; 
        10'b0110000101: data <= 22'h000496; 
        10'b0110000110: data <= 22'h3ff9e5; 
        10'b0110000111: data <= 22'h3fff98; 
        10'b0110001000: data <= 22'h000215; 
        10'b0110001001: data <= 22'h3ffcae; 
        10'b0110001010: data <= 22'h000059; 
        10'b0110001011: data <= 22'h3ff798; 
        10'b0110001100: data <= 22'h3ff001; 
        10'b0110001101: data <= 22'h3fbd91; 
        10'b0110001110: data <= 22'h3fabf5; 
        10'b0110001111: data <= 22'h3fbb7c; 
        10'b0110010000: data <= 22'h3fe485; 
        10'b0110010001: data <= 22'h3ffb42; 
        10'b0110010010: data <= 22'h001122; 
        10'b0110010011: data <= 22'h0016ac; 
        10'b0110010100: data <= 22'h001ae7; 
        10'b0110010101: data <= 22'h0029dc; 
        10'b0110010110: data <= 22'h0002db; 
        10'b0110010111: data <= 22'h3fe532; 
        10'b0110011000: data <= 22'h3fec16; 
        10'b0110011001: data <= 22'h3fdd7e; 
        10'b0110011010: data <= 22'h3ffa32; 
        10'b0110011011: data <= 22'h3fe9cf; 
        10'b0110011100: data <= 22'h3ff8fc; 
        10'b0110011101: data <= 22'h3fe66f; 
        10'b0110011110: data <= 22'h3fd20b; 
        10'b0110011111: data <= 22'h3fde96; 
        10'b0110100000: data <= 22'h3ff977; 
        10'b0110100001: data <= 22'h001044; 
        10'b0110100010: data <= 22'h001276; 
        10'b0110100011: data <= 22'h3ff5be; 
        10'b0110100100: data <= 22'h3ff8d0; 
        10'b0110100101: data <= 22'h3ffa52; 
        10'b0110100110: data <= 22'h3ff897; 
        10'b0110100111: data <= 22'h000f2f; 
        10'b0110101000: data <= 22'h00075a; 
        10'b0110101001: data <= 22'h000351; 
        10'b0110101010: data <= 22'h0011f8; 
        10'b0110101011: data <= 22'h00150c; 
        10'b0110101100: data <= 22'h00271d; 
        10'b0110101101: data <= 22'h001ba3; 
        10'b0110101110: data <= 22'h002125; 
        10'b0110101111: data <= 22'h00137b; 
        10'b0110110000: data <= 22'h00113f; 
        10'b0110110001: data <= 22'h002872; 
        10'b0110110010: data <= 22'h000302; 
        10'b0110110011: data <= 22'h000fdf; 
        10'b0110110100: data <= 22'h000244; 
        10'b0110110101: data <= 22'h3fdfec; 
        10'b0110110110: data <= 22'h3fe17b; 
        10'b0110110111: data <= 22'h3fed47; 
        10'b0110111000: data <= 22'h3ff25a; 
        10'b0110111001: data <= 22'h3feb5c; 
        10'b0110111010: data <= 22'h3fd65c; 
        10'b0110111011: data <= 22'h3fea93; 
        10'b0110111100: data <= 22'h000ccd; 
        10'b0110111101: data <= 22'h0015d2; 
        10'b0110111110: data <= 22'h000bc9; 
        10'b0110111111: data <= 22'h3ff455; 
        10'b0111000000: data <= 22'h3ff717; 
        10'b0111000001: data <= 22'h3ff229; 
        10'b0111000010: data <= 22'h3ff050; 
        10'b0111000011: data <= 22'h001027; 
        10'b0111000100: data <= 22'h0021e1; 
        10'b0111000101: data <= 22'h00374f; 
        10'b0111000110: data <= 22'h003857; 
        10'b0111000111: data <= 22'h002187; 
        10'b0111001000: data <= 22'h000de7; 
        10'b0111001001: data <= 22'h001cec; 
        10'b0111001010: data <= 22'h001adc; 
        10'b0111001011: data <= 22'h001888; 
        10'b0111001100: data <= 22'h00328a; 
        10'b0111001101: data <= 22'h002c82; 
        10'b0111001110: data <= 22'h000957; 
        10'b0111001111: data <= 22'h3ffaae; 
        10'b0111010000: data <= 22'h3fffcc; 
        10'b0111010001: data <= 22'h3feb2b; 
        10'b0111010010: data <= 22'h3fedc8; 
        10'b0111010011: data <= 22'h3fe00b; 
        10'b0111010100: data <= 22'h3ff4a4; 
        10'b0111010101: data <= 22'h0001ba; 
        10'b0111010110: data <= 22'h000707; 
        10'b0111010111: data <= 22'h000ed9; 
        10'b0111011000: data <= 22'h002f32; 
        10'b0111011001: data <= 22'h003a74; 
        10'b0111011010: data <= 22'h0009c9; 
        10'b0111011011: data <= 22'h3ff6db; 
        10'b0111011100: data <= 22'h3ff872; 
        10'b0111011101: data <= 22'h0002ab; 
        10'b0111011110: data <= 22'h3ffa1d; 
        10'b0111011111: data <= 22'h001395; 
        10'b0111100000: data <= 22'h0039db; 
        10'b0111100001: data <= 22'h00509b; 
        10'b0111100010: data <= 22'h0049aa; 
        10'b0111100011: data <= 22'h003279; 
        10'b0111100100: data <= 22'h002320; 
        10'b0111100101: data <= 22'h002a97; 
        10'b0111100110: data <= 22'h00417e; 
        10'b0111100111: data <= 22'h0035ae; 
        10'b0111101000: data <= 22'h003d8f; 
        10'b0111101001: data <= 22'h001cce; 
        10'b0111101010: data <= 22'h000ed6; 
        10'b0111101011: data <= 22'h001403; 
        10'b0111101100: data <= 22'h001436; 
        10'b0111101101: data <= 22'h3ffce0; 
        10'b0111101110: data <= 22'h000d1c; 
        10'b0111101111: data <= 22'h3ff7a3; 
        10'b0111110000: data <= 22'h00182e; 
        10'b0111110001: data <= 22'h0019cc; 
        10'b0111110010: data <= 22'h00132b; 
        10'b0111110011: data <= 22'h001a92; 
        10'b0111110100: data <= 22'h004b9e; 
        10'b0111110101: data <= 22'h004196; 
        10'b0111110110: data <= 22'h000ef8; 
        10'b0111110111: data <= 22'h0001fd; 
        10'b0111111000: data <= 22'h3ffe4c; 
        10'b0111111001: data <= 22'h3fff13; 
        10'b0111111010: data <= 22'h3fec15; 
        10'b0111111011: data <= 22'h000545; 
        10'b0111111100: data <= 22'h003eb4; 
        10'b0111111101: data <= 22'h0069f4; 
        10'b0111111110: data <= 22'h0063a9; 
        10'b0111111111: data <= 22'h0047bd; 
        10'b1000000000: data <= 22'h002fdb; 
        10'b1000000001: data <= 22'h003532; 
        10'b1000000010: data <= 22'h00514d; 
        10'b1000000011: data <= 22'h004974; 
        10'b1000000100: data <= 22'h007502; 
        10'b1000000101: data <= 22'h005567; 
        10'b1000000110: data <= 22'h004a95; 
        10'b1000000111: data <= 22'h00244b; 
        10'b1000001000: data <= 22'h0018fa; 
        10'b1000001001: data <= 22'h002de2; 
        10'b1000001010: data <= 22'h001d9a; 
        10'b1000001011: data <= 22'h001428; 
        10'b1000001100: data <= 22'h003621; 
        10'b1000001101: data <= 22'h0037eb; 
        10'b1000001110: data <= 22'h003cf2; 
        10'b1000001111: data <= 22'h005087; 
        10'b1000010000: data <= 22'h0063ee; 
        10'b1000010001: data <= 22'h0039a0; 
        10'b1000010010: data <= 22'h3ffa79; 
        10'b1000010011: data <= 22'h3ff41f; 
        10'b1000010100: data <= 22'h3ff5e2; 
        10'b1000010101: data <= 22'h3ff68d; 
        10'b1000010110: data <= 22'h3ff218; 
        10'b1000010111: data <= 22'h3fffc4; 
        10'b1000011000: data <= 22'h002274; 
        10'b1000011001: data <= 22'h00405d; 
        10'b1000011010: data <= 22'h005148; 
        10'b1000011011: data <= 22'h00467a; 
        10'b1000011100: data <= 22'h00410f; 
        10'b1000011101: data <= 22'h0044de; 
        10'b1000011110: data <= 22'h0041ea; 
        10'b1000011111: data <= 22'h004600; 
        10'b1000100000: data <= 22'h004e58; 
        10'b1000100001: data <= 22'h003c43; 
        10'b1000100010: data <= 22'h002707; 
        10'b1000100011: data <= 22'h001281; 
        10'b1000100100: data <= 22'h001cbf; 
        10'b1000100101: data <= 22'h0031ec; 
        10'b1000100110: data <= 22'h00181e; 
        10'b1000100111: data <= 22'h001790; 
        10'b1000101000: data <= 22'h002837; 
        10'b1000101001: data <= 22'h00322f; 
        10'b1000101010: data <= 22'h004188; 
        10'b1000101011: data <= 22'h00464a; 
        10'b1000101100: data <= 22'h003c94; 
        10'b1000101101: data <= 22'h001fbb; 
        10'b1000101110: data <= 22'h0002af; 
        10'b1000101111: data <= 22'h0000bb; 
        10'b1000110000: data <= 22'h3ff372; 
        10'b1000110001: data <= 22'h3fff05; 
        10'b1000110010: data <= 22'h3ffca7; 
        10'b1000110011: data <= 22'h3feebf; 
        10'b1000110100: data <= 22'h001e93; 
        10'b1000110101: data <= 22'h0025c4; 
        10'b1000110110: data <= 22'h003aa0; 
        10'b1000110111: data <= 22'h005187; 
        10'b1000111000: data <= 22'h004d71; 
        10'b1000111001: data <= 22'h00334f; 
        10'b1000111010: data <= 22'h003155; 
        10'b1000111011: data <= 22'h005293; 
        10'b1000111100: data <= 22'h002de9; 
        10'b1000111101: data <= 22'h000f33; 
        10'b1000111110: data <= 22'h000a2f; 
        10'b1000111111: data <= 22'h000c82; 
        10'b1001000000: data <= 22'h00102f; 
        10'b1001000001: data <= 22'h0000bb; 
        10'b1001000010: data <= 22'h0023b3; 
        10'b1001000011: data <= 22'h0037c0; 
        10'b1001000100: data <= 22'h0025d4; 
        10'b1001000101: data <= 22'h0035ce; 
        10'b1001000110: data <= 22'h004aee; 
        10'b1001000111: data <= 22'h004101; 
        10'b1001001000: data <= 22'h002eca; 
        10'b1001001001: data <= 22'h00162f; 
        10'b1001001010: data <= 22'h3fffb8; 
        10'b1001001011: data <= 22'h3ffdf0; 
        10'b1001001100: data <= 22'h3ffb15; 
        10'b1001001101: data <= 22'h3ff405; 
        10'b1001001110: data <= 22'h3ffdda; 
        10'b1001001111: data <= 22'h3ff919; 
        10'b1001010000: data <= 22'h000664; 
        10'b1001010001: data <= 22'h00103d; 
        10'b1001010010: data <= 22'h0028aa; 
        10'b1001010011: data <= 22'h002db0; 
        10'b1001010100: data <= 22'h002846; 
        10'b1001010101: data <= 22'h003244; 
        10'b1001010110: data <= 22'h002c77; 
        10'b1001010111: data <= 22'h002ba9; 
        10'b1001011000: data <= 22'h001124; 
        10'b1001011001: data <= 22'h000829; 
        10'b1001011010: data <= 22'h3ffb92; 
        10'b1001011011: data <= 22'h0001e4; 
        10'b1001011100: data <= 22'h0015b8; 
        10'b1001011101: data <= 22'h0017cc; 
        10'b1001011110: data <= 22'h003421; 
        10'b1001011111: data <= 22'h0036d7; 
        10'b1001100000: data <= 22'h00180f; 
        10'b1001100001: data <= 22'h0035c7; 
        10'b1001100010: data <= 22'h00426e; 
        10'b1001100011: data <= 22'h004bac; 
        10'b1001100100: data <= 22'h00254a; 
        10'b1001100101: data <= 22'h000eca; 
        10'b1001100110: data <= 22'h00036a; 
        10'b1001100111: data <= 22'h3ffe56; 
        10'b1001101000: data <= 22'h3ff35b; 
        10'b1001101001: data <= 22'h3ffc9d; 
        10'b1001101010: data <= 22'h3ff51a; 
        10'b1001101011: data <= 22'h000396; 
        10'b1001101100: data <= 22'h000cca; 
        10'b1001101101: data <= 22'h00049e; 
        10'b1001101110: data <= 22'h001bae; 
        10'b1001101111: data <= 22'h001847; 
        10'b1001110000: data <= 22'h0016a3; 
        10'b1001110001: data <= 22'h001fcb; 
        10'b1001110010: data <= 22'h001f91; 
        10'b1001110011: data <= 22'h00256d; 
        10'b1001110100: data <= 22'h00040d; 
        10'b1001110101: data <= 22'h3fe26f; 
        10'b1001110110: data <= 22'h3fdac8; 
        10'b1001110111: data <= 22'h3feaed; 
        10'b1001111000: data <= 22'h3fec26; 
        10'b1001111001: data <= 22'h000f6c; 
        10'b1001111010: data <= 22'h003076; 
        10'b1001111011: data <= 22'h003dde; 
        10'b1001111100: data <= 22'h003841; 
        10'b1001111101: data <= 22'h0035d2; 
        10'b1001111110: data <= 22'h002ebb; 
        10'b1001111111: data <= 22'h00338a; 
        10'b1010000000: data <= 22'h001327; 
        10'b1010000001: data <= 22'h3ffde1; 
        10'b1010000010: data <= 22'h3ffcbb; 
        10'b1010000011: data <= 22'h3ff707; 
        10'b1010000100: data <= 22'h3ffcef; 
        10'b1010000101: data <= 22'h3ffd50; 
        10'b1010000110: data <= 22'h3ffa6b; 
        10'b1010000111: data <= 22'h3ff981; 
        10'b1010001000: data <= 22'h3ff8bf; 
        10'b1010001001: data <= 22'h3ff19a; 
        10'b1010001010: data <= 22'h3fee54; 
        10'b1010001011: data <= 22'h3ff0a7; 
        10'b1010001100: data <= 22'h3fe6d4; 
        10'b1010001101: data <= 22'h3ff13c; 
        10'b1010001110: data <= 22'h3ff621; 
        10'b1010001111: data <= 22'h000cb9; 
        10'b1010010000: data <= 22'h00012b; 
        10'b1010010001: data <= 22'h3fec31; 
        10'b1010010010: data <= 22'h3fe531; 
        10'b1010010011: data <= 22'h3fdd00; 
        10'b1010010100: data <= 22'h3fda01; 
        10'b1010010101: data <= 22'h3fec33; 
        10'b1010010110: data <= 22'h0007c2; 
        10'b1010010111: data <= 22'h00306e; 
        10'b1010011000: data <= 22'h002a64; 
        10'b1010011001: data <= 22'h0033e9; 
        10'b1010011010: data <= 22'h002541; 
        10'b1010011011: data <= 22'h000e3c; 
        10'b1010011100: data <= 22'h00089c; 
        10'b1010011101: data <= 22'h00057d; 
        10'b1010011110: data <= 22'h3ffec9; 
        10'b1010011111: data <= 22'h3ff956; 
        10'b1010100000: data <= 22'h3ffb3f; 
        10'b1010100001: data <= 22'h3ff62e; 
        10'b1010100010: data <= 22'h3fff85; 
        10'b1010100011: data <= 22'h3ffe53; 
        10'b1010100100: data <= 22'h3ff59a; 
        10'b1010100101: data <= 22'h3fe4e5; 
        10'b1010100110: data <= 22'h3fcba0; 
        10'b1010100111: data <= 22'h3fd8d8; 
        10'b1010101000: data <= 22'h3fd7b2; 
        10'b1010101001: data <= 22'h3fd4fd; 
        10'b1010101010: data <= 22'h3fd552; 
        10'b1010101011: data <= 22'h3fdf4f; 
        10'b1010101100: data <= 22'h3fdf0e; 
        10'b1010101101: data <= 22'h3fee1c; 
        10'b1010101110: data <= 22'h3fe8a6; 
        10'b1010101111: data <= 22'h3fdeb8; 
        10'b1010110000: data <= 22'h3fe067; 
        10'b1010110001: data <= 22'h3fe73a; 
        10'b1010110010: data <= 22'h3fe1b7; 
        10'b1010110011: data <= 22'h3fefa5; 
        10'b1010110100: data <= 22'h3ff188; 
        10'b1010110101: data <= 22'h3ff19f; 
        10'b1010110110: data <= 22'h3ff796; 
        10'b1010110111: data <= 22'h3ff958; 
        10'b1010111000: data <= 22'h3fff00; 
        10'b1010111001: data <= 22'h000567; 
        10'b1010111010: data <= 22'h3ff4b1; 
        10'b1010111011: data <= 22'h3ff503; 
        10'b1010111100: data <= 22'h3fff87; 
        10'b1010111101: data <= 22'h3ff1d9; 
        10'b1010111110: data <= 22'h3ff8cc; 
        10'b1010111111: data <= 22'h3ff758; 
        10'b1011000000: data <= 22'h3ff4d4; 
        10'b1011000001: data <= 22'h3fece7; 
        10'b1011000010: data <= 22'h3fe693; 
        10'b1011000011: data <= 22'h3fd94c; 
        10'b1011000100: data <= 22'h3fd509; 
        10'b1011000101: data <= 22'h3fd829; 
        10'b1011000110: data <= 22'h3fdbed; 
        10'b1011000111: data <= 22'h3fd20f; 
        10'b1011001000: data <= 22'h3fe13a; 
        10'b1011001001: data <= 22'h3fe324; 
        10'b1011001010: data <= 22'h3fd9b7; 
        10'b1011001011: data <= 22'h3fe074; 
        10'b1011001100: data <= 22'h3fe896; 
        10'b1011001101: data <= 22'h3fea0b; 
        10'b1011001110: data <= 22'h3ff79c; 
        10'b1011001111: data <= 22'h3febed; 
        10'b1011010000: data <= 22'h3ff8ca; 
        10'b1011010001: data <= 22'h3ff83f; 
        10'b1011010010: data <= 22'h3fffab; 
        10'b1011010011: data <= 22'h3ff52c; 
        10'b1011010100: data <= 22'h3ffbf0; 
        10'b1011010101: data <= 22'h3ff56a; 
        10'b1011010110: data <= 22'h3ff23f; 
        10'b1011010111: data <= 22'h3ff59a; 
        10'b1011011000: data <= 22'h3ff2bf; 
        10'b1011011001: data <= 22'h3ff79f; 
        10'b1011011010: data <= 22'h3ff9ea; 
        10'b1011011011: data <= 22'h0000a1; 
        10'b1011011100: data <= 22'h3ffdd5; 
        10'b1011011101: data <= 22'h3ff95c; 
        10'b1011011110: data <= 22'h3ffd56; 
        10'b1011011111: data <= 22'h3fff87; 
        10'b1011100000: data <= 22'h3ff914; 
        10'b1011100001: data <= 22'h0000cc; 
        10'b1011100010: data <= 22'h3fffc1; 
        10'b1011100011: data <= 22'h000074; 
        10'b1011100100: data <= 22'h000147; 
        10'b1011100101: data <= 22'h3ffbf0; 
        10'b1011100110: data <= 22'h3ff6d2; 
        10'b1011100111: data <= 22'h3ff0f9; 
        10'b1011101000: data <= 22'h3ff81a; 
        10'b1011101001: data <= 22'h3ffbd0; 
        10'b1011101010: data <= 22'h3ffaff; 
        10'b1011101011: data <= 22'h3ff54b; 
        10'b1011101100: data <= 22'h000163; 
        10'b1011101101: data <= 22'h3fffbd; 
        10'b1011101110: data <= 22'h3ff567; 
        10'b1011101111: data <= 22'h3ff7a4; 
        10'b1011110000: data <= 22'h3ff28d; 
        10'b1011110001: data <= 22'h00009b; 
        10'b1011110010: data <= 22'h00006e; 
        10'b1011110011: data <= 22'h3fff48; 
        10'b1011110100: data <= 22'h3ffedf; 
        10'b1011110101: data <= 22'h3ff63a; 
        10'b1011110110: data <= 22'h3ff3d2; 
        10'b1011110111: data <= 22'h3ffb2b; 
        10'b1011111000: data <= 22'h3ff260; 
        10'b1011111001: data <= 22'h0002d2; 
        10'b1011111010: data <= 22'h00028c; 
        10'b1011111011: data <= 22'h3ff813; 
        10'b1011111100: data <= 22'h3fff2a; 
        10'b1011111101: data <= 22'h3ff546; 
        10'b1011111110: data <= 22'h0001de; 
        10'b1011111111: data <= 22'h3ff208; 
        10'b1100000000: data <= 22'h3fff43; 
        10'b1100000001: data <= 22'h3ff93e; 
        10'b1100000010: data <= 22'h3ffcdc; 
        10'b1100000011: data <= 22'h3ff420; 
        10'b1100000100: data <= 22'h3ffb1a; 
        10'b1100000101: data <= 22'h3ff8b5; 
        10'b1100000110: data <= 22'h3ffbd3; 
        10'b1100000111: data <= 22'h3ffacb; 
        10'b1100001000: data <= 22'h3ffe73; 
        10'b1100001001: data <= 22'h3ff17d; 
        10'b1100001010: data <= 22'h3ff9c2; 
        10'b1100001011: data <= 22'h00007b; 
        10'b1100001100: data <= 22'h3ff17b; 
        10'b1100001101: data <= 22'h3ffa81; 
        10'b1100001110: data <= 22'h3ffdec; 
        10'b1100001111: data <= 22'h3ff83a; 
      endcase 
    end 
  end 
endgenerate 
assign dout = data; 
endmodule
