`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// WEIGHT MEMORY
// This code create bram for 1 of 10 weights strings
// and send element with input address from the string to out.
//////////////////////////////////////////////////////////////////////////////////

module ROM_weights_9 #( 
    parameter int BITS = 24 // bit depth
)(
    input logic clk, // clock
    input logic [9:0] address, // address of current element from string
    output [BITS-1:0] dout // current element from string
);

(* rom_style = "block" *) reg [BITS-1:0] data;

always @(posedge clk)
begin
case(address)
10'b0000000000: data <= 24'h000091; 
10'b0000000001: data <= 24'h00007f; 
10'b0000000010: data <= 24'hffffd9; 
10'b0000000011: data <= 24'h000059; 
10'b0000000100: data <= 24'h000052; 
10'b0000000101: data <= 24'h000085; 
10'b0000000110: data <= 24'hffffce; 
10'b0000000111: data <= 24'h000019; 
10'b0000001000: data <= 24'h000099; 
10'b0000001001: data <= 24'hffffc2; 
10'b0000001010: data <= 24'hffffee; 
10'b0000001011: data <= 24'h000043; 
10'b0000001100: data <= 24'h0000c1; 
10'b0000001101: data <= 24'h00007e; 
10'b0000001110: data <= 24'hffffb1; 
10'b0000001111: data <= 24'hffffdc; 
10'b0000010000: data <= 24'hffffd8; 
10'b0000010001: data <= 24'h00004c; 
10'b0000010010: data <= 24'h00008b; 
10'b0000010011: data <= 24'h00000a; 
10'b0000010100: data <= 24'h00000e; 
10'b0000010101: data <= 24'hfffff6; 
10'b0000010110: data <= 24'hffffc2; 
10'b0000010111: data <= 24'h000016; 
10'b0000011000: data <= 24'h00009c; 
10'b0000011001: data <= 24'h00002f; 
10'b0000011010: data <= 24'hffffb9; 
10'b0000011011: data <= 24'h00004e; 
10'b0000011100: data <= 24'h000082; 
10'b0000011101: data <= 24'h00006c; 
10'b0000011110: data <= 24'h000034; 
10'b0000011111: data <= 24'hffffe2; 
10'b0000100000: data <= 24'hffffb5; 
10'b0000100001: data <= 24'hffffc3; 
10'b0000100010: data <= 24'hfffff4; 
10'b0000100011: data <= 24'h0000c2; 
10'b0000100100: data <= 24'hffffb7; 
10'b0000100101: data <= 24'h00009d; 
10'b0000100110: data <= 24'h00003d; 
10'b0000100111: data <= 24'h000061; 
10'b0000101000: data <= 24'h00004c; 
10'b0000101001: data <= 24'h00006e; 
10'b0000101010: data <= 24'h000003; 
10'b0000101011: data <= 24'hffffab; 
10'b0000101100: data <= 24'hffffd4; 
10'b0000101101: data <= 24'h000078; 
10'b0000101110: data <= 24'hfffffb; 
10'b0000101111: data <= 24'h000022; 
10'b0000110000: data <= 24'h000098; 
10'b0000110001: data <= 24'hfffff5; 
10'b0000110010: data <= 24'h00001b; 
10'b0000110011: data <= 24'h00000e; 
10'b0000110100: data <= 24'h000054; 
10'b0000110101: data <= 24'h0000a3; 
10'b0000110110: data <= 24'hfffffe; 
10'b0000110111: data <= 24'h000023; 
10'b0000111000: data <= 24'h0000ab; 
10'b0000111001: data <= 24'h0000b0; 
10'b0000111010: data <= 24'h00000d; 
10'b0000111011: data <= 24'h000078; 
10'b0000111100: data <= 24'h000091; 
10'b0000111101: data <= 24'hfffff9; 
10'b0000111110: data <= 24'hffffef; 
10'b0000111111: data <= 24'h000034; 
10'b0001000000: data <= 24'h000092; 
10'b0001000001: data <= 24'hffffeb; 
10'b0001000010: data <= 24'hffffd4; 
10'b0001000011: data <= 24'h00006f; 
10'b0001000100: data <= 24'h000042; 
10'b0001000101: data <= 24'h00008b; 
10'b0001000110: data <= 24'hffffae; 
10'b0001000111: data <= 24'h000093; 
10'b0001001000: data <= 24'hffffcb; 
10'b0001001001: data <= 24'hffffc8; 
10'b0001001010: data <= 24'h00000d; 
10'b0001001011: data <= 24'hffffba; 
10'b0001001100: data <= 24'h0000a9; 
10'b0001001101: data <= 24'hffffd4; 
10'b0001001110: data <= 24'hffffc3; 
10'b0001001111: data <= 24'h0000a8; 
10'b0001010000: data <= 24'h00001e; 
10'b0001010001: data <= 24'h00001d; 
10'b0001010010: data <= 24'h000025; 
10'b0001010011: data <= 24'h00004b; 
10'b0001010100: data <= 24'h0000d1; 
10'b0001010101: data <= 24'h000007; 
10'b0001010110: data <= 24'hffffed; 
10'b0001010111: data <= 24'h00003e; 
10'b0001011000: data <= 24'h000042; 
10'b0001011001: data <= 24'hffffbb; 
10'b0001011010: data <= 24'h0000ab; 
10'b0001011011: data <= 24'h00005e; 
10'b0001011100: data <= 24'hffffde; 
10'b0001011101: data <= 24'h0000ad; 
10'b0001011110: data <= 24'h000036; 
10'b0001011111: data <= 24'h000088; 
10'b0001100000: data <= 24'hfffff2; 
10'b0001100001: data <= 24'hffff64; 
10'b0001100010: data <= 24'hfffff2; 
10'b0001100011: data <= 24'hffff13; 
10'b0001100100: data <= 24'hffffe3; 
10'b0001100101: data <= 24'hffff85; 
10'b0001100110: data <= 24'h000029; 
10'b0001100111: data <= 24'h000019; 
10'b0001101000: data <= 24'h000035; 
10'b0001101001: data <= 24'hfffff3; 
10'b0001101010: data <= 24'h000088; 
10'b0001101011: data <= 24'hffffef; 
10'b0001101100: data <= 24'hffffec; 
10'b0001101101: data <= 24'h0000bb; 
10'b0001101110: data <= 24'h000046; 
10'b0001101111: data <= 24'h000077; 
10'b0001110000: data <= 24'h000017; 
10'b0001110001: data <= 24'h000027; 
10'b0001110010: data <= 24'h000009; 
10'b0001110011: data <= 24'hffffd8; 
10'b0001110100: data <= 24'hffffbd; 
10'b0001110101: data <= 24'h000079; 
10'b0001110110: data <= 24'h000053; 
10'b0001110111: data <= 24'hfffff1; 
10'b0001111000: data <= 24'hffff96; 
10'b0001111001: data <= 24'h000028; 
10'b0001111010: data <= 24'hffff51; 
10'b0001111011: data <= 24'hffff09; 
10'b0001111100: data <= 24'hfffea5; 
10'b0001111101: data <= 24'hfffd8a; 
10'b0001111110: data <= 24'hfffcdf; 
10'b0001111111: data <= 24'hfffbd1; 
10'b0010000000: data <= 24'hfffce8; 
10'b0010000001: data <= 24'hfffce6; 
10'b0010000010: data <= 24'hfffdb1; 
10'b0010000011: data <= 24'hfffefc; 
10'b0010000100: data <= 24'hffff86; 
10'b0010000101: data <= 24'hffffa8; 
10'b0010000110: data <= 24'h00001d; 
10'b0010000111: data <= 24'h000095; 
10'b0010001000: data <= 24'h000075; 
10'b0010001001: data <= 24'h00006c; 
10'b0010001010: data <= 24'h000001; 
10'b0010001011: data <= 24'h000005; 
10'b0010001100: data <= 24'h000091; 
10'b0010001101: data <= 24'h000067; 
10'b0010001110: data <= 24'h000078; 
10'b0010001111: data <= 24'h00004c; 
10'b0010010000: data <= 24'h00005c; 
10'b0010010001: data <= 24'hffff8e; 
10'b0010010010: data <= 24'hffff9a; 
10'b0010010011: data <= 24'hffff8f; 
10'b0010010100: data <= 24'hfffe94; 
10'b0010010101: data <= 24'hfffe9c; 
10'b0010010110: data <= 24'hfffe7f; 
10'b0010010111: data <= 24'hfffe05; 
10'b0010011000: data <= 24'hfffd85; 
10'b0010011001: data <= 24'hfffd11; 
10'b0010011010: data <= 24'hfffb85; 
10'b0010011011: data <= 24'hfffb2a; 
10'b0010011100: data <= 24'hfff9e3; 
10'b0010011101: data <= 24'hfffbf8; 
10'b0010011110: data <= 24'hfffd76; 
10'b0010011111: data <= 24'hfffec5; 
10'b0010100000: data <= 24'hfffeb4; 
10'b0010100001: data <= 24'hfffe4f; 
10'b0010100010: data <= 24'hfffe6d; 
10'b0010100011: data <= 24'hfffee1; 
10'b0010100100: data <= 24'hffff8e; 
10'b0010100101: data <= 24'hffffcb; 
10'b0010100110: data <= 24'h000012; 
10'b0010100111: data <= 24'h000065; 
10'b0010101000: data <= 24'h000082; 
10'b0010101001: data <= 24'h000086; 
10'b0010101010: data <= 24'hffffac; 
10'b0010101011: data <= 24'h000087; 
10'b0010101100: data <= 24'h000056; 
10'b0010101101: data <= 24'hfffe7d; 
10'b0010101110: data <= 24'hfffe29; 
10'b0010101111: data <= 24'hfffdd5; 
10'b0010110000: data <= 24'hfffd8f; 
10'b0010110001: data <= 24'hfffd01; 
10'b0010110010: data <= 24'hfffdcd; 
10'b0010110011: data <= 24'hffff4c; 
10'b0010110100: data <= 24'h00002d; 
10'b0010110101: data <= 24'h0002b5; 
10'b0010110110: data <= 24'h000409; 
10'b0010110111: data <= 24'h000336; 
10'b0010111000: data <= 24'h000240; 
10'b0010111001: data <= 24'h0001de; 
10'b0010111010: data <= 24'h00025f; 
10'b0010111011: data <= 24'hffff9a; 
10'b0010111100: data <= 24'hffff6e; 
10'b0010111101: data <= 24'hfffe32; 
10'b0010111110: data <= 24'hfffcc5; 
10'b0010111111: data <= 24'hfffcfe; 
10'b0011000000: data <= 24'hfffe47; 
10'b0011000001: data <= 24'hffff29; 
10'b0011000010: data <= 24'hffffdf; 
10'b0011000011: data <= 24'h000046; 
10'b0011000100: data <= 24'h0000c7; 
10'b0011000101: data <= 24'hfffff9; 
10'b0011000110: data <= 24'hffffbf; 
10'b0011000111: data <= 24'hffffb8; 
10'b0011001000: data <= 24'hfffe46; 
10'b0011001001: data <= 24'hfffd60; 
10'b0011001010: data <= 24'hfffce8; 
10'b0011001011: data <= 24'hfffc52; 
10'b0011001100: data <= 24'hfffc85; 
10'b0011001101: data <= 24'hfffec6; 
10'b0011001110: data <= 24'hffffe6; 
10'b0011001111: data <= 24'h0000f4; 
10'b0011010000: data <= 24'h0003ab; 
10'b0011010001: data <= 24'h000460; 
10'b0011010010: data <= 24'h000600; 
10'b0011010011: data <= 24'h000608; 
10'b0011010100: data <= 24'h000646; 
10'b0011010101: data <= 24'h0002d8; 
10'b0011010110: data <= 24'h000224; 
10'b0011010111: data <= 24'h00003b; 
10'b0011011000: data <= 24'h00008e; 
10'b0011011001: data <= 24'h0000a1; 
10'b0011011010: data <= 24'hfffdd7; 
10'b0011011011: data <= 24'hfffc21; 
10'b0011011100: data <= 24'hfffdb8; 
10'b0011011101: data <= 24'hffff6e; 
10'b0011011110: data <= 24'hffff6a; 
10'b0011011111: data <= 24'h000083; 
10'b0011100000: data <= 24'h0000c2; 
10'b0011100001: data <= 24'h0000c3; 
10'b0011100010: data <= 24'h000063; 
10'b0011100011: data <= 24'hffffc4; 
10'b0011100100: data <= 24'hfffe34; 
10'b0011100101: data <= 24'hfffd47; 
10'b0011100110: data <= 24'hfffcd5; 
10'b0011100111: data <= 24'hfffb92; 
10'b0011101000: data <= 24'hfffed4; 
10'b0011101001: data <= 24'hffff75; 
10'b0011101010: data <= 24'hffff5f; 
10'b0011101011: data <= 24'hfffebd; 
10'b0011101100: data <= 24'hffffe7; 
10'b0011101101: data <= 24'h0001c2; 
10'b0011101110: data <= 24'h000524; 
10'b0011101111: data <= 24'h0002d7; 
10'b0011110000: data <= 24'h0002e4; 
10'b0011110001: data <= 24'h000097; 
10'b0011110010: data <= 24'h00003a; 
10'b0011110011: data <= 24'h000027; 
10'b0011110100: data <= 24'hffff0d; 
10'b0011110101: data <= 24'h00007e; 
10'b0011110110: data <= 24'hfffec8; 
10'b0011110111: data <= 24'hfffce9; 
10'b0011111000: data <= 24'hfffd64; 
10'b0011111001: data <= 24'hfffec0; 
10'b0011111010: data <= 24'hffff74; 
10'b0011111011: data <= 24'h0000b5; 
10'b0011111100: data <= 24'h00003b; 
10'b0011111101: data <= 24'h000023; 
10'b0011111110: data <= 24'h00000d; 
10'b0011111111: data <= 24'hfffeb7; 
10'b0100000000: data <= 24'hfffd32; 
10'b0100000001: data <= 24'hfffdd9; 
10'b0100000010: data <= 24'hffff64; 
10'b0100000011: data <= 24'hfffec4; 
10'b0100000100: data <= 24'hffff44; 
10'b0100000101: data <= 24'hffffab; 
10'b0100000110: data <= 24'h000151; 
10'b0100000111: data <= 24'h0000cb; 
10'b0100001000: data <= 24'h00003c; 
10'b0100001001: data <= 24'h000220; 
10'b0100001010: data <= 24'h00038e; 
10'b0100001011: data <= 24'h00032c; 
10'b0100001100: data <= 24'hffffe0; 
10'b0100001101: data <= 24'hffff17; 
10'b0100001110: data <= 24'h000009; 
10'b0100001111: data <= 24'hfffe1b; 
10'b0100010000: data <= 24'hffff32; 
10'b0100010001: data <= 24'hfffe04; 
10'b0100010010: data <= 24'hfffde0; 
10'b0100010011: data <= 24'hfffdbc; 
10'b0100010100: data <= 24'hfffe74; 
10'b0100010101: data <= 24'hffff53; 
10'b0100010110: data <= 24'hffff82; 
10'b0100010111: data <= 24'h0000a0; 
10'b0100011000: data <= 24'h000023; 
10'b0100011001: data <= 24'hfffff9; 
10'b0100011010: data <= 24'hffffb3; 
10'b0100011011: data <= 24'hffff82; 
10'b0100011100: data <= 24'hfffdd7; 
10'b0100011101: data <= 24'hfffedf; 
10'b0100011110: data <= 24'h00010e; 
10'b0100011111: data <= 24'h000161; 
10'b0100100000: data <= 24'h0002cd; 
10'b0100100001: data <= 24'h0002c8; 
10'b0100100010: data <= 24'h000265; 
10'b0100100011: data <= 24'h00039b; 
10'b0100100100: data <= 24'h0001d1; 
10'b0100100101: data <= 24'h00006d; 
10'b0100100110: data <= 24'h000077; 
10'b0100100111: data <= 24'hfffe2d; 
10'b0100101000: data <= 24'hfffee9; 
10'b0100101001: data <= 24'hffffc9; 
10'b0100101010: data <= 24'h000145; 
10'b0100101011: data <= 24'hfffff9; 
10'b0100101100: data <= 24'h000106; 
10'b0100101101: data <= 24'hffff64; 
10'b0100101110: data <= 24'hfffebf; 
10'b0100101111: data <= 24'hfffed1; 
10'b0100110000: data <= 24'hfffe7f; 
10'b0100110001: data <= 24'hffff92; 
10'b0100110010: data <= 24'hffff6e; 
10'b0100110011: data <= 24'h00005c; 
10'b0100110100: data <= 24'hffffe2; 
10'b0100110101: data <= 24'h000025; 
10'b0100110110: data <= 24'hffffad; 
10'b0100110111: data <= 24'hffffcb; 
10'b0100111000: data <= 24'hffff68; 
10'b0100111001: data <= 24'h0001fd; 
10'b0100111010: data <= 24'h000499; 
10'b0100111011: data <= 24'h00036f; 
10'b0100111100: data <= 24'h000564; 
10'b0100111101: data <= 24'h000229; 
10'b0100111110: data <= 24'h00023e; 
10'b0100111111: data <= 24'h0003da; 
10'b0101000000: data <= 24'hfffec6; 
10'b0101000001: data <= 24'hfffef5; 
10'b0101000010: data <= 24'hffff70; 
10'b0101000011: data <= 24'h000046; 
10'b0101000100: data <= 24'h00017d; 
10'b0101000101: data <= 24'h000536; 
10'b0101000110: data <= 24'h000276; 
10'b0101000111: data <= 24'h00027f; 
10'b0101001000: data <= 24'h000418; 
10'b0101001001: data <= 24'h0002f6; 
10'b0101001010: data <= 24'h0001bb; 
10'b0101001011: data <= 24'h00005c; 
10'b0101001100: data <= 24'hffffb8; 
10'b0101001101: data <= 24'hffff4b; 
10'b0101001110: data <= 24'hfffff8; 
10'b0101001111: data <= 24'h000001; 
10'b0101010000: data <= 24'h000053; 
10'b0101010001: data <= 24'h0000ac; 
10'b0101010010: data <= 24'hffff8a; 
10'b0101010011: data <= 24'hffff43; 
10'b0101010100: data <= 24'h0001ad; 
10'b0101010101: data <= 24'h00045c; 
10'b0101010110: data <= 24'h00050b; 
10'b0101010111: data <= 24'h0002fe; 
10'b0101011000: data <= 24'h0003bd; 
10'b0101011001: data <= 24'h000493; 
10'b0101011010: data <= 24'h0002ec; 
10'b0101011011: data <= 24'h000009; 
10'b0101011100: data <= 24'hfffd12; 
10'b0101011101: data <= 24'h00028a; 
10'b0101011110: data <= 24'h00057c; 
10'b0101011111: data <= 24'h000457; 
10'b0101100000: data <= 24'h0003b6; 
10'b0101100001: data <= 24'h0005ac; 
10'b0101100010: data <= 24'h0005b6; 
10'b0101100011: data <= 24'h0005ed; 
10'b0101100100: data <= 24'h000618; 
10'b0101100101: data <= 24'h000412; 
10'b0101100110: data <= 24'h0001f5; 
10'b0101100111: data <= 24'h00000d; 
10'b0101101000: data <= 24'hffff18; 
10'b0101101001: data <= 24'h000026; 
10'b0101101010: data <= 24'h000054; 
10'b0101101011: data <= 24'h00005b; 
10'b0101101100: data <= 24'h0000c1; 
10'b0101101101: data <= 24'h000077; 
10'b0101101110: data <= 24'hffff5e; 
10'b0101101111: data <= 24'h00003d; 
10'b0101110000: data <= 24'h000289; 
10'b0101110001: data <= 24'h0003d1; 
10'b0101110010: data <= 24'h000398; 
10'b0101110011: data <= 24'h00025c; 
10'b0101110100: data <= 24'h0002f7; 
10'b0101110101: data <= 24'h0001e7; 
10'b0101110110: data <= 24'h0001b8; 
10'b0101110111: data <= 24'hffff1c; 
10'b0101111000: data <= 24'hfffe76; 
10'b0101111001: data <= 24'h0003fd; 
10'b0101111010: data <= 24'h000579; 
10'b0101111011: data <= 24'h0003f7; 
10'b0101111100: data <= 24'h000492; 
10'b0101111101: data <= 24'h000419; 
10'b0101111110: data <= 24'h00059f; 
10'b0101111111: data <= 24'h0005b8; 
10'b0110000000: data <= 24'h000478; 
10'b0110000001: data <= 24'h00029c; 
10'b0110000010: data <= 24'h000026; 
10'b0110000011: data <= 24'hfffe39; 
10'b0110000100: data <= 24'hfffef7; 
10'b0110000101: data <= 24'hffffae; 
10'b0110000110: data <= 24'h000056; 
10'b0110000111: data <= 24'h000058; 
10'b0110001000: data <= 24'h000027; 
10'b0110001001: data <= 24'h000013; 
10'b0110001010: data <= 24'h000085; 
10'b0110001011: data <= 24'h000054; 
10'b0110001100: data <= 24'h000129; 
10'b0110001101: data <= 24'h000118; 
10'b0110001110: data <= 24'h0002fb; 
10'b0110001111: data <= 24'h000216; 
10'b0110010000: data <= 24'h000103; 
10'b0110010001: data <= 24'hfffffd; 
10'b0110010010: data <= 24'h00005f; 
10'b0110010011: data <= 24'hffffd1; 
10'b0110010100: data <= 24'hfffee0; 
10'b0110010101: data <= 24'h00014b; 
10'b0110010110: data <= 24'h0000bc; 
10'b0110010111: data <= 24'h000380; 
10'b0110011000: data <= 24'h0003b6; 
10'b0110011001: data <= 24'h0003b7; 
10'b0110011010: data <= 24'h000288; 
10'b0110011011: data <= 24'h0001a0; 
10'b0110011100: data <= 24'h000208; 
10'b0110011101: data <= 24'h00000a; 
10'b0110011110: data <= 24'hfffdf3; 
10'b0110011111: data <= 24'hfffd06; 
10'b0110100000: data <= 24'hfffec5; 
10'b0110100001: data <= 24'h000035; 
10'b0110100010: data <= 24'h00001e; 
10'b0110100011: data <= 24'h000024; 
10'b0110100100: data <= 24'h000092; 
10'b0110100101: data <= 24'h000085; 
10'b0110100110: data <= 24'h000058; 
10'b0110100111: data <= 24'hffff95; 
10'b0110101000: data <= 24'h000016; 
10'b0110101001: data <= 24'h000153; 
10'b0110101010: data <= 24'h000145; 
10'b0110101011: data <= 24'h0000d7; 
10'b0110101100: data <= 24'h0000db; 
10'b0110101101: data <= 24'hfffe6e; 
10'b0110101110: data <= 24'hffff45; 
10'b0110101111: data <= 24'hffff44; 
10'b0110110000: data <= 24'hfffee7; 
10'b0110110001: data <= 24'hffff27; 
10'b0110110010: data <= 24'hfffef9; 
10'b0110110011: data <= 24'h0003d3; 
10'b0110110100: data <= 24'h000599; 
10'b0110110101: data <= 24'h00055d; 
10'b0110110110: data <= 24'h0002af; 
10'b0110110111: data <= 24'h000042; 
10'b0110111000: data <= 24'hfffed5; 
10'b0110111001: data <= 24'hfffced; 
10'b0110111010: data <= 24'hfffc2a; 
10'b0110111011: data <= 24'hfffd42; 
10'b0110111100: data <= 24'hfffec8; 
10'b0110111101: data <= 24'h000006; 
10'b0110111110: data <= 24'h000050; 
10'b0110111111: data <= 24'hfffff5; 
10'b0111000000: data <= 24'h0000a8; 
10'b0111000001: data <= 24'h00000e; 
10'b0111000010: data <= 24'hffff88; 
10'b0111000011: data <= 24'hffffe1; 
10'b0111000100: data <= 24'h00000b; 
10'b0111000101: data <= 24'h000066; 
10'b0111000110: data <= 24'hfffefa; 
10'b0111000111: data <= 24'h0000cf; 
10'b0111001000: data <= 24'h00024d; 
10'b0111001001: data <= 24'hffff76; 
10'b0111001010: data <= 24'h00014e; 
10'b0111001011: data <= 24'h0001da; 
10'b0111001100: data <= 24'hffffbf; 
10'b0111001101: data <= 24'hfffde5; 
10'b0111001110: data <= 24'hffffa6; 
10'b0111001111: data <= 24'h00021f; 
10'b0111010000: data <= 24'h0003d2; 
10'b0111010001: data <= 24'h0003cb; 
10'b0111010010: data <= 24'h0000f3; 
10'b0111010011: data <= 24'hfffdd8; 
10'b0111010100: data <= 24'hfffc6b; 
10'b0111010101: data <= 24'hfffb0d; 
10'b0111010110: data <= 24'hfffc86; 
10'b0111010111: data <= 24'hfffd2d; 
10'b0111011000: data <= 24'hfffe22; 
10'b0111011001: data <= 24'h000010; 
10'b0111011010: data <= 24'hffff98; 
10'b0111011011: data <= 24'h00005a; 
10'b0111011100: data <= 24'h000038; 
10'b0111011101: data <= 24'hffffdb; 
10'b0111011110: data <= 24'hffff7c; 
10'b0111011111: data <= 24'hffff40; 
10'b0111100000: data <= 24'hfffe98; 
10'b0111100001: data <= 24'hfffe4a; 
10'b0111100010: data <= 24'hfffe97; 
10'b0111100011: data <= 24'h0000a3; 
10'b0111100100: data <= 24'h00013d; 
10'b0111100101: data <= 24'h000169; 
10'b0111100110: data <= 24'h000227; 
10'b0111100111: data <= 24'h000322; 
10'b0111101000: data <= 24'h0001e9; 
10'b0111101001: data <= 24'h0000e3; 
10'b0111101010: data <= 24'h000137; 
10'b0111101011: data <= 24'h00031d; 
10'b0111101100: data <= 24'h0000ed; 
10'b0111101101: data <= 24'hffff5e; 
10'b0111101110: data <= 24'hfffea0; 
10'b0111101111: data <= 24'hfffcd7; 
10'b0111110000: data <= 24'hfffce1; 
10'b0111110001: data <= 24'hfffca4; 
10'b0111110010: data <= 24'hfffcd7; 
10'b0111110011: data <= 24'hfffdac; 
10'b0111110100: data <= 24'hfffe4e; 
10'b0111110101: data <= 24'h00002b; 
10'b0111110110: data <= 24'h00002d; 
10'b0111110111: data <= 24'hffffda; 
10'b0111111000: data <= 24'h00009b; 
10'b0111111001: data <= 24'h000000; 
10'b0111111010: data <= 24'hffffa5; 
10'b0111111011: data <= 24'hffffdc; 
10'b0111111100: data <= 24'hfffec3; 
10'b0111111101: data <= 24'hfffd29; 
10'b0111111110: data <= 24'hfffd1b; 
10'b0111111111: data <= 24'hfffd29; 
10'b1000000000: data <= 24'hfffecf; 
10'b1000000001: data <= 24'h000079; 
10'b1000000010: data <= 24'h00036e; 
10'b1000000011: data <= 24'h0002c6; 
10'b1000000100: data <= 24'hfffe4f; 
10'b1000000101: data <= 24'hfffe48; 
10'b1000000110: data <= 24'h00001b; 
10'b1000000111: data <= 24'h000210; 
10'b1000001000: data <= 24'hfffebd; 
10'b1000001001: data <= 24'hfffe8f; 
10'b1000001010: data <= 24'hfffd4d; 
10'b1000001011: data <= 24'hfffe60; 
10'b1000001100: data <= 24'hfffe7a; 
10'b1000001101: data <= 24'hfffd9f; 
10'b1000001110: data <= 24'hfffd80; 
10'b1000001111: data <= 24'hfffd61; 
10'b1000010000: data <= 24'hfffe26; 
10'b1000010001: data <= 24'hffffb5; 
10'b1000010010: data <= 24'h00000a; 
10'b1000010011: data <= 24'h00008e; 
10'b1000010100: data <= 24'h000065; 
10'b1000010101: data <= 24'h0000c9; 
10'b1000010110: data <= 24'h000024; 
10'b1000010111: data <= 24'hffff52; 
10'b1000011000: data <= 24'hfffedd; 
10'b1000011001: data <= 24'hfffdfd; 
10'b1000011010: data <= 24'hfffcd3; 
10'b1000011011: data <= 24'hfffcbd; 
10'b1000011100: data <= 24'hfffca0; 
10'b1000011101: data <= 24'hfffca7; 
10'b1000011110: data <= 24'hfffc41; 
10'b1000011111: data <= 24'hfffcd6; 
10'b1000100000: data <= 24'hfffbe7; 
10'b1000100001: data <= 24'hfffd23; 
10'b1000100010: data <= 24'hfffd96; 
10'b1000100011: data <= 24'hfffd41; 
10'b1000100100: data <= 24'hfffda1; 
10'b1000100101: data <= 24'hffff3a; 
10'b1000100110: data <= 24'hfffe32; 
10'b1000100111: data <= 24'hffff7f; 
10'b1000101000: data <= 24'hfffecb; 
10'b1000101001: data <= 24'hfffe92; 
10'b1000101010: data <= 24'hfffea7; 
10'b1000101011: data <= 24'hfffecd; 
10'b1000101100: data <= 24'hffff3f; 
10'b1000101101: data <= 24'h000038; 
10'b1000101110: data <= 24'hffffc3; 
10'b1000101111: data <= 24'h000016; 
10'b1000110000: data <= 24'hffffda; 
10'b1000110001: data <= 24'h00001c; 
10'b1000110010: data <= 24'h000055; 
10'b1000110011: data <= 24'h000007; 
10'b1000110100: data <= 24'hfffed3; 
10'b1000110101: data <= 24'hfffe0f; 
10'b1000110110: data <= 24'hfffd0f; 
10'b1000110111: data <= 24'hfffb64; 
10'b1000111000: data <= 24'hfffab8; 
10'b1000111001: data <= 24'hfffa14; 
10'b1000111010: data <= 24'hfff7fb; 
10'b1000111011: data <= 24'hfff9dd; 
10'b1000111100: data <= 24'hfffa05; 
10'b1000111101: data <= 24'hfffe0b; 
10'b1000111110: data <= 24'hfffd41; 
10'b1000111111: data <= 24'hfffeb6; 
10'b1001000000: data <= 24'hfffe74; 
10'b1001000001: data <= 24'hffff95; 
10'b1001000010: data <= 24'hfffd5f; 
10'b1001000011: data <= 24'hffff22; 
10'b1001000100: data <= 24'hfffef5; 
10'b1001000101: data <= 24'hfffe53; 
10'b1001000110: data <= 24'hffff87; 
10'b1001000111: data <= 24'hffff33; 
10'b1001001000: data <= 24'h000015; 
10'b1001001001: data <= 24'h0000ab; 
10'b1001001010: data <= 24'h000067; 
10'b1001001011: data <= 24'h000020; 
10'b1001001100: data <= 24'h00000e; 
10'b1001001101: data <= 24'h000000; 
10'b1001001110: data <= 24'h0000ab; 
10'b1001001111: data <= 24'hffff4b; 
10'b1001010000: data <= 24'hffff36; 
10'b1001010001: data <= 24'hfffe16; 
10'b1001010010: data <= 24'hfffd4c; 
10'b1001010011: data <= 24'hfffbd4; 
10'b1001010100: data <= 24'hfffb44; 
10'b1001010101: data <= 24'hfffaca; 
10'b1001010110: data <= 24'hfffa8a; 
10'b1001010111: data <= 24'hfffb17; 
10'b1001011000: data <= 24'hfffcdf; 
10'b1001011001: data <= 24'hfffce9; 
10'b1001011010: data <= 24'hfffcdc; 
10'b1001011011: data <= 24'hfffe33; 
10'b1001011100: data <= 24'hfffe0c; 
10'b1001011101: data <= 24'hfffd10; 
10'b1001011110: data <= 24'hfffc75; 
10'b1001011111: data <= 24'hfffe80; 
10'b1001100000: data <= 24'hffff2a; 
10'b1001100001: data <= 24'hffff84; 
10'b1001100010: data <= 24'h00003d; 
10'b1001100011: data <= 24'hffffef; 
10'b1001100100: data <= 24'h00004d; 
10'b1001100101: data <= 24'h000069; 
10'b1001100110: data <= 24'h000006; 
10'b1001100111: data <= 24'h00000d; 
10'b1001101000: data <= 24'h000083; 
10'b1001101001: data <= 24'h000021; 
10'b1001101010: data <= 24'h000025; 
10'b1001101011: data <= 24'h00007e; 
10'b1001101100: data <= 24'hffffaf; 
10'b1001101101: data <= 24'hfffe74; 
10'b1001101110: data <= 24'hfffd87; 
10'b1001101111: data <= 24'hfffca3; 
10'b1001110000: data <= 24'hfffd7f; 
10'b1001110001: data <= 24'hfffd62; 
10'b1001110010: data <= 24'hfffd25; 
10'b1001110011: data <= 24'hfffe12; 
10'b1001110100: data <= 24'hfffdd5; 
10'b1001110101: data <= 24'hfffd1d; 
10'b1001110110: data <= 24'hfffd93; 
10'b1001110111: data <= 24'hfffc9a; 
10'b1001111000: data <= 24'hfffc3e; 
10'b1001111001: data <= 24'hfffc51; 
10'b1001111010: data <= 24'hfffcef; 
10'b1001111011: data <= 24'hfffd46; 
10'b1001111100: data <= 24'hffff41; 
10'b1001111101: data <= 24'h0000eb; 
10'b1001111110: data <= 24'h000082; 
10'b1001111111: data <= 24'h0000a2; 
10'b1010000000: data <= 24'h000109; 
10'b1010000001: data <= 24'h000038; 
10'b1010000010: data <= 24'h00003e; 
10'b1010000011: data <= 24'h000061; 
10'b1010000100: data <= 24'h00009a; 
10'b1010000101: data <= 24'h000079; 
10'b1010000110: data <= 24'h00002d; 
10'b1010000111: data <= 24'hffffc4; 
10'b1010001000: data <= 24'hffff91; 
10'b1010001001: data <= 24'hfffeac; 
10'b1010001010: data <= 24'hfffe74; 
10'b1010001011: data <= 24'hfffdf5; 
10'b1010001100: data <= 24'hffffd8; 
10'b1010001101: data <= 24'hffff2c; 
10'b1010001110: data <= 24'hffff57; 
10'b1010001111: data <= 24'hfffd86; 
10'b1010010000: data <= 24'hfffdfb; 
10'b1010010001: data <= 24'hfffd74; 
10'b1010010010: data <= 24'hfffdd9; 
10'b1010010011: data <= 24'hfffc53; 
10'b1010010100: data <= 24'hfffc08; 
10'b1010010101: data <= 24'hfffc82; 
10'b1010010110: data <= 24'hfffdd3; 
10'b1010010111: data <= 24'hffffca; 
10'b1010011000: data <= 24'h0000da; 
10'b1010011001: data <= 24'h0001fa; 
10'b1010011010: data <= 24'h0002da; 
10'b1010011011: data <= 24'h000263; 
10'b1010011100: data <= 24'h00011e; 
10'b1010011101: data <= 24'hffffec; 
10'b1010011110: data <= 24'h0000cd; 
10'b1010011111: data <= 24'hffffe8; 
10'b1010100000: data <= 24'hffffff; 
10'b1010100001: data <= 24'hffffaf; 
10'b1010100010: data <= 24'hffffea; 
10'b1010100011: data <= 24'h0000ad; 
10'b1010100100: data <= 24'h00007c; 
10'b1010100101: data <= 24'h0000c3; 
10'b1010100110: data <= 24'h00008d; 
10'b1010100111: data <= 24'h0000cd; 
10'b1010101000: data <= 24'h000122; 
10'b1010101001: data <= 24'h00009d; 
10'b1010101010: data <= 24'hffff99; 
10'b1010101011: data <= 24'hfffebb; 
10'b1010101100: data <= 24'hffffe9; 
10'b1010101101: data <= 24'hfffe0d; 
10'b1010101110: data <= 24'hfffd89; 
10'b1010101111: data <= 24'hfffd66; 
10'b1010110000: data <= 24'hfffed2; 
10'b1010110001: data <= 24'h0000db; 
10'b1010110010: data <= 24'h000176; 
10'b1010110011: data <= 24'h000183; 
10'b1010110100: data <= 24'h000373; 
10'b1010110101: data <= 24'h0003b6; 
10'b1010110110: data <= 24'h000223; 
10'b1010110111: data <= 24'h00014e; 
10'b1010111000: data <= 24'h000108; 
10'b1010111001: data <= 24'hffffcc; 
10'b1010111010: data <= 24'h000076; 
10'b1010111011: data <= 24'hfffff8; 
10'b1010111100: data <= 24'h00002b; 
10'b1010111101: data <= 24'h0000ab; 
10'b1010111110: data <= 24'h0000ac; 
10'b1010111111: data <= 24'hffffee; 
10'b1011000000: data <= 24'h000010; 
10'b1011000001: data <= 24'h000125; 
10'b1011000010: data <= 24'h0000de; 
10'b1011000011: data <= 24'h000281; 
10'b1011000100: data <= 24'h0002bf; 
10'b1011000101: data <= 24'h0002cb; 
10'b1011000110: data <= 24'h00026b; 
10'b1011000111: data <= 24'h0000f6; 
10'b1011001000: data <= 24'h00028b; 
10'b1011001001: data <= 24'h000245; 
10'b1011001010: data <= 24'h00022c; 
10'b1011001011: data <= 24'h00020b; 
10'b1011001100: data <= 24'h0003d1; 
10'b1011001101: data <= 24'h000425; 
10'b1011001110: data <= 24'h00048f; 
10'b1011001111: data <= 24'h0004c2; 
10'b1011010000: data <= 24'h000550; 
10'b1011010001: data <= 24'h0003c5; 
10'b1011010010: data <= 24'h000178; 
10'b1011010011: data <= 24'h0000b3; 
10'b1011010100: data <= 24'hffffe8; 
10'b1011010101: data <= 24'hfffff2; 
10'b1011010110: data <= 24'h000032; 
10'b1011010111: data <= 24'h00002a; 
10'b1011011000: data <= 24'h000007; 
10'b1011011001: data <= 24'h00009c; 
10'b1011011010: data <= 24'h00002a; 
10'b1011011011: data <= 24'hffffc7; 
10'b1011011100: data <= 24'h00009d; 
10'b1011011101: data <= 24'h0000f3; 
10'b1011011110: data <= 24'h000155; 
10'b1011011111: data <= 24'h0001da; 
10'b1011100000: data <= 24'h00021c; 
10'b1011100001: data <= 24'h000332; 
10'b1011100010: data <= 24'h00034c; 
10'b1011100011: data <= 24'h0003b4; 
10'b1011100100: data <= 24'h000463; 
10'b1011100101: data <= 24'h00046d; 
10'b1011100110: data <= 24'h00056b; 
10'b1011100111: data <= 24'h000320; 
10'b1011101000: data <= 24'h000224; 
10'b1011101001: data <= 24'h0001cf; 
10'b1011101010: data <= 24'h0002ab; 
10'b1011101011: data <= 24'h0002e1; 
10'b1011101100: data <= 24'h000217; 
10'b1011101101: data <= 24'h000175; 
10'b1011101110: data <= 24'h00009b; 
10'b1011101111: data <= 24'h000038; 
10'b1011110000: data <= 24'h000023; 
10'b1011110001: data <= 24'h00003e; 
10'b1011110010: data <= 24'hffffc5; 
10'b1011110011: data <= 24'h000022; 
10'b1011110100: data <= 24'hffffdb; 
10'b1011110101: data <= 24'h000047; 
10'b1011110110: data <= 24'hffffc0; 
10'b1011110111: data <= 24'h0000bd; 
10'b1011111000: data <= 24'h00006d; 
10'b1011111001: data <= 24'h00003c; 
10'b1011111010: data <= 24'hffffe5; 
10'b1011111011: data <= 24'h0000b8; 
10'b1011111100: data <= 24'h00009b; 
10'b1011111101: data <= 24'h00006a; 
10'b1011111110: data <= 24'hffffde; 
10'b1011111111: data <= 24'hffffda; 
10'b1100000000: data <= 24'h000025; 
10'b1100000001: data <= 24'hffffde; 
10'b1100000010: data <= 24'h000028; 
10'b1100000011: data <= 24'h000076; 
10'b1100000100: data <= 24'h00000b; 
10'b1100000101: data <= 24'h000040; 
10'b1100000110: data <= 24'h0000d2; 
10'b1100000111: data <= 24'h0000bb; 
10'b1100001000: data <= 24'h000069; 
10'b1100001001: data <= 24'h000040; 
10'b1100001010: data <= 24'hffffcc; 
10'b1100001011: data <= 24'h0000cf; 
10'b1100001100: data <= 24'h000071; 
10'b1100001101: data <= 24'hffffda; 
10'b1100001110: data <= 24'h00000e; 
10'b1100001111: data <= 24'hffffeb; 
endcase
end

assign dout = data;

endmodule