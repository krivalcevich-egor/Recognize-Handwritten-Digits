`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// WEIGHT MEMORY
// This code create bram for 1 of 10 weights strings
// and send element with input address from the string to out.
//////////////////////////////////////////////////////////////////////////////////

module ROM_weights_7 #( 
    parameter int BITS = 24 // bit depth
)(
    input logic clk, // clock
    input logic [9:0] address, // address of current element from string
    output [BITS-1:0] dout // current element from string
);

(* rom_style = "block" *) reg [BITS-1:0] data;

always @(posedge clk)
begin
case(address)
10'b0000000000: data <= 24'h00000c; 
10'b0000000001: data <= 24'h000010; 
10'b0000000010: data <= 24'h000079; 
10'b0000000011: data <= 24'h00002f; 
10'b0000000100: data <= 24'h0000c6; 
10'b0000000101: data <= 24'hffffa8; 
10'b0000000110: data <= 24'hffffc5; 
10'b0000000111: data <= 24'h000040; 
10'b0000001000: data <= 24'h000098; 
10'b0000001001: data <= 24'h000095; 
10'b0000001010: data <= 24'hffffac; 
10'b0000001011: data <= 24'h000028; 
10'b0000001100: data <= 24'h00002b; 
10'b0000001101: data <= 24'hffffea; 
10'b0000001110: data <= 24'h00009f; 
10'b0000001111: data <= 24'h00002b; 
10'b0000010000: data <= 24'h000003; 
10'b0000010001: data <= 24'hfffffa; 
10'b0000010010: data <= 24'h000011; 
10'b0000010011: data <= 24'h000037; 
10'b0000010100: data <= 24'h000066; 
10'b0000010101: data <= 24'h0000c2; 
10'b0000010110: data <= 24'hffffcc; 
10'b0000010111: data <= 24'h00008f; 
10'b0000011000: data <= 24'hffffec; 
10'b0000011001: data <= 24'h000066; 
10'b0000011010: data <= 24'hfffff8; 
10'b0000011011: data <= 24'hffffff; 
10'b0000011100: data <= 24'h0000b7; 
10'b0000011101: data <= 24'hffffd9; 
10'b0000011110: data <= 24'h000029; 
10'b0000011111: data <= 24'h0000b4; 
10'b0000100000: data <= 24'h000045; 
10'b0000100001: data <= 24'h000007; 
10'b0000100010: data <= 24'h0000b3; 
10'b0000100011: data <= 24'h000038; 
10'b0000100100: data <= 24'h000011; 
10'b0000100101: data <= 24'hffffe2; 
10'b0000100110: data <= 24'hffffe8; 
10'b0000100111: data <= 24'hffffa2; 
10'b0000101000: data <= 24'h00009a; 
10'b0000101001: data <= 24'hfffff5; 
10'b0000101010: data <= 24'h0000b8; 
10'b0000101011: data <= 24'hffffd0; 
10'b0000101100: data <= 24'h000050; 
10'b0000101101: data <= 24'h00008b; 
10'b0000101110: data <= 24'h00009c; 
10'b0000101111: data <= 24'h00007c; 
10'b0000110000: data <= 24'h000004; 
10'b0000110001: data <= 24'h00007b; 
10'b0000110010: data <= 24'hfffffc; 
10'b0000110011: data <= 24'h0000c2; 
10'b0000110100: data <= 24'h000096; 
10'b0000110101: data <= 24'hffffca; 
10'b0000110110: data <= 24'hffffcb; 
10'b0000110111: data <= 24'h00004f; 
10'b0000111000: data <= 24'h0000ad; 
10'b0000111001: data <= 24'h0000aa; 
10'b0000111010: data <= 24'h000086; 
10'b0000111011: data <= 24'hffffe7; 
10'b0000111100: data <= 24'h00009b; 
10'b0000111101: data <= 24'hffffb6; 
10'b0000111110: data <= 24'hffffc3; 
10'b0000111111: data <= 24'h00007a; 
10'b0001000000: data <= 24'h000067; 
10'b0001000001: data <= 24'hffffc4; 
10'b0001000010: data <= 24'hfffff3; 
10'b0001000011: data <= 24'h00004c; 
10'b0001000100: data <= 24'hffffeb; 
10'b0001000101: data <= 24'hffffd8; 
10'b0001000110: data <= 24'h000030; 
10'b0001000111: data <= 24'h00009c; 
10'b0001001000: data <= 24'h00007e; 
10'b0001001001: data <= 24'h000017; 
10'b0001001010: data <= 24'h00003e; 
10'b0001001011: data <= 24'h0000b1; 
10'b0001001100: data <= 24'h000096; 
10'b0001001101: data <= 24'h0000ae; 
10'b0001001110: data <= 24'hffffa9; 
10'b0001001111: data <= 24'h000087; 
10'b0001010000: data <= 24'h000033; 
10'b0001010001: data <= 24'h000078; 
10'b0001010010: data <= 24'h000067; 
10'b0001010011: data <= 24'h000098; 
10'b0001010100: data <= 24'hfffff2; 
10'b0001010101: data <= 24'h00000a; 
10'b0001010110: data <= 24'h00009e; 
10'b0001010111: data <= 24'hffffe8; 
10'b0001011000: data <= 24'h000012; 
10'b0001011001: data <= 24'hfffff5; 
10'b0001011010: data <= 24'hffffc6; 
10'b0001011011: data <= 24'h000067; 
10'b0001011100: data <= 24'h000001; 
10'b0001011101: data <= 24'h000067; 
10'b0001011110: data <= 24'hffffab; 
10'b0001011111: data <= 24'h000015; 
10'b0001100000: data <= 24'h000053; 
10'b0001100001: data <= 24'hffff8e; 
10'b0001100010: data <= 24'h00005e; 
10'b0001100011: data <= 24'hffffb3; 
10'b0001100100: data <= 24'hffff58; 
10'b0001100101: data <= 24'hffff77; 
10'b0001100110: data <= 24'hffff8a; 
10'b0001100111: data <= 24'hffffb1; 
10'b0001101000: data <= 24'hffffec; 
10'b0001101001: data <= 24'hffffb7; 
10'b0001101010: data <= 24'h000040; 
10'b0001101011: data <= 24'hfffff8; 
10'b0001101100: data <= 24'h00004d; 
10'b0001101101: data <= 24'h0000c3; 
10'b0001101110: data <= 24'hffffc0; 
10'b0001101111: data <= 24'h000051; 
10'b0001110000: data <= 24'h0000bd; 
10'b0001110001: data <= 24'hffffbb; 
10'b0001110010: data <= 24'h000069; 
10'b0001110011: data <= 24'hffffb0; 
10'b0001110100: data <= 24'h00002c; 
10'b0001110101: data <= 24'hffffdc; 
10'b0001110110: data <= 24'h000008; 
10'b0001110111: data <= 24'hffffb2; 
10'b0001111000: data <= 24'h00003b; 
10'b0001111001: data <= 24'hffffe4; 
10'b0001111010: data <= 24'hffff47; 
10'b0001111011: data <= 24'hfffe9b; 
10'b0001111100: data <= 24'hfffe89; 
10'b0001111101: data <= 24'hfffe9a; 
10'b0001111110: data <= 24'hfffe55; 
10'b0001111111: data <= 24'hfffd41; 
10'b0010000000: data <= 24'hfffe61; 
10'b0010000001: data <= 24'hfffec8; 
10'b0010000010: data <= 24'hfffef1; 
10'b0010000011: data <= 24'hffffb7; 
10'b0010000100: data <= 24'hffff35; 
10'b0010000101: data <= 24'h00005e; 
10'b0010000110: data <= 24'h00000e; 
10'b0010000111: data <= 24'hffff9e; 
10'b0010001000: data <= 24'h0000b3; 
10'b0010001001: data <= 24'hfffffa; 
10'b0010001010: data <= 24'h0000b0; 
10'b0010001011: data <= 24'h0000aa; 
10'b0010001100: data <= 24'h0000a1; 
10'b0010001101: data <= 24'h000006; 
10'b0010001110: data <= 24'h00009b; 
10'b0010001111: data <= 24'hffffd6; 
10'b0010010000: data <= 24'hffff86; 
10'b0010010001: data <= 24'hffffeb; 
10'b0010010010: data <= 24'hffffa3; 
10'b0010010011: data <= 24'hffffde; 
10'b0010010100: data <= 24'hffff92; 
10'b0010010101: data <= 24'hffff00; 
10'b0010010110: data <= 24'hfffd8a; 
10'b0010010111: data <= 24'hfffcfb; 
10'b0010011000: data <= 24'hfffc33; 
10'b0010011001: data <= 24'hfffb8d; 
10'b0010011010: data <= 24'hfffa72; 
10'b0010011011: data <= 24'hfffa7d; 
10'b0010011100: data <= 24'hfffa38; 
10'b0010011101: data <= 24'hfffae6; 
10'b0010011110: data <= 24'hfffbae; 
10'b0010011111: data <= 24'hfffcb6; 
10'b0010100000: data <= 24'hfffdaa; 
10'b0010100001: data <= 24'hffff2b; 
10'b0010100010: data <= 24'hfffeb6; 
10'b0010100011: data <= 24'hffffd7; 
10'b0010100100: data <= 24'h000090; 
10'b0010100101: data <= 24'h000073; 
10'b0010100110: data <= 24'hffffe2; 
10'b0010100111: data <= 24'h000006; 
10'b0010101000: data <= 24'h000086; 
10'b0010101001: data <= 24'h0000b8; 
10'b0010101010: data <= 24'h00000d; 
10'b0010101011: data <= 24'h00001e; 
10'b0010101100: data <= 24'h0000c7; 
10'b0010101101: data <= 24'h0000ec; 
10'b0010101110: data <= 24'h000115; 
10'b0010101111: data <= 24'h0001a1; 
10'b0010110000: data <= 24'h00026a; 
10'b0010110001: data <= 24'h0001ef; 
10'b0010110010: data <= 24'h00020f; 
10'b0010110011: data <= 24'h00005f; 
10'b0010110100: data <= 24'hfffe59; 
10'b0010110101: data <= 24'hfffc89; 
10'b0010110110: data <= 24'hfffc62; 
10'b0010110111: data <= 24'hfffe1f; 
10'b0010111000: data <= 24'hfffedc; 
10'b0010111001: data <= 24'hfffea6; 
10'b0010111010: data <= 24'hfffe5c; 
10'b0010111011: data <= 24'hfffe1a; 
10'b0010111100: data <= 24'hfffd20; 
10'b0010111101: data <= 24'hfffeec; 
10'b0010111110: data <= 24'hfffdfc; 
10'b0010111111: data <= 24'hfffe89; 
10'b0011000000: data <= 24'hffff05; 
10'b0011000001: data <= 24'hffffac; 
10'b0011000010: data <= 24'hffffa9; 
10'b0011000011: data <= 24'h000014; 
10'b0011000100: data <= 24'h00007a; 
10'b0011000101: data <= 24'h0000b9; 
10'b0011000110: data <= 24'h000098; 
10'b0011000111: data <= 24'h000168; 
10'b0011001000: data <= 24'h0001b5; 
10'b0011001001: data <= 24'h000189; 
10'b0011001010: data <= 24'h000239; 
10'b0011001011: data <= 24'h000365; 
10'b0011001100: data <= 24'h0004a7; 
10'b0011001101: data <= 24'h0003af; 
10'b0011001110: data <= 24'h00028b; 
10'b0011001111: data <= 24'h0002cd; 
10'b0011010000: data <= 24'h0002fc; 
10'b0011010001: data <= 24'h000093; 
10'b0011010010: data <= 24'h00006c; 
10'b0011010011: data <= 24'h000111; 
10'b0011010100: data <= 24'h000326; 
10'b0011010101: data <= 24'h000380; 
10'b0011010110: data <= 24'h00025f; 
10'b0011010111: data <= 24'h0001e7; 
10'b0011011000: data <= 24'h000077; 
10'b0011011001: data <= 24'hffff79; 
10'b0011011010: data <= 24'h00003f; 
10'b0011011011: data <= 24'hffff6f; 
10'b0011011100: data <= 24'hffff78; 
10'b0011011101: data <= 24'hfffff9; 
10'b0011011110: data <= 24'h000060; 
10'b0011011111: data <= 24'hffffdc; 
10'b0011100000: data <= 24'hffffa3; 
10'b0011100001: data <= 24'h0000c2; 
10'b0011100010: data <= 24'h00004b; 
10'b0011100011: data <= 24'h000130; 
10'b0011100100: data <= 24'h000268; 
10'b0011100101: data <= 24'h00022b; 
10'b0011100110: data <= 24'h0002e8; 
10'b0011100111: data <= 24'h000537; 
10'b0011101000: data <= 24'h000383; 
10'b0011101001: data <= 24'h00026b; 
10'b0011101010: data <= 24'h000313; 
10'b0011101011: data <= 24'h00041f; 
10'b0011101100: data <= 24'h0003eb; 
10'b0011101101: data <= 24'h0001f8; 
10'b0011101110: data <= 24'h000127; 
10'b0011101111: data <= 24'h000199; 
10'b0011110000: data <= 24'h0002c7; 
10'b0011110001: data <= 24'h000445; 
10'b0011110010: data <= 24'h0002ed; 
10'b0011110011: data <= 24'h000281; 
10'b0011110100: data <= 24'h000200; 
10'b0011110101: data <= 24'h00000c; 
10'b0011110110: data <= 24'h000136; 
10'b0011110111: data <= 24'h000107; 
10'b0011111000: data <= 24'hffff44; 
10'b0011111001: data <= 24'hffffa6; 
10'b0011111010: data <= 24'h000068; 
10'b0011111011: data <= 24'h0000a0; 
10'b0011111100: data <= 24'h000052; 
10'b0011111101: data <= 24'h00009a; 
10'b0011111110: data <= 24'h0000cf; 
10'b0011111111: data <= 24'h0001b7; 
10'b0100000000: data <= 24'h00025b; 
10'b0100000001: data <= 24'h0002ad; 
10'b0100000010: data <= 24'h0000fb; 
10'b0100000011: data <= 24'h00014e; 
10'b0100000100: data <= 24'h00017b; 
10'b0100000101: data <= 24'h0000fb; 
10'b0100000110: data <= 24'h000266; 
10'b0100000111: data <= 24'h0002f1; 
10'b0100001000: data <= 24'h0003c0; 
10'b0100001001: data <= 24'h00030d; 
10'b0100001010: data <= 24'h00045f; 
10'b0100001011: data <= 24'h000561; 
10'b0100001100: data <= 24'h0004f4; 
10'b0100001101: data <= 24'h000587; 
10'b0100001110: data <= 24'h00039c; 
10'b0100001111: data <= 24'h0003ad; 
10'b0100010000: data <= 24'h000317; 
10'b0100010001: data <= 24'h000294; 
10'b0100010010: data <= 24'h000138; 
10'b0100010011: data <= 24'hffff8e; 
10'b0100010100: data <= 24'hffff40; 
10'b0100010101: data <= 24'hffffa2; 
10'b0100010110: data <= 24'h000054; 
10'b0100010111: data <= 24'hffffd5; 
10'b0100011000: data <= 24'h000020; 
10'b0100011001: data <= 24'h0000a8; 
10'b0100011010: data <= 24'h0000bb; 
10'b0100011011: data <= 24'h000221; 
10'b0100011100: data <= 24'h000271; 
10'b0100011101: data <= 24'h000207; 
10'b0100011110: data <= 24'h000060; 
10'b0100011111: data <= 24'h00009c; 
10'b0100100000: data <= 24'hffff2e; 
10'b0100100001: data <= 24'hfffff8; 
10'b0100100010: data <= 24'h00017d; 
10'b0100100011: data <= 24'h00029f; 
10'b0100100100: data <= 24'h0001d3; 
10'b0100100101: data <= 24'h00043e; 
10'b0100100110: data <= 24'h000576; 
10'b0100100111: data <= 24'h0006b5; 
10'b0100101000: data <= 24'h0007a2; 
10'b0100101001: data <= 24'h0005a9; 
10'b0100101010: data <= 24'h000475; 
10'b0100101011: data <= 24'h0004a3; 
10'b0100101100: data <= 24'h000412; 
10'b0100101101: data <= 24'h000376; 
10'b0100101110: data <= 24'h000188; 
10'b0100101111: data <= 24'hffff60; 
10'b0100110000: data <= 24'hfffef8; 
10'b0100110001: data <= 24'hffff95; 
10'b0100110010: data <= 24'h000014; 
10'b0100110011: data <= 24'hffffd8; 
10'b0100110100: data <= 24'h000094; 
10'b0100110101: data <= 24'h000068; 
10'b0100110110: data <= 24'h0000bd; 
10'b0100110111: data <= 24'h00022e; 
10'b0100111000: data <= 24'h0002a1; 
10'b0100111001: data <= 24'h00014e; 
10'b0100111010: data <= 24'h000079; 
10'b0100111011: data <= 24'h00006d; 
10'b0100111100: data <= 24'h00001f; 
10'b0100111101: data <= 24'h000194; 
10'b0100111110: data <= 24'h0000d0; 
10'b0100111111: data <= 24'h000107; 
10'b0101000000: data <= 24'h0001b2; 
10'b0101000001: data <= 24'h0001ae; 
10'b0101000010: data <= 24'h0001c0; 
10'b0101000011: data <= 24'h000522; 
10'b0101000100: data <= 24'h0006aa; 
10'b0101000101: data <= 24'h000471; 
10'b0101000110: data <= 24'h00047c; 
10'b0101000111: data <= 24'h000373; 
10'b0101001000: data <= 24'h00035a; 
10'b0101001001: data <= 24'h00021b; 
10'b0101001010: data <= 24'h000186; 
10'b0101001011: data <= 24'hffff79; 
10'b0101001100: data <= 24'hfffe76; 
10'b0101001101: data <= 24'hfffff5; 
10'b0101001110: data <= 24'h000026; 
10'b0101001111: data <= 24'h0000ad; 
10'b0101010000: data <= 24'h000084; 
10'b0101010001: data <= 24'hfffff6; 
10'b0101010010: data <= 24'h00005e; 
10'b0101010011: data <= 24'h000160; 
10'b0101010100: data <= 24'h00018b; 
10'b0101010101: data <= 24'h000041; 
10'b0101010110: data <= 24'h000058; 
10'b0101010111: data <= 24'h000178; 
10'b0101011000: data <= 24'h000102; 
10'b0101011001: data <= 24'hfffff1; 
10'b0101011010: data <= 24'hfffecd; 
10'b0101011011: data <= 24'hfffcce; 
10'b0101011100: data <= 24'hfff93f; 
10'b0101011101: data <= 24'hfff58c; 
10'b0101011110: data <= 24'hfff82d; 
10'b0101011111: data <= 24'h00002c; 
10'b0101100000: data <= 24'h00046b; 
10'b0101100001: data <= 24'h000403; 
10'b0101100010: data <= 24'h000194; 
10'b0101100011: data <= 24'h000091; 
10'b0101100100: data <= 24'h00001b; 
10'b0101100101: data <= 24'hffff6c; 
10'b0101100110: data <= 24'hffff7a; 
10'b0101100111: data <= 24'hffff0e; 
10'b0101101000: data <= 24'hffff52; 
10'b0101101001: data <= 24'h0000a3; 
10'b0101101010: data <= 24'h000073; 
10'b0101101011: data <= 24'h000001; 
10'b0101101100: data <= 24'h00008f; 
10'b0101101101: data <= 24'h000054; 
10'b0101101110: data <= 24'h00009a; 
10'b0101101111: data <= 24'h00013f; 
10'b0101110000: data <= 24'h000077; 
10'b0101110001: data <= 24'h000033; 
10'b0101110010: data <= 24'hffff97; 
10'b0101110011: data <= 24'h000045; 
10'b0101110100: data <= 24'hffffd0; 
10'b0101110101: data <= 24'hfffefa; 
10'b0101110110: data <= 24'hfffca6; 
10'b0101110111: data <= 24'hfff8ef; 
10'b0101111000: data <= 24'hfff397; 
10'b0101111001: data <= 24'hfff224; 
10'b0101111010: data <= 24'hfff895; 
10'b0101111011: data <= 24'hffff07; 
10'b0101111100: data <= 24'h000242; 
10'b0101111101: data <= 24'h000174; 
10'b0101111110: data <= 24'h000051; 
10'b0101111111: data <= 24'h0000a9; 
10'b0110000000: data <= 24'hfffea4; 
10'b0110000001: data <= 24'hfffe43; 
10'b0110000010: data <= 24'hffff98; 
10'b0110000011: data <= 24'h000021; 
10'b0110000100: data <= 24'hffffab; 
10'b0110000101: data <= 24'hffffbc; 
10'b0110000110: data <= 24'h00005a; 
10'b0110000111: data <= 24'hffffa8; 
10'b0110001000: data <= 24'hffffda; 
10'b0110001001: data <= 24'h00004c; 
10'b0110001010: data <= 24'h00011e; 
10'b0110001011: data <= 24'h000164; 
10'b0110001100: data <= 24'h0000e2; 
10'b0110001101: data <= 24'h000106; 
10'b0110001110: data <= 24'hffffa9; 
10'b0110001111: data <= 24'hffff49; 
10'b0110010000: data <= 24'hfffe6d; 
10'b0110010001: data <= 24'hfffc51; 
10'b0110010010: data <= 24'hfffa95; 
10'b0110010011: data <= 24'hfff79f; 
10'b0110010100: data <= 24'hfff543; 
10'b0110010101: data <= 24'hfff6f1; 
10'b0110010110: data <= 24'hfffcae; 
10'b0110010111: data <= 24'h000014; 
10'b0110011000: data <= 24'h0000b1; 
10'b0110011001: data <= 24'h00016e; 
10'b0110011010: data <= 24'h00041b; 
10'b0110011011: data <= 24'h00046a; 
10'b0110011100: data <= 24'h0002a8; 
10'b0110011101: data <= 24'h0001b2; 
10'b0110011110: data <= 24'h0001b5; 
10'b0110011111: data <= 24'h00017b; 
10'b0110100000: data <= 24'h000080; 
10'b0110100001: data <= 24'h000026; 
10'b0110100010: data <= 24'hffffc4; 
10'b0110100011: data <= 24'hffffc9; 
10'b0110100100: data <= 24'h00005c; 
10'b0110100101: data <= 24'h000088; 
10'b0110100110: data <= 24'h000032; 
10'b0110100111: data <= 24'h000087; 
10'b0110101000: data <= 24'h000086; 
10'b0110101001: data <= 24'hfffe83; 
10'b0110101010: data <= 24'hffff56; 
10'b0110101011: data <= 24'hffff14; 
10'b0110101100: data <= 24'hfffc0c; 
10'b0110101101: data <= 24'hfffb34; 
10'b0110101110: data <= 24'hfff99f; 
10'b0110101111: data <= 24'hfff8b1; 
10'b0110110000: data <= 24'hfff80a; 
10'b0110110001: data <= 24'hfffa22; 
10'b0110110010: data <= 24'hfffc93; 
10'b0110110011: data <= 24'h00001b; 
10'b0110110100: data <= 24'h000060; 
10'b0110110101: data <= 24'h000595; 
10'b0110110110: data <= 24'h000689; 
10'b0110110111: data <= 24'h000563; 
10'b0110111000: data <= 24'h0004c9; 
10'b0110111001: data <= 24'h00041d; 
10'b0110111010: data <= 24'h0002a9; 
10'b0110111011: data <= 24'h000134; 
10'b0110111100: data <= 24'hfffff3; 
10'b0110111101: data <= 24'hffffab; 
10'b0110111110: data <= 24'h000017; 
10'b0110111111: data <= 24'h000093; 
10'b0111000000: data <= 24'h00005b; 
10'b0111000001: data <= 24'h0000b5; 
10'b0111000010: data <= 24'hfffff1; 
10'b0111000011: data <= 24'h0000be; 
10'b0111000100: data <= 24'h000096; 
10'b0111000101: data <= 24'hffff56; 
10'b0111000110: data <= 24'hffff0f; 
10'b0111000111: data <= 24'hffffdd; 
10'b0111001000: data <= 24'hfffcd1; 
10'b0111001001: data <= 24'hfffc68; 
10'b0111001010: data <= 24'hfffa37; 
10'b0111001011: data <= 24'hfff91f; 
10'b0111001100: data <= 24'hfffbb0; 
10'b0111001101: data <= 24'hfffd97; 
10'b0111001110: data <= 24'hfffc81; 
10'b0111001111: data <= 24'h0001cd; 
10'b0111010000: data <= 24'h00022d; 
10'b0111010001: data <= 24'h0004b9; 
10'b0111010010: data <= 24'h00040c; 
10'b0111010011: data <= 24'h00043e; 
10'b0111010100: data <= 24'h000360; 
10'b0111010101: data <= 24'h000292; 
10'b0111010110: data <= 24'h000082; 
10'b0111010111: data <= 24'hfffef1; 
10'b0111011000: data <= 24'hffff58; 
10'b0111011001: data <= 24'hffffa0; 
10'b0111011010: data <= 24'h000067; 
10'b0111011011: data <= 24'h0000b3; 
10'b0111011100: data <= 24'h000006; 
10'b0111011101: data <= 24'h000017; 
10'b0111011110: data <= 24'h00006e; 
10'b0111011111: data <= 24'hfffff8; 
10'b0111100000: data <= 24'h000024; 
10'b0111100001: data <= 24'hffff93; 
10'b0111100010: data <= 24'hfffddb; 
10'b0111100011: data <= 24'hfffd2c; 
10'b0111100100: data <= 24'hfffc74; 
10'b0111100101: data <= 24'hfffd12; 
10'b0111100110: data <= 24'hfffc1e; 
10'b0111100111: data <= 24'hfffd1e; 
10'b0111101000: data <= 24'hffff14; 
10'b0111101001: data <= 24'h0000b8; 
10'b0111101010: data <= 24'h000068; 
10'b0111101011: data <= 24'h0000b7; 
10'b0111101100: data <= 24'hffff93; 
10'b0111101101: data <= 24'h000123; 
10'b0111101110: data <= 24'h000103; 
10'b0111101111: data <= 24'h0000b8; 
10'b0111110000: data <= 24'h000062; 
10'b0111110001: data <= 24'hffff69; 
10'b0111110010: data <= 24'hfffeb2; 
10'b0111110011: data <= 24'hffff6a; 
10'b0111110100: data <= 24'hffff7d; 
10'b0111110101: data <= 24'hffff99; 
10'b0111110110: data <= 24'hffffc9; 
10'b0111110111: data <= 24'hffffce; 
10'b0111111000: data <= 24'hffffce; 
10'b0111111001: data <= 24'hfffff0; 
10'b0111111010: data <= 24'h00007c; 
10'b0111111011: data <= 24'h000026; 
10'b0111111100: data <= 24'hffff22; 
10'b0111111101: data <= 24'hfffdef; 
10'b0111111110: data <= 24'hfffc96; 
10'b0111111111: data <= 24'hfffbc0; 
10'b1000000000: data <= 24'hfffc0e; 
10'b1000000001: data <= 24'hfffc4e; 
10'b1000000010: data <= 24'hfffb41; 
10'b1000000011: data <= 24'hfffe5e; 
10'b1000000100: data <= 24'hffff82; 
10'b1000000101: data <= 24'h00000f; 
10'b1000000110: data <= 24'h000156; 
10'b1000000111: data <= 24'hfffe97; 
10'b1000001000: data <= 24'hfffe45; 
10'b1000001001: data <= 24'hffff0b; 
10'b1000001010: data <= 24'hfffdd2; 
10'b1000001011: data <= 24'hfffeaa; 
10'b1000001100: data <= 24'hfffdc1; 
10'b1000001101: data <= 24'hfffc8d; 
10'b1000001110: data <= 24'hfffd7a; 
10'b1000001111: data <= 24'hfffe68; 
10'b1000010000: data <= 24'hfffebf; 
10'b1000010001: data <= 24'h000021; 
10'b1000010010: data <= 24'hffffdd; 
10'b1000010011: data <= 24'h000008; 
10'b1000010100: data <= 24'h0000ad; 
10'b1000010101: data <= 24'h0000b9; 
10'b1000010110: data <= 24'h0000aa; 
10'b1000010111: data <= 24'h000055; 
10'b1000011000: data <= 24'hffff6a; 
10'b1000011001: data <= 24'hfffd50; 
10'b1000011010: data <= 24'hfffbb3; 
10'b1000011011: data <= 24'hfffb62; 
10'b1000011100: data <= 24'hfffb43; 
10'b1000011101: data <= 24'hfffb3b; 
10'b1000011110: data <= 24'hfffcc5; 
10'b1000011111: data <= 24'hfffdad; 
10'b1000100000: data <= 24'hfffe9c; 
10'b1000100001: data <= 24'h00009a; 
10'b1000100010: data <= 24'h0001e4; 
10'b1000100011: data <= 24'hfffe07; 
10'b1000100100: data <= 24'hfffe13; 
10'b1000100101: data <= 24'hfffd92; 
10'b1000100110: data <= 24'hfffc23; 
10'b1000100111: data <= 24'hfffc57; 
10'b1000101000: data <= 24'hfffb7f; 
10'b1000101001: data <= 24'hfffbd7; 
10'b1000101010: data <= 24'hfffcd5; 
10'b1000101011: data <= 24'hfffdd2; 
10'b1000101100: data <= 24'hfffee5; 
10'b1000101101: data <= 24'hffff97; 
10'b1000101110: data <= 24'h0000b2; 
10'b1000101111: data <= 24'hffffb0; 
10'b1000110000: data <= 24'hffffa4; 
10'b1000110001: data <= 24'hffffd6; 
10'b1000110010: data <= 24'h000049; 
10'b1000110011: data <= 24'hffffe2; 
10'b1000110100: data <= 24'hffff52; 
10'b1000110101: data <= 24'hfffded; 
10'b1000110110: data <= 24'hfffbaa; 
10'b1000110111: data <= 24'hfffb7b; 
10'b1000111000: data <= 24'hfffbbc; 
10'b1000111001: data <= 24'hfffbd6; 
10'b1000111010: data <= 24'hfffd19; 
10'b1000111011: data <= 24'hfffd01; 
10'b1000111100: data <= 24'h000038; 
10'b1000111101: data <= 24'h00004c; 
10'b1000111110: data <= 24'h000101; 
10'b1000111111: data <= 24'hfffd5b; 
10'b1001000000: data <= 24'hfffcb2; 
10'b1001000001: data <= 24'hfffbaf; 
10'b1001000010: data <= 24'hfffa0b; 
10'b1001000011: data <= 24'hfffc36; 
10'b1001000100: data <= 24'hfffac7; 
10'b1001000101: data <= 24'hfffc05; 
10'b1001000110: data <= 24'hfffd1f; 
10'b1001000111: data <= 24'hfffec6; 
10'b1001001000: data <= 24'hffff2f; 
10'b1001001001: data <= 24'h00009e; 
10'b1001001010: data <= 24'h000096; 
10'b1001001011: data <= 24'h000066; 
10'b1001001100: data <= 24'h00008e; 
10'b1001001101: data <= 24'h000095; 
10'b1001001110: data <= 24'h000021; 
10'b1001001111: data <= 24'hffff3d; 
10'b1001010000: data <= 24'hffff9d; 
10'b1001010001: data <= 24'hfffe27; 
10'b1001010010: data <= 24'hfffdd5; 
10'b1001010011: data <= 24'hfffce1; 
10'b1001010100: data <= 24'hfffd30; 
10'b1001010101: data <= 24'hfffe54; 
10'b1001010110: data <= 24'hfffd9f; 
10'b1001010111: data <= 24'hfffe0f; 
10'b1001011000: data <= 24'hffff22; 
10'b1001011001: data <= 24'h00001e; 
10'b1001011010: data <= 24'hffff7b; 
10'b1001011011: data <= 24'hfffe38; 
10'b1001011100: data <= 24'hfffdf3; 
10'b1001011101: data <= 24'hfffbbe; 
10'b1001011110: data <= 24'hfffbc3; 
10'b1001011111: data <= 24'hfffbc0; 
10'b1001100000: data <= 24'hfffb86; 
10'b1001100001: data <= 24'hfffc36; 
10'b1001100010: data <= 24'hfffdc6; 
10'b1001100011: data <= 24'hfffe51; 
10'b1001100100: data <= 24'hffffed; 
10'b1001100101: data <= 24'h000042; 
10'b1001100110: data <= 24'h000090; 
10'b1001100111: data <= 24'hffffe1; 
10'b1001101000: data <= 24'h000031; 
10'b1001101001: data <= 24'h00000b; 
10'b1001101010: data <= 24'h000026; 
10'b1001101011: data <= 24'hffff88; 
10'b1001101100: data <= 24'hffffc9; 
10'b1001101101: data <= 24'h000046; 
10'b1001101110: data <= 24'hffff53; 
10'b1001101111: data <= 24'h000056; 
10'b1001110000: data <= 24'h000089; 
10'b1001110001: data <= 24'hffff25; 
10'b1001110010: data <= 24'hfffe5f; 
10'b1001110011: data <= 24'hfffd39; 
10'b1001110100: data <= 24'hfffd67; 
10'b1001110101: data <= 24'hfffef4; 
10'b1001110110: data <= 24'h000050; 
10'b1001110111: data <= 24'h00004e; 
10'b1001111000: data <= 24'hfffe63; 
10'b1001111001: data <= 24'hfffe00; 
10'b1001111010: data <= 24'hfffc98; 
10'b1001111011: data <= 24'hfffc98; 
10'b1001111100: data <= 24'hfffc29; 
10'b1001111101: data <= 24'hfffca4; 
10'b1001111110: data <= 24'hfffe4b; 
10'b1001111111: data <= 24'hffff6c; 
10'b1010000000: data <= 24'h00005f; 
10'b1010000001: data <= 24'hffffa3; 
10'b1010000010: data <= 24'h00002d; 
10'b1010000011: data <= 24'h000003; 
10'b1010000100: data <= 24'h000043; 
10'b1010000101: data <= 24'h000088; 
10'b1010000110: data <= 24'hffff97; 
10'b1010000111: data <= 24'hffffa1; 
10'b1010001000: data <= 24'h0000b4; 
10'b1010001001: data <= 24'h0000f1; 
10'b1010001010: data <= 24'h00020d; 
10'b1010001011: data <= 24'h0002bc; 
10'b1010001100: data <= 24'h00014e; 
10'b1010001101: data <= 24'h000043; 
10'b1010001110: data <= 24'hffff32; 
10'b1010001111: data <= 24'hfffe24; 
10'b1010010000: data <= 24'hfffe7b; 
10'b1010010001: data <= 24'h00001b; 
10'b1010010010: data <= 24'h000111; 
10'b1010010011: data <= 24'h0000fb; 
10'b1010010100: data <= 24'hffff97; 
10'b1010010101: data <= 24'hffff65; 
10'b1010010110: data <= 24'hfffdd2; 
10'b1010010111: data <= 24'hfffcf5; 
10'b1010011000: data <= 24'hfffce3; 
10'b1010011001: data <= 24'hfffd92; 
10'b1010011010: data <= 24'hfffdff; 
10'b1010011011: data <= 24'hfffeb1; 
10'b1010011100: data <= 24'hffff6c; 
10'b1010011101: data <= 24'h00000b; 
10'b1010011110: data <= 24'h00000a; 
10'b1010011111: data <= 24'hffffc9; 
10'b1010100000: data <= 24'hffffff; 
10'b1010100001: data <= 24'hffffee; 
10'b1010100010: data <= 24'h000032; 
10'b1010100011: data <= 24'h000075; 
10'b1010100100: data <= 24'h0000fa; 
10'b1010100101: data <= 24'h000240; 
10'b1010100110: data <= 24'h000367; 
10'b1010100111: data <= 24'h0003d6; 
10'b1010101000: data <= 24'h000342; 
10'b1010101001: data <= 24'h0001ae; 
10'b1010101010: data <= 24'h00039f; 
10'b1010101011: data <= 24'h000223; 
10'b1010101100: data <= 24'h0001db; 
10'b1010101101: data <= 24'h00029d; 
10'b1010101110: data <= 24'h00019c; 
10'b1010101111: data <= 24'h000252; 
10'b1010110000: data <= 24'h000160; 
10'b1010110001: data <= 24'h000112; 
10'b1010110010: data <= 24'hffffee; 
10'b1010110011: data <= 24'hffff00; 
10'b1010110100: data <= 24'hfffef0; 
10'b1010110101: data <= 24'hfffeb6; 
10'b1010110110: data <= 24'hfffe8b; 
10'b1010110111: data <= 24'hfffead; 
10'b1010111000: data <= 24'h000034; 
10'b1010111001: data <= 24'hffffe5; 
10'b1010111010: data <= 24'hffffa7; 
10'b1010111011: data <= 24'h000066; 
10'b1010111100: data <= 24'hffffa5; 
10'b1010111101: data <= 24'h000053; 
10'b1010111110: data <= 24'h000096; 
10'b1010111111: data <= 24'h00008d; 
10'b1011000000: data <= 24'h000052; 
10'b1011000001: data <= 24'h00011f; 
10'b1011000010: data <= 24'h0001a9; 
10'b1011000011: data <= 24'h000291; 
10'b1011000100: data <= 24'h0003f7; 
10'b1011000101: data <= 24'h0003df; 
10'b1011000110: data <= 24'h000495; 
10'b1011000111: data <= 24'h000444; 
10'b1011001000: data <= 24'h0003cd; 
10'b1011001001: data <= 24'h000303; 
10'b1011001010: data <= 24'h000313; 
10'b1011001011: data <= 24'h000342; 
10'b1011001100: data <= 24'h0002bb; 
10'b1011001101: data <= 24'h00028d; 
10'b1011001110: data <= 24'h00020f; 
10'b1011001111: data <= 24'h0000b5; 
10'b1011010000: data <= 24'hffff22; 
10'b1011010001: data <= 24'h00001e; 
10'b1011010010: data <= 24'hffff92; 
10'b1011010011: data <= 24'hffffaf; 
10'b1011010100: data <= 24'hffffe6; 
10'b1011010101: data <= 24'h000032; 
10'b1011010110: data <= 24'h0000c7; 
10'b1011010111: data <= 24'h000081; 
10'b1011011000: data <= 24'hffffb9; 
10'b1011011001: data <= 24'h000026; 
10'b1011011010: data <= 24'h0000bc; 
10'b1011011011: data <= 24'hffffe0; 
10'b1011011100: data <= 24'hffffc0; 
10'b1011011101: data <= 24'h0000b0; 
10'b1011011110: data <= 24'h00000d; 
10'b1011011111: data <= 24'h0000a1; 
10'b1011100000: data <= 24'h000099; 
10'b1011100001: data <= 24'h000015; 
10'b1011100010: data <= 24'h0000dd; 
10'b1011100011: data <= 24'h000145; 
10'b1011100100: data <= 24'h00005e; 
10'b1011100101: data <= 24'h000117; 
10'b1011100110: data <= 24'h000257; 
10'b1011100111: data <= 24'h0002e4; 
10'b1011101000: data <= 24'h000247; 
10'b1011101001: data <= 24'h0002ec; 
10'b1011101010: data <= 24'h0001aa; 
10'b1011101011: data <= 24'h0000c9; 
10'b1011101100: data <= 24'h000007; 
10'b1011101101: data <= 24'h00004d; 
10'b1011101110: data <= 24'hffffeb; 
10'b1011101111: data <= 24'h00002b; 
10'b1011110000: data <= 24'h000009; 
10'b1011110001: data <= 24'hffffce; 
10'b1011110010: data <= 24'hfffff4; 
10'b1011110011: data <= 24'hffffe7; 
10'b1011110100: data <= 24'hffffa3; 
10'b1011110101: data <= 24'h00004c; 
10'b1011110110: data <= 24'h000033; 
10'b1011110111: data <= 24'h00005e; 
10'b1011111000: data <= 24'h000080; 
10'b1011111001: data <= 24'h00004d; 
10'b1011111010: data <= 24'h000021; 
10'b1011111011: data <= 24'h00000e; 
10'b1011111100: data <= 24'h0000d2; 
10'b1011111101: data <= 24'h000081; 
10'b1011111110: data <= 24'h000026; 
10'b1011111111: data <= 24'h000082; 
10'b1100000000: data <= 24'h00003f; 
10'b1100000001: data <= 24'h0000f3; 
10'b1100000010: data <= 24'h000091; 
10'b1100000011: data <= 24'h00006f; 
10'b1100000100: data <= 24'h000152; 
10'b1100000101: data <= 24'h000072; 
10'b1100000110: data <= 24'h000065; 
10'b1100000111: data <= 24'h0000eb; 
10'b1100001000: data <= 24'h00001c; 
10'b1100001001: data <= 24'hffffd8; 
10'b1100001010: data <= 24'h0000bf; 
10'b1100001011: data <= 24'h000069; 
10'b1100001100: data <= 24'h000031; 
10'b1100001101: data <= 24'hffffdd; 
10'b1100001110: data <= 24'hffffb2; 
10'b1100001111: data <= 24'h00007f; 
endcase
end

assign dout = data;

endmodule