`timescale 1ns / 1ps 
 
////////////////////////////////////////////////////////////////////////////////// 
// WEIGHT MEMORY (ROM) 
////////////////////////////////////////////////////////////////////////////////// 
module ROM_weights_8 #( 
    parameter int WGHT_INT = 6, // integer part 
    parameter int WGHT_FRC = 16 // fractional part 
)( 
    input logic clk, // clock 
    input logic [9:0] address,
    output [WGHT_INT + WGHT_FRC-1:0] dout 
); 

(* rom_style = "block" *) reg [WGHT_INT + WGHT_FRC-1:0] data;
generate 
  if (WGHT_FRC == 1) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 7'h00; 
        10'b0000000001: data <= 7'h00; 
        10'b0000000010: data <= 7'h00; 
        10'b0000000011: data <= 7'h00; 
        10'b0000000100: data <= 7'h00; 
        10'b0000000101: data <= 7'h00; 
        10'b0000000110: data <= 7'h00; 
        10'b0000000111: data <= 7'h00; 
        10'b0000001000: data <= 7'h00; 
        10'b0000001001: data <= 7'h00; 
        10'b0000001010: data <= 7'h00; 
        10'b0000001011: data <= 7'h00; 
        10'b0000001100: data <= 7'h00; 
        10'b0000001101: data <= 7'h00; 
        10'b0000001110: data <= 7'h00; 
        10'b0000001111: data <= 7'h00; 
        10'b0000010000: data <= 7'h00; 
        10'b0000010001: data <= 7'h00; 
        10'b0000010010: data <= 7'h00; 
        10'b0000010011: data <= 7'h00; 
        10'b0000010100: data <= 7'h00; 
        10'b0000010101: data <= 7'h00; 
        10'b0000010110: data <= 7'h00; 
        10'b0000010111: data <= 7'h00; 
        10'b0000011000: data <= 7'h00; 
        10'b0000011001: data <= 7'h00; 
        10'b0000011010: data <= 7'h00; 
        10'b0000011011: data <= 7'h00; 
        10'b0000011100: data <= 7'h00; 
        10'b0000011101: data <= 7'h00; 
        10'b0000011110: data <= 7'h00; 
        10'b0000011111: data <= 7'h00; 
        10'b0000100000: data <= 7'h00; 
        10'b0000100001: data <= 7'h00; 
        10'b0000100010: data <= 7'h00; 
        10'b0000100011: data <= 7'h00; 
        10'b0000100100: data <= 7'h00; 
        10'b0000100101: data <= 7'h00; 
        10'b0000100110: data <= 7'h00; 
        10'b0000100111: data <= 7'h00; 
        10'b0000101000: data <= 7'h00; 
        10'b0000101001: data <= 7'h00; 
        10'b0000101010: data <= 7'h00; 
        10'b0000101011: data <= 7'h00; 
        10'b0000101100: data <= 7'h00; 
        10'b0000101101: data <= 7'h00; 
        10'b0000101110: data <= 7'h00; 
        10'b0000101111: data <= 7'h00; 
        10'b0000110000: data <= 7'h00; 
        10'b0000110001: data <= 7'h00; 
        10'b0000110010: data <= 7'h00; 
        10'b0000110011: data <= 7'h00; 
        10'b0000110100: data <= 7'h00; 
        10'b0000110101: data <= 7'h00; 
        10'b0000110110: data <= 7'h00; 
        10'b0000110111: data <= 7'h00; 
        10'b0000111000: data <= 7'h00; 
        10'b0000111001: data <= 7'h00; 
        10'b0000111010: data <= 7'h00; 
        10'b0000111011: data <= 7'h00; 
        10'b0000111100: data <= 7'h00; 
        10'b0000111101: data <= 7'h00; 
        10'b0000111110: data <= 7'h00; 
        10'b0000111111: data <= 7'h00; 
        10'b0001000000: data <= 7'h00; 
        10'b0001000001: data <= 7'h00; 
        10'b0001000010: data <= 7'h00; 
        10'b0001000011: data <= 7'h00; 
        10'b0001000100: data <= 7'h00; 
        10'b0001000101: data <= 7'h00; 
        10'b0001000110: data <= 7'h00; 
        10'b0001000111: data <= 7'h00; 
        10'b0001001000: data <= 7'h00; 
        10'b0001001001: data <= 7'h00; 
        10'b0001001010: data <= 7'h00; 
        10'b0001001011: data <= 7'h00; 
        10'b0001001100: data <= 7'h00; 
        10'b0001001101: data <= 7'h00; 
        10'b0001001110: data <= 7'h00; 
        10'b0001001111: data <= 7'h00; 
        10'b0001010000: data <= 7'h00; 
        10'b0001010001: data <= 7'h00; 
        10'b0001010010: data <= 7'h00; 
        10'b0001010011: data <= 7'h00; 
        10'b0001010100: data <= 7'h00; 
        10'b0001010101: data <= 7'h00; 
        10'b0001010110: data <= 7'h00; 
        10'b0001010111: data <= 7'h00; 
        10'b0001011000: data <= 7'h00; 
        10'b0001011001: data <= 7'h00; 
        10'b0001011010: data <= 7'h00; 
        10'b0001011011: data <= 7'h00; 
        10'b0001011100: data <= 7'h00; 
        10'b0001011101: data <= 7'h00; 
        10'b0001011110: data <= 7'h00; 
        10'b0001011111: data <= 7'h00; 
        10'b0001100000: data <= 7'h00; 
        10'b0001100001: data <= 7'h00; 
        10'b0001100010: data <= 7'h00; 
        10'b0001100011: data <= 7'h00; 
        10'b0001100100: data <= 7'h00; 
        10'b0001100101: data <= 7'h00; 
        10'b0001100110: data <= 7'h00; 
        10'b0001100111: data <= 7'h00; 
        10'b0001101000: data <= 7'h00; 
        10'b0001101001: data <= 7'h00; 
        10'b0001101010: data <= 7'h00; 
        10'b0001101011: data <= 7'h00; 
        10'b0001101100: data <= 7'h00; 
        10'b0001101101: data <= 7'h00; 
        10'b0001101110: data <= 7'h00; 
        10'b0001101111: data <= 7'h00; 
        10'b0001110000: data <= 7'h00; 
        10'b0001110001: data <= 7'h00; 
        10'b0001110010: data <= 7'h00; 
        10'b0001110011: data <= 7'h00; 
        10'b0001110100: data <= 7'h00; 
        10'b0001110101: data <= 7'h00; 
        10'b0001110110: data <= 7'h00; 
        10'b0001110111: data <= 7'h00; 
        10'b0001111000: data <= 7'h00; 
        10'b0001111001: data <= 7'h00; 
        10'b0001111010: data <= 7'h00; 
        10'b0001111011: data <= 7'h00; 
        10'b0001111100: data <= 7'h00; 
        10'b0001111101: data <= 7'h00; 
        10'b0001111110: data <= 7'h00; 
        10'b0001111111: data <= 7'h00; 
        10'b0010000000: data <= 7'h00; 
        10'b0010000001: data <= 7'h00; 
        10'b0010000010: data <= 7'h00; 
        10'b0010000011: data <= 7'h00; 
        10'b0010000100: data <= 7'h00; 
        10'b0010000101: data <= 7'h00; 
        10'b0010000110: data <= 7'h00; 
        10'b0010000111: data <= 7'h00; 
        10'b0010001000: data <= 7'h00; 
        10'b0010001001: data <= 7'h00; 
        10'b0010001010: data <= 7'h00; 
        10'b0010001011: data <= 7'h00; 
        10'b0010001100: data <= 7'h00; 
        10'b0010001101: data <= 7'h00; 
        10'b0010001110: data <= 7'h00; 
        10'b0010001111: data <= 7'h00; 
        10'b0010010000: data <= 7'h00; 
        10'b0010010001: data <= 7'h00; 
        10'b0010010010: data <= 7'h00; 
        10'b0010010011: data <= 7'h00; 
        10'b0010010100: data <= 7'h00; 
        10'b0010010101: data <= 7'h00; 
        10'b0010010110: data <= 7'h00; 
        10'b0010010111: data <= 7'h00; 
        10'b0010011000: data <= 7'h00; 
        10'b0010011001: data <= 7'h00; 
        10'b0010011010: data <= 7'h00; 
        10'b0010011011: data <= 7'h00; 
        10'b0010011100: data <= 7'h00; 
        10'b0010011101: data <= 7'h00; 
        10'b0010011110: data <= 7'h00; 
        10'b0010011111: data <= 7'h00; 
        10'b0010100000: data <= 7'h00; 
        10'b0010100001: data <= 7'h00; 
        10'b0010100010: data <= 7'h00; 
        10'b0010100011: data <= 7'h00; 
        10'b0010100100: data <= 7'h00; 
        10'b0010100101: data <= 7'h00; 
        10'b0010100110: data <= 7'h00; 
        10'b0010100111: data <= 7'h00; 
        10'b0010101000: data <= 7'h00; 
        10'b0010101001: data <= 7'h00; 
        10'b0010101010: data <= 7'h00; 
        10'b0010101011: data <= 7'h00; 
        10'b0010101100: data <= 7'h00; 
        10'b0010101101: data <= 7'h00; 
        10'b0010101110: data <= 7'h00; 
        10'b0010101111: data <= 7'h00; 
        10'b0010110000: data <= 7'h00; 
        10'b0010110001: data <= 7'h00; 
        10'b0010110010: data <= 7'h00; 
        10'b0010110011: data <= 7'h00; 
        10'b0010110100: data <= 7'h00; 
        10'b0010110101: data <= 7'h00; 
        10'b0010110110: data <= 7'h00; 
        10'b0010110111: data <= 7'h00; 
        10'b0010111000: data <= 7'h00; 
        10'b0010111001: data <= 7'h00; 
        10'b0010111010: data <= 7'h00; 
        10'b0010111011: data <= 7'h00; 
        10'b0010111100: data <= 7'h00; 
        10'b0010111101: data <= 7'h00; 
        10'b0010111110: data <= 7'h00; 
        10'b0010111111: data <= 7'h00; 
        10'b0011000000: data <= 7'h00; 
        10'b0011000001: data <= 7'h00; 
        10'b0011000010: data <= 7'h00; 
        10'b0011000011: data <= 7'h00; 
        10'b0011000100: data <= 7'h00; 
        10'b0011000101: data <= 7'h00; 
        10'b0011000110: data <= 7'h00; 
        10'b0011000111: data <= 7'h00; 
        10'b0011001000: data <= 7'h00; 
        10'b0011001001: data <= 7'h00; 
        10'b0011001010: data <= 7'h00; 
        10'b0011001011: data <= 7'h00; 
        10'b0011001100: data <= 7'h00; 
        10'b0011001101: data <= 7'h00; 
        10'b0011001110: data <= 7'h00; 
        10'b0011001111: data <= 7'h00; 
        10'b0011010000: data <= 7'h00; 
        10'b0011010001: data <= 7'h00; 
        10'b0011010010: data <= 7'h00; 
        10'b0011010011: data <= 7'h00; 
        10'b0011010100: data <= 7'h00; 
        10'b0011010101: data <= 7'h00; 
        10'b0011010110: data <= 7'h00; 
        10'b0011010111: data <= 7'h00; 
        10'b0011011000: data <= 7'h00; 
        10'b0011011001: data <= 7'h00; 
        10'b0011011010: data <= 7'h00; 
        10'b0011011011: data <= 7'h00; 
        10'b0011011100: data <= 7'h00; 
        10'b0011011101: data <= 7'h00; 
        10'b0011011110: data <= 7'h00; 
        10'b0011011111: data <= 7'h00; 
        10'b0011100000: data <= 7'h00; 
        10'b0011100001: data <= 7'h00; 
        10'b0011100010: data <= 7'h00; 
        10'b0011100011: data <= 7'h00; 
        10'b0011100100: data <= 7'h00; 
        10'b0011100101: data <= 7'h00; 
        10'b0011100110: data <= 7'h00; 
        10'b0011100111: data <= 7'h00; 
        10'b0011101000: data <= 7'h00; 
        10'b0011101001: data <= 7'h00; 
        10'b0011101010: data <= 7'h00; 
        10'b0011101011: data <= 7'h00; 
        10'b0011101100: data <= 7'h00; 
        10'b0011101101: data <= 7'h00; 
        10'b0011101110: data <= 7'h00; 
        10'b0011101111: data <= 7'h00; 
        10'b0011110000: data <= 7'h00; 
        10'b0011110001: data <= 7'h00; 
        10'b0011110010: data <= 7'h00; 
        10'b0011110011: data <= 7'h00; 
        10'b0011110100: data <= 7'h00; 
        10'b0011110101: data <= 7'h00; 
        10'b0011110110: data <= 7'h00; 
        10'b0011110111: data <= 7'h00; 
        10'b0011111000: data <= 7'h00; 
        10'b0011111001: data <= 7'h00; 
        10'b0011111010: data <= 7'h00; 
        10'b0011111011: data <= 7'h00; 
        10'b0011111100: data <= 7'h00; 
        10'b0011111101: data <= 7'h00; 
        10'b0011111110: data <= 7'h00; 
        10'b0011111111: data <= 7'h00; 
        10'b0100000000: data <= 7'h00; 
        10'b0100000001: data <= 7'h00; 
        10'b0100000010: data <= 7'h00; 
        10'b0100000011: data <= 7'h00; 
        10'b0100000100: data <= 7'h00; 
        10'b0100000101: data <= 7'h00; 
        10'b0100000110: data <= 7'h00; 
        10'b0100000111: data <= 7'h00; 
        10'b0100001000: data <= 7'h00; 
        10'b0100001001: data <= 7'h00; 
        10'b0100001010: data <= 7'h00; 
        10'b0100001011: data <= 7'h7f; 
        10'b0100001100: data <= 7'h00; 
        10'b0100001101: data <= 7'h00; 
        10'b0100001110: data <= 7'h00; 
        10'b0100001111: data <= 7'h00; 
        10'b0100010000: data <= 7'h00; 
        10'b0100010001: data <= 7'h00; 
        10'b0100010010: data <= 7'h00; 
        10'b0100010011: data <= 7'h00; 
        10'b0100010100: data <= 7'h00; 
        10'b0100010101: data <= 7'h00; 
        10'b0100010110: data <= 7'h00; 
        10'b0100010111: data <= 7'h00; 
        10'b0100011000: data <= 7'h00; 
        10'b0100011001: data <= 7'h00; 
        10'b0100011010: data <= 7'h00; 
        10'b0100011011: data <= 7'h00; 
        10'b0100011100: data <= 7'h00; 
        10'b0100011101: data <= 7'h00; 
        10'b0100011110: data <= 7'h00; 
        10'b0100011111: data <= 7'h00; 
        10'b0100100000: data <= 7'h00; 
        10'b0100100001: data <= 7'h00; 
        10'b0100100010: data <= 7'h01; 
        10'b0100100011: data <= 7'h00; 
        10'b0100100100: data <= 7'h00; 
        10'b0100100101: data <= 7'h00; 
        10'b0100100110: data <= 7'h00; 
        10'b0100100111: data <= 7'h7f; 
        10'b0100101000: data <= 7'h00; 
        10'b0100101001: data <= 7'h00; 
        10'b0100101010: data <= 7'h00; 
        10'b0100101011: data <= 7'h00; 
        10'b0100101100: data <= 7'h00; 
        10'b0100101101: data <= 7'h00; 
        10'b0100101110: data <= 7'h00; 
        10'b0100101111: data <= 7'h00; 
        10'b0100110000: data <= 7'h00; 
        10'b0100110001: data <= 7'h00; 
        10'b0100110010: data <= 7'h00; 
        10'b0100110011: data <= 7'h00; 
        10'b0100110100: data <= 7'h00; 
        10'b0100110101: data <= 7'h00; 
        10'b0100110110: data <= 7'h00; 
        10'b0100110111: data <= 7'h00; 
        10'b0100111000: data <= 7'h00; 
        10'b0100111001: data <= 7'h00; 
        10'b0100111010: data <= 7'h01; 
        10'b0100111011: data <= 7'h01; 
        10'b0100111100: data <= 7'h01; 
        10'b0100111101: data <= 7'h01; 
        10'b0100111110: data <= 7'h00; 
        10'b0100111111: data <= 7'h00; 
        10'b0101000000: data <= 7'h00; 
        10'b0101000001: data <= 7'h01; 
        10'b0101000010: data <= 7'h01; 
        10'b0101000011: data <= 7'h00; 
        10'b0101000100: data <= 7'h00; 
        10'b0101000101: data <= 7'h00; 
        10'b0101000110: data <= 7'h00; 
        10'b0101000111: data <= 7'h00; 
        10'b0101001000: data <= 7'h00; 
        10'b0101001001: data <= 7'h00; 
        10'b0101001010: data <= 7'h01; 
        10'b0101001011: data <= 7'h01; 
        10'b0101001100: data <= 7'h00; 
        10'b0101001101: data <= 7'h00; 
        10'b0101001110: data <= 7'h00; 
        10'b0101001111: data <= 7'h00; 
        10'b0101010000: data <= 7'h00; 
        10'b0101010001: data <= 7'h00; 
        10'b0101010010: data <= 7'h00; 
        10'b0101010011: data <= 7'h00; 
        10'b0101010100: data <= 7'h00; 
        10'b0101010101: data <= 7'h00; 
        10'b0101010110: data <= 7'h00; 
        10'b0101010111: data <= 7'h00; 
        10'b0101011000: data <= 7'h00; 
        10'b0101011001: data <= 7'h00; 
        10'b0101011010: data <= 7'h00; 
        10'b0101011011: data <= 7'h00; 
        10'b0101011100: data <= 7'h00; 
        10'b0101011101: data <= 7'h01; 
        10'b0101011110: data <= 7'h01; 
        10'b0101011111: data <= 7'h00; 
        10'b0101100000: data <= 7'h00; 
        10'b0101100001: data <= 7'h00; 
        10'b0101100010: data <= 7'h00; 
        10'b0101100011: data <= 7'h00; 
        10'b0101100100: data <= 7'h00; 
        10'b0101100101: data <= 7'h01; 
        10'b0101100110: data <= 7'h01; 
        10'b0101100111: data <= 7'h01; 
        10'b0101101000: data <= 7'h00; 
        10'b0101101001: data <= 7'h00; 
        10'b0101101010: data <= 7'h00; 
        10'b0101101011: data <= 7'h00; 
        10'b0101101100: data <= 7'h00; 
        10'b0101101101: data <= 7'h00; 
        10'b0101101110: data <= 7'h00; 
        10'b0101101111: data <= 7'h00; 
        10'b0101110000: data <= 7'h00; 
        10'b0101110001: data <= 7'h00; 
        10'b0101110010: data <= 7'h00; 
        10'b0101110011: data <= 7'h00; 
        10'b0101110100: data <= 7'h00; 
        10'b0101110101: data <= 7'h00; 
        10'b0101110110: data <= 7'h00; 
        10'b0101110111: data <= 7'h00; 
        10'b0101111000: data <= 7'h00; 
        10'b0101111001: data <= 7'h01; 
        10'b0101111010: data <= 7'h00; 
        10'b0101111011: data <= 7'h01; 
        10'b0101111100: data <= 7'h00; 
        10'b0101111101: data <= 7'h00; 
        10'b0101111110: data <= 7'h00; 
        10'b0101111111: data <= 7'h00; 
        10'b0110000000: data <= 7'h00; 
        10'b0110000001: data <= 7'h00; 
        10'b0110000010: data <= 7'h00; 
        10'b0110000011: data <= 7'h00; 
        10'b0110000100: data <= 7'h00; 
        10'b0110000101: data <= 7'h00; 
        10'b0110000110: data <= 7'h00; 
        10'b0110000111: data <= 7'h00; 
        10'b0110001000: data <= 7'h00; 
        10'b0110001001: data <= 7'h00; 
        10'b0110001010: data <= 7'h00; 
        10'b0110001011: data <= 7'h00; 
        10'b0110001100: data <= 7'h00; 
        10'b0110001101: data <= 7'h00; 
        10'b0110001110: data <= 7'h00; 
        10'b0110001111: data <= 7'h00; 
        10'b0110010000: data <= 7'h7f; 
        10'b0110010001: data <= 7'h00; 
        10'b0110010010: data <= 7'h00; 
        10'b0110010011: data <= 7'h00; 
        10'b0110010100: data <= 7'h00; 
        10'b0110010101: data <= 7'h01; 
        10'b0110010110: data <= 7'h00; 
        10'b0110010111: data <= 7'h00; 
        10'b0110011000: data <= 7'h00; 
        10'b0110011001: data <= 7'h00; 
        10'b0110011010: data <= 7'h00; 
        10'b0110011011: data <= 7'h00; 
        10'b0110011100: data <= 7'h00; 
        10'b0110011101: data <= 7'h00; 
        10'b0110011110: data <= 7'h00; 
        10'b0110011111: data <= 7'h00; 
        10'b0110100000: data <= 7'h00; 
        10'b0110100001: data <= 7'h00; 
        10'b0110100010: data <= 7'h00; 
        10'b0110100011: data <= 7'h00; 
        10'b0110100100: data <= 7'h00; 
        10'b0110100101: data <= 7'h00; 
        10'b0110100110: data <= 7'h00; 
        10'b0110100111: data <= 7'h00; 
        10'b0110101000: data <= 7'h00; 
        10'b0110101001: data <= 7'h00; 
        10'b0110101010: data <= 7'h00; 
        10'b0110101011: data <= 7'h7f; 
        10'b0110101100: data <= 7'h7f; 
        10'b0110101101: data <= 7'h00; 
        10'b0110101110: data <= 7'h00; 
        10'b0110101111: data <= 7'h00; 
        10'b0110110000: data <= 7'h00; 
        10'b0110110001: data <= 7'h00; 
        10'b0110110010: data <= 7'h00; 
        10'b0110110011: data <= 7'h00; 
        10'b0110110100: data <= 7'h00; 
        10'b0110110101: data <= 7'h00; 
        10'b0110110110: data <= 7'h00; 
        10'b0110110111: data <= 7'h00; 
        10'b0110111000: data <= 7'h7f; 
        10'b0110111001: data <= 7'h00; 
        10'b0110111010: data <= 7'h00; 
        10'b0110111011: data <= 7'h00; 
        10'b0110111100: data <= 7'h00; 
        10'b0110111101: data <= 7'h00; 
        10'b0110111110: data <= 7'h00; 
        10'b0110111111: data <= 7'h00; 
        10'b0111000000: data <= 7'h00; 
        10'b0111000001: data <= 7'h00; 
        10'b0111000010: data <= 7'h00; 
        10'b0111000011: data <= 7'h00; 
        10'b0111000100: data <= 7'h00; 
        10'b0111000101: data <= 7'h00; 
        10'b0111000110: data <= 7'h00; 
        10'b0111000111: data <= 7'h00; 
        10'b0111001000: data <= 7'h00; 
        10'b0111001001: data <= 7'h00; 
        10'b0111001010: data <= 7'h00; 
        10'b0111001011: data <= 7'h00; 
        10'b0111001100: data <= 7'h00; 
        10'b0111001101: data <= 7'h00; 
        10'b0111001110: data <= 7'h00; 
        10'b0111001111: data <= 7'h00; 
        10'b0111010000: data <= 7'h00; 
        10'b0111010001: data <= 7'h00; 
        10'b0111010010: data <= 7'h00; 
        10'b0111010011: data <= 7'h00; 
        10'b0111010100: data <= 7'h00; 
        10'b0111010101: data <= 7'h7f; 
        10'b0111010110: data <= 7'h00; 
        10'b0111010111: data <= 7'h00; 
        10'b0111011000: data <= 7'h00; 
        10'b0111011001: data <= 7'h00; 
        10'b0111011010: data <= 7'h00; 
        10'b0111011011: data <= 7'h00; 
        10'b0111011100: data <= 7'h00; 
        10'b0111011101: data <= 7'h00; 
        10'b0111011110: data <= 7'h00; 
        10'b0111011111: data <= 7'h00; 
        10'b0111100000: data <= 7'h00; 
        10'b0111100001: data <= 7'h00; 
        10'b0111100010: data <= 7'h00; 
        10'b0111100011: data <= 7'h00; 
        10'b0111100100: data <= 7'h00; 
        10'b0111100101: data <= 7'h01; 
        10'b0111100110: data <= 7'h00; 
        10'b0111100111: data <= 7'h00; 
        10'b0111101000: data <= 7'h01; 
        10'b0111101001: data <= 7'h00; 
        10'b0111101010: data <= 7'h00; 
        10'b0111101011: data <= 7'h00; 
        10'b0111101100: data <= 7'h00; 
        10'b0111101101: data <= 7'h00; 
        10'b0111101110: data <= 7'h7f; 
        10'b0111101111: data <= 7'h00; 
        10'b0111110000: data <= 7'h00; 
        10'b0111110001: data <= 7'h00; 
        10'b0111110010: data <= 7'h00; 
        10'b0111110011: data <= 7'h00; 
        10'b0111110100: data <= 7'h00; 
        10'b0111110101: data <= 7'h00; 
        10'b0111110110: data <= 7'h00; 
        10'b0111110111: data <= 7'h00; 
        10'b0111111000: data <= 7'h00; 
        10'b0111111001: data <= 7'h00; 
        10'b0111111010: data <= 7'h00; 
        10'b0111111011: data <= 7'h00; 
        10'b0111111100: data <= 7'h00; 
        10'b0111111101: data <= 7'h00; 
        10'b0111111110: data <= 7'h00; 
        10'b0111111111: data <= 7'h00; 
        10'b1000000000: data <= 7'h00; 
        10'b1000000001: data <= 7'h01; 
        10'b1000000010: data <= 7'h00; 
        10'b1000000011: data <= 7'h01; 
        10'b1000000100: data <= 7'h00; 
        10'b1000000101: data <= 7'h00; 
        10'b1000000110: data <= 7'h00; 
        10'b1000000111: data <= 7'h00; 
        10'b1000001000: data <= 7'h00; 
        10'b1000001001: data <= 7'h00; 
        10'b1000001010: data <= 7'h00; 
        10'b1000001011: data <= 7'h00; 
        10'b1000001100: data <= 7'h00; 
        10'b1000001101: data <= 7'h00; 
        10'b1000001110: data <= 7'h00; 
        10'b1000001111: data <= 7'h00; 
        10'b1000010000: data <= 7'h00; 
        10'b1000010001: data <= 7'h00; 
        10'b1000010010: data <= 7'h00; 
        10'b1000010011: data <= 7'h00; 
        10'b1000010100: data <= 7'h00; 
        10'b1000010101: data <= 7'h00; 
        10'b1000010110: data <= 7'h00; 
        10'b1000010111: data <= 7'h00; 
        10'b1000011000: data <= 7'h00; 
        10'b1000011001: data <= 7'h00; 
        10'b1000011010: data <= 7'h00; 
        10'b1000011011: data <= 7'h00; 
        10'b1000011100: data <= 7'h00; 
        10'b1000011101: data <= 7'h00; 
        10'b1000011110: data <= 7'h00; 
        10'b1000011111: data <= 7'h00; 
        10'b1000100000: data <= 7'h00; 
        10'b1000100001: data <= 7'h00; 
        10'b1000100010: data <= 7'h00; 
        10'b1000100011: data <= 7'h00; 
        10'b1000100100: data <= 7'h00; 
        10'b1000100101: data <= 7'h00; 
        10'b1000100110: data <= 7'h00; 
        10'b1000100111: data <= 7'h00; 
        10'b1000101000: data <= 7'h00; 
        10'b1000101001: data <= 7'h00; 
        10'b1000101010: data <= 7'h00; 
        10'b1000101011: data <= 7'h00; 
        10'b1000101100: data <= 7'h00; 
        10'b1000101101: data <= 7'h00; 
        10'b1000101110: data <= 7'h00; 
        10'b1000101111: data <= 7'h00; 
        10'b1000110000: data <= 7'h00; 
        10'b1000110001: data <= 7'h00; 
        10'b1000110010: data <= 7'h00; 
        10'b1000110011: data <= 7'h00; 
        10'b1000110100: data <= 7'h00; 
        10'b1000110101: data <= 7'h00; 
        10'b1000110110: data <= 7'h00; 
        10'b1000110111: data <= 7'h00; 
        10'b1000111000: data <= 7'h00; 
        10'b1000111001: data <= 7'h00; 
        10'b1000111010: data <= 7'h00; 
        10'b1000111011: data <= 7'h00; 
        10'b1000111100: data <= 7'h00; 
        10'b1000111101: data <= 7'h00; 
        10'b1000111110: data <= 7'h00; 
        10'b1000111111: data <= 7'h00; 
        10'b1001000000: data <= 7'h00; 
        10'b1001000001: data <= 7'h00; 
        10'b1001000010: data <= 7'h00; 
        10'b1001000011: data <= 7'h00; 
        10'b1001000100: data <= 7'h00; 
        10'b1001000101: data <= 7'h00; 
        10'b1001000110: data <= 7'h00; 
        10'b1001000111: data <= 7'h00; 
        10'b1001001000: data <= 7'h00; 
        10'b1001001001: data <= 7'h00; 
        10'b1001001010: data <= 7'h00; 
        10'b1001001011: data <= 7'h00; 
        10'b1001001100: data <= 7'h00; 
        10'b1001001101: data <= 7'h00; 
        10'b1001001110: data <= 7'h00; 
        10'b1001001111: data <= 7'h00; 
        10'b1001010000: data <= 7'h00; 
        10'b1001010001: data <= 7'h00; 
        10'b1001010010: data <= 7'h00; 
        10'b1001010011: data <= 7'h00; 
        10'b1001010100: data <= 7'h00; 
        10'b1001010101: data <= 7'h00; 
        10'b1001010110: data <= 7'h00; 
        10'b1001010111: data <= 7'h00; 
        10'b1001011000: data <= 7'h00; 
        10'b1001011001: data <= 7'h00; 
        10'b1001011010: data <= 7'h00; 
        10'b1001011011: data <= 7'h00; 
        10'b1001011100: data <= 7'h00; 
        10'b1001011101: data <= 7'h00; 
        10'b1001011110: data <= 7'h00; 
        10'b1001011111: data <= 7'h00; 
        10'b1001100000: data <= 7'h00; 
        10'b1001100001: data <= 7'h00; 
        10'b1001100010: data <= 7'h00; 
        10'b1001100011: data <= 7'h00; 
        10'b1001100100: data <= 7'h00; 
        10'b1001100101: data <= 7'h00; 
        10'b1001100110: data <= 7'h00; 
        10'b1001100111: data <= 7'h00; 
        10'b1001101000: data <= 7'h00; 
        10'b1001101001: data <= 7'h00; 
        10'b1001101010: data <= 7'h00; 
        10'b1001101011: data <= 7'h00; 
        10'b1001101100: data <= 7'h00; 
        10'b1001101101: data <= 7'h00; 
        10'b1001101110: data <= 7'h00; 
        10'b1001101111: data <= 7'h00; 
        10'b1001110000: data <= 7'h00; 
        10'b1001110001: data <= 7'h00; 
        10'b1001110010: data <= 7'h00; 
        10'b1001110011: data <= 7'h00; 
        10'b1001110100: data <= 7'h00; 
        10'b1001110101: data <= 7'h00; 
        10'b1001110110: data <= 7'h00; 
        10'b1001110111: data <= 7'h00; 
        10'b1001111000: data <= 7'h00; 
        10'b1001111001: data <= 7'h00; 
        10'b1001111010: data <= 7'h00; 
        10'b1001111011: data <= 7'h00; 
        10'b1001111100: data <= 7'h00; 
        10'b1001111101: data <= 7'h00; 
        10'b1001111110: data <= 7'h00; 
        10'b1001111111: data <= 7'h00; 
        10'b1010000000: data <= 7'h00; 
        10'b1010000001: data <= 7'h00; 
        10'b1010000010: data <= 7'h00; 
        10'b1010000011: data <= 7'h00; 
        10'b1010000100: data <= 7'h00; 
        10'b1010000101: data <= 7'h00; 
        10'b1010000110: data <= 7'h00; 
        10'b1010000111: data <= 7'h00; 
        10'b1010001000: data <= 7'h00; 
        10'b1010001001: data <= 7'h7f; 
        10'b1010001010: data <= 7'h00; 
        10'b1010001011: data <= 7'h00; 
        10'b1010001100: data <= 7'h00; 
        10'b1010001101: data <= 7'h00; 
        10'b1010001110: data <= 7'h00; 
        10'b1010001111: data <= 7'h00; 
        10'b1010010000: data <= 7'h00; 
        10'b1010010001: data <= 7'h01; 
        10'b1010010010: data <= 7'h01; 
        10'b1010010011: data <= 7'h00; 
        10'b1010010100: data <= 7'h00; 
        10'b1010010101: data <= 7'h00; 
        10'b1010010110: data <= 7'h00; 
        10'b1010010111: data <= 7'h00; 
        10'b1010011000: data <= 7'h00; 
        10'b1010011001: data <= 7'h00; 
        10'b1010011010: data <= 7'h00; 
        10'b1010011011: data <= 7'h00; 
        10'b1010011100: data <= 7'h00; 
        10'b1010011101: data <= 7'h00; 
        10'b1010011110: data <= 7'h00; 
        10'b1010011111: data <= 7'h00; 
        10'b1010100000: data <= 7'h00; 
        10'b1010100001: data <= 7'h00; 
        10'b1010100010: data <= 7'h00; 
        10'b1010100011: data <= 7'h00; 
        10'b1010100100: data <= 7'h00; 
        10'b1010100101: data <= 7'h00; 
        10'b1010100110: data <= 7'h7f; 
        10'b1010100111: data <= 7'h00; 
        10'b1010101000: data <= 7'h00; 
        10'b1010101001: data <= 7'h00; 
        10'b1010101010: data <= 7'h00; 
        10'b1010101011: data <= 7'h00; 
        10'b1010101100: data <= 7'h00; 
        10'b1010101101: data <= 7'h00; 
        10'b1010101110: data <= 7'h00; 
        10'b1010101111: data <= 7'h01; 
        10'b1010110000: data <= 7'h01; 
        10'b1010110001: data <= 7'h00; 
        10'b1010110010: data <= 7'h01; 
        10'b1010110011: data <= 7'h00; 
        10'b1010110100: data <= 7'h00; 
        10'b1010110101: data <= 7'h00; 
        10'b1010110110: data <= 7'h00; 
        10'b1010110111: data <= 7'h00; 
        10'b1010111000: data <= 7'h00; 
        10'b1010111001: data <= 7'h00; 
        10'b1010111010: data <= 7'h00; 
        10'b1010111011: data <= 7'h00; 
        10'b1010111100: data <= 7'h00; 
        10'b1010111101: data <= 7'h00; 
        10'b1010111110: data <= 7'h00; 
        10'b1010111111: data <= 7'h00; 
        10'b1011000000: data <= 7'h00; 
        10'b1011000001: data <= 7'h00; 
        10'b1011000010: data <= 7'h00; 
        10'b1011000011: data <= 7'h00; 
        10'b1011000100: data <= 7'h00; 
        10'b1011000101: data <= 7'h00; 
        10'b1011000110: data <= 7'h00; 
        10'b1011000111: data <= 7'h00; 
        10'b1011001000: data <= 7'h00; 
        10'b1011001001: data <= 7'h00; 
        10'b1011001010: data <= 7'h00; 
        10'b1011001011: data <= 7'h00; 
        10'b1011001100: data <= 7'h00; 
        10'b1011001101: data <= 7'h00; 
        10'b1011001110: data <= 7'h00; 
        10'b1011001111: data <= 7'h00; 
        10'b1011010000: data <= 7'h00; 
        10'b1011010001: data <= 7'h00; 
        10'b1011010010: data <= 7'h00; 
        10'b1011010011: data <= 7'h00; 
        10'b1011010100: data <= 7'h00; 
        10'b1011010101: data <= 7'h00; 
        10'b1011010110: data <= 7'h00; 
        10'b1011010111: data <= 7'h00; 
        10'b1011011000: data <= 7'h00; 
        10'b1011011001: data <= 7'h00; 
        10'b1011011010: data <= 7'h00; 
        10'b1011011011: data <= 7'h00; 
        10'b1011011100: data <= 7'h00; 
        10'b1011011101: data <= 7'h00; 
        10'b1011011110: data <= 7'h00; 
        10'b1011011111: data <= 7'h00; 
        10'b1011100000: data <= 7'h00; 
        10'b1011100001: data <= 7'h00; 
        10'b1011100010: data <= 7'h00; 
        10'b1011100011: data <= 7'h00; 
        10'b1011100100: data <= 7'h00; 
        10'b1011100101: data <= 7'h00; 
        10'b1011100110: data <= 7'h00; 
        10'b1011100111: data <= 7'h00; 
        10'b1011101000: data <= 7'h00; 
        10'b1011101001: data <= 7'h00; 
        10'b1011101010: data <= 7'h00; 
        10'b1011101011: data <= 7'h00; 
        10'b1011101100: data <= 7'h00; 
        10'b1011101101: data <= 7'h00; 
        10'b1011101110: data <= 7'h00; 
        10'b1011101111: data <= 7'h00; 
        10'b1011110000: data <= 7'h00; 
        10'b1011110001: data <= 7'h00; 
        10'b1011110010: data <= 7'h00; 
        10'b1011110011: data <= 7'h00; 
        10'b1011110100: data <= 7'h00; 
        10'b1011110101: data <= 7'h00; 
        10'b1011110110: data <= 7'h00; 
        10'b1011110111: data <= 7'h00; 
        10'b1011111000: data <= 7'h00; 
        10'b1011111001: data <= 7'h00; 
        10'b1011111010: data <= 7'h00; 
        10'b1011111011: data <= 7'h00; 
        10'b1011111100: data <= 7'h00; 
        10'b1011111101: data <= 7'h00; 
        10'b1011111110: data <= 7'h00; 
        10'b1011111111: data <= 7'h00; 
        10'b1100000000: data <= 7'h00; 
        10'b1100000001: data <= 7'h00; 
        10'b1100000010: data <= 7'h00; 
        10'b1100000011: data <= 7'h00; 
        10'b1100000100: data <= 7'h00; 
        10'b1100000101: data <= 7'h00; 
        10'b1100000110: data <= 7'h00; 
        10'b1100000111: data <= 7'h00; 
        10'b1100001000: data <= 7'h00; 
        10'b1100001001: data <= 7'h00; 
        10'b1100001010: data <= 7'h00; 
        10'b1100001011: data <= 7'h00; 
        10'b1100001100: data <= 7'h00; 
        10'b1100001101: data <= 7'h00; 
        10'b1100001110: data <= 7'h00; 
        10'b1100001111: data <= 7'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 2) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 8'h00; 
        10'b0000000001: data <= 8'h00; 
        10'b0000000010: data <= 8'h00; 
        10'b0000000011: data <= 8'h00; 
        10'b0000000100: data <= 8'h00; 
        10'b0000000101: data <= 8'h00; 
        10'b0000000110: data <= 8'h00; 
        10'b0000000111: data <= 8'h00; 
        10'b0000001000: data <= 8'h00; 
        10'b0000001001: data <= 8'h00; 
        10'b0000001010: data <= 8'h00; 
        10'b0000001011: data <= 8'h00; 
        10'b0000001100: data <= 8'h00; 
        10'b0000001101: data <= 8'h00; 
        10'b0000001110: data <= 8'h00; 
        10'b0000001111: data <= 8'h00; 
        10'b0000010000: data <= 8'h00; 
        10'b0000010001: data <= 8'h00; 
        10'b0000010010: data <= 8'h00; 
        10'b0000010011: data <= 8'h00; 
        10'b0000010100: data <= 8'h00; 
        10'b0000010101: data <= 8'h00; 
        10'b0000010110: data <= 8'h00; 
        10'b0000010111: data <= 8'h00; 
        10'b0000011000: data <= 8'h00; 
        10'b0000011001: data <= 8'h00; 
        10'b0000011010: data <= 8'h00; 
        10'b0000011011: data <= 8'h00; 
        10'b0000011100: data <= 8'h00; 
        10'b0000011101: data <= 8'h00; 
        10'b0000011110: data <= 8'h00; 
        10'b0000011111: data <= 8'h00; 
        10'b0000100000: data <= 8'h00; 
        10'b0000100001: data <= 8'h00; 
        10'b0000100010: data <= 8'h00; 
        10'b0000100011: data <= 8'h00; 
        10'b0000100100: data <= 8'h00; 
        10'b0000100101: data <= 8'h00; 
        10'b0000100110: data <= 8'h00; 
        10'b0000100111: data <= 8'h00; 
        10'b0000101000: data <= 8'h00; 
        10'b0000101001: data <= 8'h00; 
        10'b0000101010: data <= 8'h00; 
        10'b0000101011: data <= 8'h00; 
        10'b0000101100: data <= 8'h00; 
        10'b0000101101: data <= 8'h00; 
        10'b0000101110: data <= 8'h00; 
        10'b0000101111: data <= 8'h00; 
        10'b0000110000: data <= 8'h00; 
        10'b0000110001: data <= 8'h00; 
        10'b0000110010: data <= 8'h00; 
        10'b0000110011: data <= 8'h00; 
        10'b0000110100: data <= 8'h00; 
        10'b0000110101: data <= 8'h00; 
        10'b0000110110: data <= 8'h00; 
        10'b0000110111: data <= 8'h00; 
        10'b0000111000: data <= 8'h00; 
        10'b0000111001: data <= 8'h00; 
        10'b0000111010: data <= 8'h00; 
        10'b0000111011: data <= 8'h00; 
        10'b0000111100: data <= 8'h00; 
        10'b0000111101: data <= 8'h00; 
        10'b0000111110: data <= 8'h00; 
        10'b0000111111: data <= 8'h00; 
        10'b0001000000: data <= 8'h00; 
        10'b0001000001: data <= 8'h00; 
        10'b0001000010: data <= 8'h00; 
        10'b0001000011: data <= 8'h00; 
        10'b0001000100: data <= 8'h00; 
        10'b0001000101: data <= 8'h00; 
        10'b0001000110: data <= 8'h00; 
        10'b0001000111: data <= 8'h00; 
        10'b0001001000: data <= 8'h00; 
        10'b0001001001: data <= 8'h00; 
        10'b0001001010: data <= 8'h00; 
        10'b0001001011: data <= 8'h00; 
        10'b0001001100: data <= 8'h00; 
        10'b0001001101: data <= 8'h00; 
        10'b0001001110: data <= 8'h00; 
        10'b0001001111: data <= 8'h00; 
        10'b0001010000: data <= 8'h00; 
        10'b0001010001: data <= 8'h00; 
        10'b0001010010: data <= 8'h00; 
        10'b0001010011: data <= 8'h00; 
        10'b0001010100: data <= 8'h00; 
        10'b0001010101: data <= 8'h00; 
        10'b0001010110: data <= 8'h00; 
        10'b0001010111: data <= 8'h00; 
        10'b0001011000: data <= 8'h00; 
        10'b0001011001: data <= 8'h00; 
        10'b0001011010: data <= 8'h00; 
        10'b0001011011: data <= 8'h00; 
        10'b0001011100: data <= 8'h00; 
        10'b0001011101: data <= 8'h00; 
        10'b0001011110: data <= 8'h00; 
        10'b0001011111: data <= 8'h00; 
        10'b0001100000: data <= 8'h00; 
        10'b0001100001: data <= 8'h00; 
        10'b0001100010: data <= 8'h00; 
        10'b0001100011: data <= 8'h00; 
        10'b0001100100: data <= 8'h00; 
        10'b0001100101: data <= 8'h00; 
        10'b0001100110: data <= 8'h00; 
        10'b0001100111: data <= 8'h00; 
        10'b0001101000: data <= 8'h00; 
        10'b0001101001: data <= 8'h00; 
        10'b0001101010: data <= 8'h00; 
        10'b0001101011: data <= 8'h00; 
        10'b0001101100: data <= 8'h00; 
        10'b0001101101: data <= 8'h00; 
        10'b0001101110: data <= 8'h00; 
        10'b0001101111: data <= 8'h00; 
        10'b0001110000: data <= 8'h00; 
        10'b0001110001: data <= 8'h00; 
        10'b0001110010: data <= 8'h00; 
        10'b0001110011: data <= 8'h00; 
        10'b0001110100: data <= 8'h00; 
        10'b0001110101: data <= 8'h00; 
        10'b0001110110: data <= 8'h00; 
        10'b0001110111: data <= 8'h00; 
        10'b0001111000: data <= 8'h00; 
        10'b0001111001: data <= 8'h00; 
        10'b0001111010: data <= 8'h00; 
        10'b0001111011: data <= 8'h00; 
        10'b0001111100: data <= 8'h00; 
        10'b0001111101: data <= 8'h00; 
        10'b0001111110: data <= 8'h01; 
        10'b0001111111: data <= 8'h01; 
        10'b0010000000: data <= 8'h00; 
        10'b0010000001: data <= 8'h00; 
        10'b0010000010: data <= 8'h00; 
        10'b0010000011: data <= 8'h00; 
        10'b0010000100: data <= 8'h00; 
        10'b0010000101: data <= 8'h00; 
        10'b0010000110: data <= 8'h00; 
        10'b0010000111: data <= 8'h00; 
        10'b0010001000: data <= 8'h00; 
        10'b0010001001: data <= 8'h00; 
        10'b0010001010: data <= 8'h00; 
        10'b0010001011: data <= 8'h00; 
        10'b0010001100: data <= 8'h00; 
        10'b0010001101: data <= 8'h00; 
        10'b0010001110: data <= 8'h00; 
        10'b0010001111: data <= 8'h00; 
        10'b0010010000: data <= 8'h00; 
        10'b0010010001: data <= 8'h00; 
        10'b0010010010: data <= 8'h00; 
        10'b0010010011: data <= 8'h00; 
        10'b0010010100: data <= 8'h00; 
        10'b0010010101: data <= 8'h00; 
        10'b0010010110: data <= 8'h00; 
        10'b0010010111: data <= 8'h00; 
        10'b0010011000: data <= 8'h01; 
        10'b0010011001: data <= 8'h01; 
        10'b0010011010: data <= 8'h01; 
        10'b0010011011: data <= 8'h00; 
        10'b0010011100: data <= 8'h00; 
        10'b0010011101: data <= 8'h01; 
        10'b0010011110: data <= 8'h00; 
        10'b0010011111: data <= 8'h00; 
        10'b0010100000: data <= 8'h00; 
        10'b0010100001: data <= 8'h00; 
        10'b0010100010: data <= 8'h00; 
        10'b0010100011: data <= 8'h00; 
        10'b0010100100: data <= 8'h00; 
        10'b0010100101: data <= 8'h00; 
        10'b0010100110: data <= 8'h00; 
        10'b0010100111: data <= 8'h00; 
        10'b0010101000: data <= 8'h00; 
        10'b0010101001: data <= 8'h00; 
        10'b0010101010: data <= 8'h00; 
        10'b0010101011: data <= 8'h00; 
        10'b0010101100: data <= 8'h00; 
        10'b0010101101: data <= 8'h00; 
        10'b0010101110: data <= 8'h00; 
        10'b0010101111: data <= 8'h00; 
        10'b0010110000: data <= 8'h00; 
        10'b0010110001: data <= 8'h00; 
        10'b0010110010: data <= 8'h00; 
        10'b0010110011: data <= 8'h00; 
        10'b0010110100: data <= 8'h00; 
        10'b0010110101: data <= 8'h00; 
        10'b0010110110: data <= 8'h00; 
        10'b0010110111: data <= 8'h01; 
        10'b0010111000: data <= 8'h00; 
        10'b0010111001: data <= 8'h00; 
        10'b0010111010: data <= 8'h00; 
        10'b0010111011: data <= 8'h00; 
        10'b0010111100: data <= 8'h00; 
        10'b0010111101: data <= 8'h00; 
        10'b0010111110: data <= 8'h00; 
        10'b0010111111: data <= 8'h00; 
        10'b0011000000: data <= 8'h00; 
        10'b0011000001: data <= 8'h00; 
        10'b0011000010: data <= 8'h00; 
        10'b0011000011: data <= 8'h00; 
        10'b0011000100: data <= 8'h00; 
        10'b0011000101: data <= 8'h00; 
        10'b0011000110: data <= 8'h00; 
        10'b0011000111: data <= 8'h00; 
        10'b0011001000: data <= 8'h00; 
        10'b0011001001: data <= 8'h00; 
        10'b0011001010: data <= 8'h00; 
        10'b0011001011: data <= 8'h00; 
        10'b0011001100: data <= 8'h00; 
        10'b0011001101: data <= 8'h00; 
        10'b0011001110: data <= 8'h00; 
        10'b0011001111: data <= 8'h00; 
        10'b0011010000: data <= 8'h00; 
        10'b0011010001: data <= 8'h00; 
        10'b0011010010: data <= 8'h00; 
        10'b0011010011: data <= 8'h00; 
        10'b0011010100: data <= 8'h00; 
        10'b0011010101: data <= 8'h00; 
        10'b0011010110: data <= 8'h00; 
        10'b0011010111: data <= 8'h00; 
        10'b0011011000: data <= 8'h00; 
        10'b0011011001: data <= 8'h00; 
        10'b0011011010: data <= 8'h00; 
        10'b0011011011: data <= 8'h01; 
        10'b0011011100: data <= 8'h01; 
        10'b0011011101: data <= 8'h00; 
        10'b0011011110: data <= 8'h00; 
        10'b0011011111: data <= 8'h00; 
        10'b0011100000: data <= 8'h00; 
        10'b0011100001: data <= 8'h00; 
        10'b0011100010: data <= 8'h00; 
        10'b0011100011: data <= 8'h00; 
        10'b0011100100: data <= 8'h00; 
        10'b0011100101: data <= 8'h00; 
        10'b0011100110: data <= 8'h00; 
        10'b0011100111: data <= 8'h00; 
        10'b0011101000: data <= 8'h00; 
        10'b0011101001: data <= 8'h01; 
        10'b0011101010: data <= 8'h00; 
        10'b0011101011: data <= 8'h00; 
        10'b0011101100: data <= 8'h00; 
        10'b0011101101: data <= 8'h01; 
        10'b0011101110: data <= 8'h00; 
        10'b0011101111: data <= 8'h00; 
        10'b0011110000: data <= 8'h00; 
        10'b0011110001: data <= 8'h00; 
        10'b0011110010: data <= 8'h00; 
        10'b0011110011: data <= 8'h00; 
        10'b0011110100: data <= 8'h00; 
        10'b0011110101: data <= 8'h01; 
        10'b0011110110: data <= 8'h00; 
        10'b0011110111: data <= 8'h01; 
        10'b0011111000: data <= 8'h01; 
        10'b0011111001: data <= 8'h00; 
        10'b0011111010: data <= 8'h00; 
        10'b0011111011: data <= 8'h00; 
        10'b0011111100: data <= 8'h00; 
        10'b0011111101: data <= 8'h00; 
        10'b0011111110: data <= 8'h00; 
        10'b0011111111: data <= 8'h00; 
        10'b0100000000: data <= 8'h00; 
        10'b0100000001: data <= 8'h00; 
        10'b0100000010: data <= 8'h00; 
        10'b0100000011: data <= 8'h01; 
        10'b0100000100: data <= 8'h01; 
        10'b0100000101: data <= 8'h01; 
        10'b0100000110: data <= 8'h00; 
        10'b0100000111: data <= 8'h01; 
        10'b0100001000: data <= 8'h00; 
        10'b0100001001: data <= 8'h00; 
        10'b0100001010: data <= 8'hff; 
        10'b0100001011: data <= 8'hff; 
        10'b0100001100: data <= 8'h00; 
        10'b0100001101: data <= 8'h00; 
        10'b0100001110: data <= 8'h00; 
        10'b0100001111: data <= 8'h00; 
        10'b0100010000: data <= 8'h00; 
        10'b0100010001: data <= 8'h00; 
        10'b0100010010: data <= 8'h01; 
        10'b0100010011: data <= 8'h01; 
        10'b0100010100: data <= 8'h00; 
        10'b0100010101: data <= 8'h00; 
        10'b0100010110: data <= 8'h00; 
        10'b0100010111: data <= 8'h00; 
        10'b0100011000: data <= 8'h00; 
        10'b0100011001: data <= 8'h00; 
        10'b0100011010: data <= 8'h00; 
        10'b0100011011: data <= 8'h00; 
        10'b0100011100: data <= 8'h00; 
        10'b0100011101: data <= 8'h00; 
        10'b0100011110: data <= 8'h00; 
        10'b0100011111: data <= 8'h01; 
        10'b0100100000: data <= 8'h01; 
        10'b0100100001: data <= 8'h01; 
        10'b0100100010: data <= 8'h01; 
        10'b0100100011: data <= 8'h01; 
        10'b0100100100: data <= 8'h01; 
        10'b0100100101: data <= 8'h00; 
        10'b0100100110: data <= 8'h00; 
        10'b0100100111: data <= 8'hff; 
        10'b0100101000: data <= 8'hff; 
        10'b0100101001: data <= 8'h00; 
        10'b0100101010: data <= 8'h00; 
        10'b0100101011: data <= 8'h00; 
        10'b0100101100: data <= 8'h00; 
        10'b0100101101: data <= 8'h01; 
        10'b0100101110: data <= 8'h01; 
        10'b0100101111: data <= 8'h01; 
        10'b0100110000: data <= 8'h00; 
        10'b0100110001: data <= 8'h00; 
        10'b0100110010: data <= 8'h00; 
        10'b0100110011: data <= 8'h00; 
        10'b0100110100: data <= 8'h00; 
        10'b0100110101: data <= 8'h00; 
        10'b0100110110: data <= 8'h00; 
        10'b0100110111: data <= 8'h00; 
        10'b0100111000: data <= 8'h00; 
        10'b0100111001: data <= 8'h01; 
        10'b0100111010: data <= 8'h01; 
        10'b0100111011: data <= 8'h01; 
        10'b0100111100: data <= 8'h01; 
        10'b0100111101: data <= 8'h01; 
        10'b0100111110: data <= 8'h01; 
        10'b0100111111: data <= 8'h00; 
        10'b0101000000: data <= 8'h01; 
        10'b0101000001: data <= 8'h01; 
        10'b0101000010: data <= 8'h02; 
        10'b0101000011: data <= 8'h00; 
        10'b0101000100: data <= 8'hff; 
        10'b0101000101: data <= 8'h00; 
        10'b0101000110: data <= 8'h00; 
        10'b0101000111: data <= 8'h00; 
        10'b0101001000: data <= 8'h01; 
        10'b0101001001: data <= 8'h01; 
        10'b0101001010: data <= 8'h01; 
        10'b0101001011: data <= 8'h01; 
        10'b0101001100: data <= 8'h01; 
        10'b0101001101: data <= 8'h00; 
        10'b0101001110: data <= 8'h00; 
        10'b0101001111: data <= 8'h00; 
        10'b0101010000: data <= 8'h00; 
        10'b0101010001: data <= 8'h00; 
        10'b0101010010: data <= 8'h00; 
        10'b0101010011: data <= 8'h00; 
        10'b0101010100: data <= 8'h00; 
        10'b0101010101: data <= 8'h01; 
        10'b0101010110: data <= 8'h01; 
        10'b0101010111: data <= 8'h01; 
        10'b0101011000: data <= 8'h01; 
        10'b0101011001: data <= 8'h01; 
        10'b0101011010: data <= 8'h00; 
        10'b0101011011: data <= 8'h00; 
        10'b0101011100: data <= 8'h00; 
        10'b0101011101: data <= 8'h02; 
        10'b0101011110: data <= 8'h02; 
        10'b0101011111: data <= 8'h00; 
        10'b0101100000: data <= 8'h00; 
        10'b0101100001: data <= 8'h00; 
        10'b0101100010: data <= 8'h00; 
        10'b0101100011: data <= 8'h00; 
        10'b0101100100: data <= 8'h01; 
        10'b0101100101: data <= 8'h01; 
        10'b0101100110: data <= 8'h01; 
        10'b0101100111: data <= 8'h01; 
        10'b0101101000: data <= 8'h01; 
        10'b0101101001: data <= 8'h00; 
        10'b0101101010: data <= 8'h00; 
        10'b0101101011: data <= 8'h00; 
        10'b0101101100: data <= 8'h00; 
        10'b0101101101: data <= 8'h00; 
        10'b0101101110: data <= 8'h00; 
        10'b0101101111: data <= 8'h00; 
        10'b0101110000: data <= 8'h00; 
        10'b0101110001: data <= 8'h00; 
        10'b0101110010: data <= 8'h00; 
        10'b0101110011: data <= 8'h00; 
        10'b0101110100: data <= 8'h00; 
        10'b0101110101: data <= 8'h00; 
        10'b0101110110: data <= 8'h00; 
        10'b0101110111: data <= 8'h00; 
        10'b0101111000: data <= 8'h01; 
        10'b0101111001: data <= 8'h01; 
        10'b0101111010: data <= 8'h00; 
        10'b0101111011: data <= 8'h01; 
        10'b0101111100: data <= 8'h00; 
        10'b0101111101: data <= 8'h00; 
        10'b0101111110: data <= 8'h00; 
        10'b0101111111: data <= 8'h00; 
        10'b0110000000: data <= 8'h00; 
        10'b0110000001: data <= 8'h00; 
        10'b0110000010: data <= 8'h00; 
        10'b0110000011: data <= 8'h00; 
        10'b0110000100: data <= 8'h00; 
        10'b0110000101: data <= 8'h00; 
        10'b0110000110: data <= 8'h00; 
        10'b0110000111: data <= 8'h00; 
        10'b0110001000: data <= 8'h00; 
        10'b0110001001: data <= 8'h00; 
        10'b0110001010: data <= 8'h00; 
        10'b0110001011: data <= 8'h00; 
        10'b0110001100: data <= 8'h00; 
        10'b0110001101: data <= 8'h00; 
        10'b0110001110: data <= 8'hff; 
        10'b0110001111: data <= 8'hff; 
        10'b0110010000: data <= 8'hff; 
        10'b0110010001: data <= 8'hff; 
        10'b0110010010: data <= 8'h00; 
        10'b0110010011: data <= 8'h01; 
        10'b0110010100: data <= 8'h01; 
        10'b0110010101: data <= 8'h01; 
        10'b0110010110: data <= 8'h01; 
        10'b0110010111: data <= 8'h01; 
        10'b0110011000: data <= 8'h00; 
        10'b0110011001: data <= 8'h00; 
        10'b0110011010: data <= 8'h00; 
        10'b0110011011: data <= 8'h00; 
        10'b0110011100: data <= 8'hff; 
        10'b0110011101: data <= 8'hff; 
        10'b0110011110: data <= 8'h00; 
        10'b0110011111: data <= 8'hff; 
        10'b0110100000: data <= 8'h00; 
        10'b0110100001: data <= 8'h00; 
        10'b0110100010: data <= 8'h00; 
        10'b0110100011: data <= 8'h00; 
        10'b0110100100: data <= 8'h00; 
        10'b0110100101: data <= 8'h00; 
        10'b0110100110: data <= 8'h00; 
        10'b0110100111: data <= 8'h00; 
        10'b0110101000: data <= 8'h00; 
        10'b0110101001: data <= 8'h00; 
        10'b0110101010: data <= 8'hff; 
        10'b0110101011: data <= 8'hff; 
        10'b0110101100: data <= 8'hff; 
        10'b0110101101: data <= 8'h00; 
        10'b0110101110: data <= 8'h00; 
        10'b0110101111: data <= 8'h00; 
        10'b0110110000: data <= 8'h01; 
        10'b0110110001: data <= 8'h01; 
        10'b0110110010: data <= 8'h01; 
        10'b0110110011: data <= 8'h00; 
        10'b0110110100: data <= 8'h00; 
        10'b0110110101: data <= 8'h00; 
        10'b0110110110: data <= 8'h00; 
        10'b0110110111: data <= 8'hff; 
        10'b0110111000: data <= 8'hff; 
        10'b0110111001: data <= 8'hff; 
        10'b0110111010: data <= 8'hff; 
        10'b0110111011: data <= 8'h00; 
        10'b0110111100: data <= 8'h00; 
        10'b0110111101: data <= 8'h00; 
        10'b0110111110: data <= 8'h00; 
        10'b0110111111: data <= 8'h00; 
        10'b0111000000: data <= 8'h00; 
        10'b0111000001: data <= 8'h00; 
        10'b0111000010: data <= 8'h00; 
        10'b0111000011: data <= 8'h00; 
        10'b0111000100: data <= 8'h00; 
        10'b0111000101: data <= 8'hff; 
        10'b0111000110: data <= 8'hff; 
        10'b0111000111: data <= 8'hff; 
        10'b0111001000: data <= 8'h00; 
        10'b0111001001: data <= 8'h00; 
        10'b0111001010: data <= 8'h00; 
        10'b0111001011: data <= 8'h00; 
        10'b0111001100: data <= 8'h01; 
        10'b0111001101: data <= 8'h01; 
        10'b0111001110: data <= 8'h00; 
        10'b0111001111: data <= 8'h00; 
        10'b0111010000: data <= 8'h00; 
        10'b0111010001: data <= 8'h00; 
        10'b0111010010: data <= 8'hff; 
        10'b0111010011: data <= 8'hff; 
        10'b0111010100: data <= 8'hff; 
        10'b0111010101: data <= 8'hff; 
        10'b0111010110: data <= 8'hff; 
        10'b0111010111: data <= 8'h00; 
        10'b0111011000: data <= 8'h00; 
        10'b0111011001: data <= 8'h00; 
        10'b0111011010: data <= 8'h00; 
        10'b0111011011: data <= 8'h00; 
        10'b0111011100: data <= 8'h00; 
        10'b0111011101: data <= 8'h00; 
        10'b0111011110: data <= 8'h00; 
        10'b0111011111: data <= 8'h00; 
        10'b0111100000: data <= 8'h00; 
        10'b0111100001: data <= 8'hff; 
        10'b0111100010: data <= 8'hff; 
        10'b0111100011: data <= 8'h00; 
        10'b0111100100: data <= 8'h01; 
        10'b0111100101: data <= 8'h01; 
        10'b0111100110: data <= 8'h00; 
        10'b0111100111: data <= 8'h01; 
        10'b0111101000: data <= 8'h01; 
        10'b0111101001: data <= 8'h01; 
        10'b0111101010: data <= 8'h00; 
        10'b0111101011: data <= 8'h00; 
        10'b0111101100: data <= 8'h00; 
        10'b0111101101: data <= 8'h00; 
        10'b0111101110: data <= 8'hff; 
        10'b0111101111: data <= 8'h00; 
        10'b0111110000: data <= 8'h00; 
        10'b0111110001: data <= 8'hff; 
        10'b0111110010: data <= 8'hff; 
        10'b0111110011: data <= 8'h00; 
        10'b0111110100: data <= 8'h00; 
        10'b0111110101: data <= 8'h00; 
        10'b0111110110: data <= 8'h00; 
        10'b0111110111: data <= 8'h00; 
        10'b0111111000: data <= 8'h00; 
        10'b0111111001: data <= 8'h00; 
        10'b0111111010: data <= 8'h00; 
        10'b0111111011: data <= 8'h00; 
        10'b0111111100: data <= 8'h00; 
        10'b0111111101: data <= 8'h00; 
        10'b0111111110: data <= 8'h00; 
        10'b0111111111: data <= 8'h00; 
        10'b1000000000: data <= 8'h01; 
        10'b1000000001: data <= 8'h01; 
        10'b1000000010: data <= 8'h01; 
        10'b1000000011: data <= 8'h01; 
        10'b1000000100: data <= 8'h01; 
        10'b1000000101: data <= 8'h00; 
        10'b1000000110: data <= 8'hff; 
        10'b1000000111: data <= 8'h00; 
        10'b1000001000: data <= 8'h00; 
        10'b1000001001: data <= 8'hff; 
        10'b1000001010: data <= 8'h00; 
        10'b1000001011: data <= 8'h00; 
        10'b1000001100: data <= 8'h00; 
        10'b1000001101: data <= 8'h00; 
        10'b1000001110: data <= 8'h00; 
        10'b1000001111: data <= 8'h00; 
        10'b1000010000: data <= 8'h00; 
        10'b1000010001: data <= 8'h00; 
        10'b1000010010: data <= 8'h00; 
        10'b1000010011: data <= 8'h00; 
        10'b1000010100: data <= 8'h00; 
        10'b1000010101: data <= 8'h00; 
        10'b1000010110: data <= 8'h00; 
        10'b1000010111: data <= 8'h00; 
        10'b1000011000: data <= 8'h00; 
        10'b1000011001: data <= 8'h00; 
        10'b1000011010: data <= 8'h00; 
        10'b1000011011: data <= 8'h00; 
        10'b1000011100: data <= 8'h00; 
        10'b1000011101: data <= 8'h01; 
        10'b1000011110: data <= 8'h00; 
        10'b1000011111: data <= 8'h00; 
        10'b1000100000: data <= 8'h00; 
        10'b1000100001: data <= 8'hff; 
        10'b1000100010: data <= 8'hff; 
        10'b1000100011: data <= 8'h00; 
        10'b1000100100: data <= 8'h00; 
        10'b1000100101: data <= 8'h00; 
        10'b1000100110: data <= 8'h00; 
        10'b1000100111: data <= 8'h00; 
        10'b1000101000: data <= 8'h00; 
        10'b1000101001: data <= 8'h00; 
        10'b1000101010: data <= 8'h00; 
        10'b1000101011: data <= 8'h00; 
        10'b1000101100: data <= 8'h00; 
        10'b1000101101: data <= 8'h00; 
        10'b1000101110: data <= 8'h00; 
        10'b1000101111: data <= 8'h00; 
        10'b1000110000: data <= 8'h00; 
        10'b1000110001: data <= 8'h00; 
        10'b1000110010: data <= 8'h00; 
        10'b1000110011: data <= 8'h00; 
        10'b1000110100: data <= 8'h00; 
        10'b1000110101: data <= 8'h00; 
        10'b1000110110: data <= 8'h00; 
        10'b1000110111: data <= 8'h01; 
        10'b1000111000: data <= 8'h00; 
        10'b1000111001: data <= 8'h00; 
        10'b1000111010: data <= 8'h00; 
        10'b1000111011: data <= 8'hff; 
        10'b1000111100: data <= 8'h00; 
        10'b1000111101: data <= 8'h00; 
        10'b1000111110: data <= 8'hff; 
        10'b1000111111: data <= 8'h00; 
        10'b1001000000: data <= 8'hff; 
        10'b1001000001: data <= 8'h00; 
        10'b1001000010: data <= 8'h00; 
        10'b1001000011: data <= 8'h00; 
        10'b1001000100: data <= 8'h00; 
        10'b1001000101: data <= 8'h00; 
        10'b1001000110: data <= 8'h00; 
        10'b1001000111: data <= 8'h00; 
        10'b1001001000: data <= 8'h00; 
        10'b1001001001: data <= 8'h00; 
        10'b1001001010: data <= 8'h00; 
        10'b1001001011: data <= 8'h00; 
        10'b1001001100: data <= 8'h00; 
        10'b1001001101: data <= 8'h00; 
        10'b1001001110: data <= 8'h00; 
        10'b1001001111: data <= 8'h00; 
        10'b1001010000: data <= 8'hff; 
        10'b1001010001: data <= 8'h00; 
        10'b1001010010: data <= 8'h00; 
        10'b1001010011: data <= 8'h01; 
        10'b1001010100: data <= 8'h00; 
        10'b1001010101: data <= 8'h00; 
        10'b1001010110: data <= 8'h00; 
        10'b1001010111: data <= 8'h00; 
        10'b1001011000: data <= 8'h00; 
        10'b1001011001: data <= 8'h00; 
        10'b1001011010: data <= 8'h00; 
        10'b1001011011: data <= 8'h00; 
        10'b1001011100: data <= 8'hff; 
        10'b1001011101: data <= 8'h00; 
        10'b1001011110: data <= 8'h00; 
        10'b1001011111: data <= 8'h00; 
        10'b1001100000: data <= 8'h00; 
        10'b1001100001: data <= 8'h00; 
        10'b1001100010: data <= 8'h00; 
        10'b1001100011: data <= 8'h00; 
        10'b1001100100: data <= 8'h00; 
        10'b1001100101: data <= 8'h00; 
        10'b1001100110: data <= 8'h00; 
        10'b1001100111: data <= 8'h00; 
        10'b1001101000: data <= 8'h00; 
        10'b1001101001: data <= 8'h00; 
        10'b1001101010: data <= 8'h00; 
        10'b1001101011: data <= 8'h00; 
        10'b1001101100: data <= 8'h00; 
        10'b1001101101: data <= 8'hff; 
        10'b1001101110: data <= 8'h00; 
        10'b1001101111: data <= 8'h00; 
        10'b1001110000: data <= 8'h00; 
        10'b1001110001: data <= 8'h00; 
        10'b1001110010: data <= 8'h00; 
        10'b1001110011: data <= 8'h00; 
        10'b1001110100: data <= 8'h01; 
        10'b1001110101: data <= 8'h01; 
        10'b1001110110: data <= 8'h01; 
        10'b1001110111: data <= 8'h00; 
        10'b1001111000: data <= 8'h00; 
        10'b1001111001: data <= 8'h00; 
        10'b1001111010: data <= 8'h00; 
        10'b1001111011: data <= 8'h00; 
        10'b1001111100: data <= 8'h00; 
        10'b1001111101: data <= 8'h00; 
        10'b1001111110: data <= 8'h00; 
        10'b1001111111: data <= 8'h00; 
        10'b1010000000: data <= 8'h00; 
        10'b1010000001: data <= 8'h00; 
        10'b1010000010: data <= 8'h00; 
        10'b1010000011: data <= 8'h00; 
        10'b1010000100: data <= 8'h00; 
        10'b1010000101: data <= 8'h00; 
        10'b1010000110: data <= 8'h00; 
        10'b1010000111: data <= 8'h00; 
        10'b1010001000: data <= 8'h00; 
        10'b1010001001: data <= 8'hff; 
        10'b1010001010: data <= 8'hff; 
        10'b1010001011: data <= 8'h00; 
        10'b1010001100: data <= 8'h00; 
        10'b1010001101: data <= 8'h00; 
        10'b1010001110: data <= 8'h00; 
        10'b1010001111: data <= 8'h00; 
        10'b1010010000: data <= 8'h01; 
        10'b1010010001: data <= 8'h01; 
        10'b1010010010: data <= 8'h01; 
        10'b1010010011: data <= 8'h01; 
        10'b1010010100: data <= 8'h01; 
        10'b1010010101: data <= 8'h01; 
        10'b1010010110: data <= 8'h00; 
        10'b1010010111: data <= 8'h01; 
        10'b1010011000: data <= 8'h00; 
        10'b1010011001: data <= 8'h00; 
        10'b1010011010: data <= 8'h00; 
        10'b1010011011: data <= 8'h00; 
        10'b1010011100: data <= 8'h00; 
        10'b1010011101: data <= 8'h00; 
        10'b1010011110: data <= 8'h00; 
        10'b1010011111: data <= 8'h00; 
        10'b1010100000: data <= 8'h00; 
        10'b1010100001: data <= 8'h00; 
        10'b1010100010: data <= 8'h00; 
        10'b1010100011: data <= 8'h00; 
        10'b1010100100: data <= 8'h00; 
        10'b1010100101: data <= 8'hff; 
        10'b1010100110: data <= 8'hff; 
        10'b1010100111: data <= 8'hff; 
        10'b1010101000: data <= 8'h00; 
        10'b1010101001: data <= 8'h00; 
        10'b1010101010: data <= 8'h00; 
        10'b1010101011: data <= 8'h00; 
        10'b1010101100: data <= 8'h00; 
        10'b1010101101: data <= 8'h00; 
        10'b1010101110: data <= 8'h00; 
        10'b1010101111: data <= 8'h01; 
        10'b1010110000: data <= 8'h01; 
        10'b1010110001: data <= 8'h01; 
        10'b1010110010: data <= 8'h01; 
        10'b1010110011: data <= 8'h01; 
        10'b1010110100: data <= 8'h00; 
        10'b1010110101: data <= 8'h00; 
        10'b1010110110: data <= 8'h00; 
        10'b1010110111: data <= 8'h00; 
        10'b1010111000: data <= 8'h00; 
        10'b1010111001: data <= 8'h00; 
        10'b1010111010: data <= 8'h00; 
        10'b1010111011: data <= 8'h00; 
        10'b1010111100: data <= 8'h00; 
        10'b1010111101: data <= 8'h00; 
        10'b1010111110: data <= 8'h00; 
        10'b1010111111: data <= 8'h00; 
        10'b1011000000: data <= 8'h00; 
        10'b1011000001: data <= 8'h00; 
        10'b1011000010: data <= 8'h00; 
        10'b1011000011: data <= 8'h00; 
        10'b1011000100: data <= 8'hff; 
        10'b1011000101: data <= 8'hff; 
        10'b1011000110: data <= 8'h00; 
        10'b1011000111: data <= 8'h00; 
        10'b1011001000: data <= 8'h00; 
        10'b1011001001: data <= 8'h00; 
        10'b1011001010: data <= 8'h00; 
        10'b1011001011: data <= 8'h00; 
        10'b1011001100: data <= 8'h00; 
        10'b1011001101: data <= 8'h00; 
        10'b1011001110: data <= 8'h00; 
        10'b1011001111: data <= 8'h00; 
        10'b1011010000: data <= 8'h00; 
        10'b1011010001: data <= 8'h00; 
        10'b1011010010: data <= 8'h00; 
        10'b1011010011: data <= 8'h00; 
        10'b1011010100: data <= 8'h00; 
        10'b1011010101: data <= 8'h00; 
        10'b1011010110: data <= 8'h00; 
        10'b1011010111: data <= 8'h00; 
        10'b1011011000: data <= 8'h00; 
        10'b1011011001: data <= 8'h00; 
        10'b1011011010: data <= 8'h00; 
        10'b1011011011: data <= 8'h00; 
        10'b1011011100: data <= 8'h00; 
        10'b1011011101: data <= 8'h00; 
        10'b1011011110: data <= 8'h00; 
        10'b1011011111: data <= 8'h00; 
        10'b1011100000: data <= 8'h00; 
        10'b1011100001: data <= 8'h00; 
        10'b1011100010: data <= 8'h00; 
        10'b1011100011: data <= 8'h00; 
        10'b1011100100: data <= 8'h00; 
        10'b1011100101: data <= 8'h00; 
        10'b1011100110: data <= 8'h00; 
        10'b1011100111: data <= 8'h00; 
        10'b1011101000: data <= 8'h00; 
        10'b1011101001: data <= 8'h00; 
        10'b1011101010: data <= 8'h00; 
        10'b1011101011: data <= 8'h00; 
        10'b1011101100: data <= 8'h00; 
        10'b1011101101: data <= 8'h00; 
        10'b1011101110: data <= 8'h00; 
        10'b1011101111: data <= 8'h00; 
        10'b1011110000: data <= 8'h00; 
        10'b1011110001: data <= 8'h00; 
        10'b1011110010: data <= 8'h00; 
        10'b1011110011: data <= 8'h00; 
        10'b1011110100: data <= 8'h00; 
        10'b1011110101: data <= 8'h00; 
        10'b1011110110: data <= 8'h00; 
        10'b1011110111: data <= 8'h00; 
        10'b1011111000: data <= 8'h00; 
        10'b1011111001: data <= 8'h00; 
        10'b1011111010: data <= 8'h00; 
        10'b1011111011: data <= 8'h00; 
        10'b1011111100: data <= 8'h00; 
        10'b1011111101: data <= 8'h00; 
        10'b1011111110: data <= 8'h00; 
        10'b1011111111: data <= 8'h00; 
        10'b1100000000: data <= 8'h00; 
        10'b1100000001: data <= 8'h00; 
        10'b1100000010: data <= 8'h00; 
        10'b1100000011: data <= 8'h00; 
        10'b1100000100: data <= 8'h00; 
        10'b1100000101: data <= 8'h00; 
        10'b1100000110: data <= 8'h00; 
        10'b1100000111: data <= 8'h00; 
        10'b1100001000: data <= 8'h00; 
        10'b1100001001: data <= 8'h00; 
        10'b1100001010: data <= 8'h00; 
        10'b1100001011: data <= 8'h00; 
        10'b1100001100: data <= 8'h00; 
        10'b1100001101: data <= 8'h00; 
        10'b1100001110: data <= 8'h00; 
        10'b1100001111: data <= 8'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 3) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 9'h000; 
        10'b0000000001: data <= 9'h000; 
        10'b0000000010: data <= 9'h000; 
        10'b0000000011: data <= 9'h000; 
        10'b0000000100: data <= 9'h000; 
        10'b0000000101: data <= 9'h000; 
        10'b0000000110: data <= 9'h000; 
        10'b0000000111: data <= 9'h000; 
        10'b0000001000: data <= 9'h000; 
        10'b0000001001: data <= 9'h000; 
        10'b0000001010: data <= 9'h000; 
        10'b0000001011: data <= 9'h000; 
        10'b0000001100: data <= 9'h000; 
        10'b0000001101: data <= 9'h000; 
        10'b0000001110: data <= 9'h000; 
        10'b0000001111: data <= 9'h000; 
        10'b0000010000: data <= 9'h000; 
        10'b0000010001: data <= 9'h000; 
        10'b0000010010: data <= 9'h000; 
        10'b0000010011: data <= 9'h000; 
        10'b0000010100: data <= 9'h000; 
        10'b0000010101: data <= 9'h000; 
        10'b0000010110: data <= 9'h000; 
        10'b0000010111: data <= 9'h000; 
        10'b0000011000: data <= 9'h000; 
        10'b0000011001: data <= 9'h000; 
        10'b0000011010: data <= 9'h000; 
        10'b0000011011: data <= 9'h000; 
        10'b0000011100: data <= 9'h000; 
        10'b0000011101: data <= 9'h000; 
        10'b0000011110: data <= 9'h000; 
        10'b0000011111: data <= 9'h000; 
        10'b0000100000: data <= 9'h000; 
        10'b0000100001: data <= 9'h000; 
        10'b0000100010: data <= 9'h000; 
        10'b0000100011: data <= 9'h000; 
        10'b0000100100: data <= 9'h000; 
        10'b0000100101: data <= 9'h000; 
        10'b0000100110: data <= 9'h000; 
        10'b0000100111: data <= 9'h000; 
        10'b0000101000: data <= 9'h000; 
        10'b0000101001: data <= 9'h000; 
        10'b0000101010: data <= 9'h000; 
        10'b0000101011: data <= 9'h000; 
        10'b0000101100: data <= 9'h000; 
        10'b0000101101: data <= 9'h000; 
        10'b0000101110: data <= 9'h000; 
        10'b0000101111: data <= 9'h000; 
        10'b0000110000: data <= 9'h000; 
        10'b0000110001: data <= 9'h000; 
        10'b0000110010: data <= 9'h000; 
        10'b0000110011: data <= 9'h000; 
        10'b0000110100: data <= 9'h000; 
        10'b0000110101: data <= 9'h000; 
        10'b0000110110: data <= 9'h000; 
        10'b0000110111: data <= 9'h000; 
        10'b0000111000: data <= 9'h000; 
        10'b0000111001: data <= 9'h000; 
        10'b0000111010: data <= 9'h000; 
        10'b0000111011: data <= 9'h000; 
        10'b0000111100: data <= 9'h000; 
        10'b0000111101: data <= 9'h000; 
        10'b0000111110: data <= 9'h000; 
        10'b0000111111: data <= 9'h000; 
        10'b0001000000: data <= 9'h000; 
        10'b0001000001: data <= 9'h000; 
        10'b0001000010: data <= 9'h000; 
        10'b0001000011: data <= 9'h000; 
        10'b0001000100: data <= 9'h000; 
        10'b0001000101: data <= 9'h000; 
        10'b0001000110: data <= 9'h000; 
        10'b0001000111: data <= 9'h000; 
        10'b0001001000: data <= 9'h1ff; 
        10'b0001001001: data <= 9'h000; 
        10'b0001001010: data <= 9'h000; 
        10'b0001001011: data <= 9'h000; 
        10'b0001001100: data <= 9'h000; 
        10'b0001001101: data <= 9'h000; 
        10'b0001001110: data <= 9'h000; 
        10'b0001001111: data <= 9'h000; 
        10'b0001010000: data <= 9'h000; 
        10'b0001010001: data <= 9'h000; 
        10'b0001010010: data <= 9'h000; 
        10'b0001010011: data <= 9'h000; 
        10'b0001010100: data <= 9'h000; 
        10'b0001010101: data <= 9'h000; 
        10'b0001010110: data <= 9'h000; 
        10'b0001010111: data <= 9'h000; 
        10'b0001011000: data <= 9'h000; 
        10'b0001011001: data <= 9'h000; 
        10'b0001011010: data <= 9'h000; 
        10'b0001011011: data <= 9'h000; 
        10'b0001011100: data <= 9'h000; 
        10'b0001011101: data <= 9'h000; 
        10'b0001011110: data <= 9'h000; 
        10'b0001011111: data <= 9'h1ff; 
        10'b0001100000: data <= 9'h1ff; 
        10'b0001100001: data <= 9'h1ff; 
        10'b0001100010: data <= 9'h1ff; 
        10'b0001100011: data <= 9'h000; 
        10'b0001100100: data <= 9'h1ff; 
        10'b0001100101: data <= 9'h1ff; 
        10'b0001100110: data <= 9'h000; 
        10'b0001100111: data <= 9'h000; 
        10'b0001101000: data <= 9'h1ff; 
        10'b0001101001: data <= 9'h000; 
        10'b0001101010: data <= 9'h000; 
        10'b0001101011: data <= 9'h000; 
        10'b0001101100: data <= 9'h000; 
        10'b0001101101: data <= 9'h000; 
        10'b0001101110: data <= 9'h000; 
        10'b0001101111: data <= 9'h000; 
        10'b0001110000: data <= 9'h000; 
        10'b0001110001: data <= 9'h000; 
        10'b0001110010: data <= 9'h000; 
        10'b0001110011: data <= 9'h000; 
        10'b0001110100: data <= 9'h000; 
        10'b0001110101: data <= 9'h000; 
        10'b0001110110: data <= 9'h000; 
        10'b0001110111: data <= 9'h000; 
        10'b0001111000: data <= 9'h000; 
        10'b0001111001: data <= 9'h000; 
        10'b0001111010: data <= 9'h000; 
        10'b0001111011: data <= 9'h000; 
        10'b0001111100: data <= 9'h001; 
        10'b0001111101: data <= 9'h000; 
        10'b0001111110: data <= 9'h001; 
        10'b0001111111: data <= 9'h001; 
        10'b0010000000: data <= 9'h000; 
        10'b0010000001: data <= 9'h000; 
        10'b0010000010: data <= 9'h000; 
        10'b0010000011: data <= 9'h000; 
        10'b0010000100: data <= 9'h000; 
        10'b0010000101: data <= 9'h000; 
        10'b0010000110: data <= 9'h1ff; 
        10'b0010000111: data <= 9'h000; 
        10'b0010001000: data <= 9'h000; 
        10'b0010001001: data <= 9'h000; 
        10'b0010001010: data <= 9'h000; 
        10'b0010001011: data <= 9'h000; 
        10'b0010001100: data <= 9'h000; 
        10'b0010001101: data <= 9'h000; 
        10'b0010001110: data <= 9'h000; 
        10'b0010001111: data <= 9'h000; 
        10'b0010010000: data <= 9'h000; 
        10'b0010010001: data <= 9'h000; 
        10'b0010010010: data <= 9'h000; 
        10'b0010010011: data <= 9'h1ff; 
        10'b0010010100: data <= 9'h000; 
        10'b0010010101: data <= 9'h000; 
        10'b0010010110: data <= 9'h1ff; 
        10'b0010010111: data <= 9'h001; 
        10'b0010011000: data <= 9'h002; 
        10'b0010011001: data <= 9'h001; 
        10'b0010011010: data <= 9'h002; 
        10'b0010011011: data <= 9'h001; 
        10'b0010011100: data <= 9'h001; 
        10'b0010011101: data <= 9'h001; 
        10'b0010011110: data <= 9'h000; 
        10'b0010011111: data <= 9'h000; 
        10'b0010100000: data <= 9'h000; 
        10'b0010100001: data <= 9'h000; 
        10'b0010100010: data <= 9'h1ff; 
        10'b0010100011: data <= 9'h1ff; 
        10'b0010100100: data <= 9'h000; 
        10'b0010100101: data <= 9'h000; 
        10'b0010100110: data <= 9'h000; 
        10'b0010100111: data <= 9'h000; 
        10'b0010101000: data <= 9'h000; 
        10'b0010101001: data <= 9'h000; 
        10'b0010101010: data <= 9'h000; 
        10'b0010101011: data <= 9'h000; 
        10'b0010101100: data <= 9'h1ff; 
        10'b0010101101: data <= 9'h000; 
        10'b0010101110: data <= 9'h1ff; 
        10'b0010101111: data <= 9'h1ff; 
        10'b0010110000: data <= 9'h000; 
        10'b0010110001: data <= 9'h000; 
        10'b0010110010: data <= 9'h000; 
        10'b0010110011: data <= 9'h000; 
        10'b0010110100: data <= 9'h001; 
        10'b0010110101: data <= 9'h001; 
        10'b0010110110: data <= 9'h001; 
        10'b0010110111: data <= 9'h001; 
        10'b0010111000: data <= 9'h001; 
        10'b0010111001: data <= 9'h001; 
        10'b0010111010: data <= 9'h000; 
        10'b0010111011: data <= 9'h001; 
        10'b0010111100: data <= 9'h000; 
        10'b0010111101: data <= 9'h000; 
        10'b0010111110: data <= 9'h001; 
        10'b0010111111: data <= 9'h001; 
        10'b0011000000: data <= 9'h000; 
        10'b0011000001: data <= 9'h000; 
        10'b0011000010: data <= 9'h000; 
        10'b0011000011: data <= 9'h000; 
        10'b0011000100: data <= 9'h000; 
        10'b0011000101: data <= 9'h000; 
        10'b0011000110: data <= 9'h000; 
        10'b0011000111: data <= 9'h000; 
        10'b0011001000: data <= 9'h1ff; 
        10'b0011001001: data <= 9'h000; 
        10'b0011001010: data <= 9'h1ff; 
        10'b0011001011: data <= 9'h000; 
        10'b0011001100: data <= 9'h001; 
        10'b0011001101: data <= 9'h000; 
        10'b0011001110: data <= 9'h000; 
        10'b0011001111: data <= 9'h000; 
        10'b0011010000: data <= 9'h1ff; 
        10'b0011010001: data <= 9'h1ff; 
        10'b0011010010: data <= 9'h1ff; 
        10'b0011010011: data <= 9'h000; 
        10'b0011010100: data <= 9'h001; 
        10'b0011010101: data <= 9'h000; 
        10'b0011010110: data <= 9'h000; 
        10'b0011010111: data <= 9'h000; 
        10'b0011011000: data <= 9'h001; 
        10'b0011011001: data <= 9'h001; 
        10'b0011011010: data <= 9'h000; 
        10'b0011011011: data <= 9'h002; 
        10'b0011011100: data <= 9'h001; 
        10'b0011011101: data <= 9'h000; 
        10'b0011011110: data <= 9'h000; 
        10'b0011011111: data <= 9'h000; 
        10'b0011100000: data <= 9'h000; 
        10'b0011100001: data <= 9'h000; 
        10'b0011100010: data <= 9'h000; 
        10'b0011100011: data <= 9'h000; 
        10'b0011100100: data <= 9'h000; 
        10'b0011100101: data <= 9'h000; 
        10'b0011100110: data <= 9'h001; 
        10'b0011100111: data <= 9'h000; 
        10'b0011101000: data <= 9'h000; 
        10'b0011101001: data <= 9'h001; 
        10'b0011101010: data <= 9'h000; 
        10'b0011101011: data <= 9'h000; 
        10'b0011101100: data <= 9'h001; 
        10'b0011101101: data <= 9'h001; 
        10'b0011101110: data <= 9'h1ff; 
        10'b0011101111: data <= 9'h1ff; 
        10'b0011110000: data <= 9'h001; 
        10'b0011110001: data <= 9'h000; 
        10'b0011110010: data <= 9'h000; 
        10'b0011110011: data <= 9'h001; 
        10'b0011110100: data <= 9'h000; 
        10'b0011110101: data <= 9'h001; 
        10'b0011110110: data <= 9'h001; 
        10'b0011110111: data <= 9'h001; 
        10'b0011111000: data <= 9'h001; 
        10'b0011111001: data <= 9'h000; 
        10'b0011111010: data <= 9'h000; 
        10'b0011111011: data <= 9'h000; 
        10'b0011111100: data <= 9'h000; 
        10'b0011111101: data <= 9'h000; 
        10'b0011111110: data <= 9'h000; 
        10'b0011111111: data <= 9'h000; 
        10'b0100000000: data <= 9'h000; 
        10'b0100000001: data <= 9'h001; 
        10'b0100000010: data <= 9'h001; 
        10'b0100000011: data <= 9'h001; 
        10'b0100000100: data <= 9'h002; 
        10'b0100000101: data <= 9'h001; 
        10'b0100000110: data <= 9'h001; 
        10'b0100000111: data <= 9'h002; 
        10'b0100001000: data <= 9'h000; 
        10'b0100001001: data <= 9'h000; 
        10'b0100001010: data <= 9'h1fe; 
        10'b0100001011: data <= 9'h1fe; 
        10'b0100001100: data <= 9'h1ff; 
        10'b0100001101: data <= 9'h000; 
        10'b0100001110: data <= 9'h000; 
        10'b0100001111: data <= 9'h000; 
        10'b0100010000: data <= 9'h001; 
        10'b0100010001: data <= 9'h001; 
        10'b0100010010: data <= 9'h001; 
        10'b0100010011: data <= 9'h001; 
        10'b0100010100: data <= 9'h000; 
        10'b0100010101: data <= 9'h000; 
        10'b0100010110: data <= 9'h000; 
        10'b0100010111: data <= 9'h000; 
        10'b0100011000: data <= 9'h000; 
        10'b0100011001: data <= 9'h000; 
        10'b0100011010: data <= 9'h000; 
        10'b0100011011: data <= 9'h000; 
        10'b0100011100: data <= 9'h000; 
        10'b0100011101: data <= 9'h001; 
        10'b0100011110: data <= 9'h001; 
        10'b0100011111: data <= 9'h002; 
        10'b0100100000: data <= 9'h001; 
        10'b0100100001: data <= 9'h002; 
        10'b0100100010: data <= 9'h002; 
        10'b0100100011: data <= 9'h001; 
        10'b0100100100: data <= 9'h001; 
        10'b0100100101: data <= 9'h001; 
        10'b0100100110: data <= 9'h000; 
        10'b0100100111: data <= 9'h1fe; 
        10'b0100101000: data <= 9'h1fe; 
        10'b0100101001: data <= 9'h1ff; 
        10'b0100101010: data <= 9'h001; 
        10'b0100101011: data <= 9'h001; 
        10'b0100101100: data <= 9'h001; 
        10'b0100101101: data <= 9'h002; 
        10'b0100101110: data <= 9'h002; 
        10'b0100101111: data <= 9'h001; 
        10'b0100110000: data <= 9'h000; 
        10'b0100110001: data <= 9'h000; 
        10'b0100110010: data <= 9'h000; 
        10'b0100110011: data <= 9'h000; 
        10'b0100110100: data <= 9'h000; 
        10'b0100110101: data <= 9'h000; 
        10'b0100110110: data <= 9'h000; 
        10'b0100110111: data <= 9'h1ff; 
        10'b0100111000: data <= 9'h000; 
        10'b0100111001: data <= 9'h001; 
        10'b0100111010: data <= 9'h002; 
        10'b0100111011: data <= 9'h003; 
        10'b0100111100: data <= 9'h002; 
        10'b0100111101: data <= 9'h003; 
        10'b0100111110: data <= 9'h002; 
        10'b0100111111: data <= 9'h001; 
        10'b0101000000: data <= 9'h001; 
        10'b0101000001: data <= 9'h003; 
        10'b0101000010: data <= 9'h003; 
        10'b0101000011: data <= 9'h000; 
        10'b0101000100: data <= 9'h1fe; 
        10'b0101000101: data <= 9'h1ff; 
        10'b0101000110: data <= 9'h1ff; 
        10'b0101000111: data <= 9'h000; 
        10'b0101001000: data <= 9'h001; 
        10'b0101001001: data <= 9'h002; 
        10'b0101001010: data <= 9'h002; 
        10'b0101001011: data <= 9'h002; 
        10'b0101001100: data <= 9'h002; 
        10'b0101001101: data <= 9'h000; 
        10'b0101001110: data <= 9'h000; 
        10'b0101001111: data <= 9'h000; 
        10'b0101010000: data <= 9'h000; 
        10'b0101010001: data <= 9'h000; 
        10'b0101010010: data <= 9'h000; 
        10'b0101010011: data <= 9'h000; 
        10'b0101010100: data <= 9'h000; 
        10'b0101010101: data <= 9'h001; 
        10'b0101010110: data <= 9'h001; 
        10'b0101010111: data <= 9'h002; 
        10'b0101011000: data <= 9'h002; 
        10'b0101011001: data <= 9'h002; 
        10'b0101011010: data <= 9'h000; 
        10'b0101011011: data <= 9'h000; 
        10'b0101011100: data <= 9'h000; 
        10'b0101011101: data <= 9'h003; 
        10'b0101011110: data <= 9'h003; 
        10'b0101011111: data <= 9'h001; 
        10'b0101100000: data <= 9'h000; 
        10'b0101100001: data <= 9'h000; 
        10'b0101100010: data <= 9'h000; 
        10'b0101100011: data <= 9'h001; 
        10'b0101100100: data <= 9'h001; 
        10'b0101100101: data <= 9'h002; 
        10'b0101100110: data <= 9'h003; 
        10'b0101100111: data <= 9'h002; 
        10'b0101101000: data <= 9'h001; 
        10'b0101101001: data <= 9'h001; 
        10'b0101101010: data <= 9'h000; 
        10'b0101101011: data <= 9'h000; 
        10'b0101101100: data <= 9'h000; 
        10'b0101101101: data <= 9'h000; 
        10'b0101101110: data <= 9'h000; 
        10'b0101101111: data <= 9'h000; 
        10'b0101110000: data <= 9'h000; 
        10'b0101110001: data <= 9'h000; 
        10'b0101110010: data <= 9'h000; 
        10'b0101110011: data <= 9'h000; 
        10'b0101110100: data <= 9'h000; 
        10'b0101110101: data <= 9'h000; 
        10'b0101110110: data <= 9'h1ff; 
        10'b0101110111: data <= 9'h000; 
        10'b0101111000: data <= 9'h001; 
        10'b0101111001: data <= 9'h003; 
        10'b0101111010: data <= 9'h001; 
        10'b0101111011: data <= 9'h002; 
        10'b0101111100: data <= 9'h001; 
        10'b0101111101: data <= 9'h1ff; 
        10'b0101111110: data <= 9'h000; 
        10'b0101111111: data <= 9'h000; 
        10'b0110000000: data <= 9'h001; 
        10'b0110000001: data <= 9'h001; 
        10'b0110000010: data <= 9'h000; 
        10'b0110000011: data <= 9'h001; 
        10'b0110000100: data <= 9'h000; 
        10'b0110000101: data <= 9'h000; 
        10'b0110000110: data <= 9'h000; 
        10'b0110000111: data <= 9'h000; 
        10'b0110001000: data <= 9'h000; 
        10'b0110001001: data <= 9'h000; 
        10'b0110001010: data <= 9'h000; 
        10'b0110001011: data <= 9'h000; 
        10'b0110001100: data <= 9'h000; 
        10'b0110001101: data <= 9'h1ff; 
        10'b0110001110: data <= 9'h1fe; 
        10'b0110001111: data <= 9'h1fe; 
        10'b0110010000: data <= 9'h1fe; 
        10'b0110010001: data <= 9'h1fe; 
        10'b0110010010: data <= 9'h000; 
        10'b0110010011: data <= 9'h001; 
        10'b0110010100: data <= 9'h001; 
        10'b0110010101: data <= 9'h002; 
        10'b0110010110: data <= 9'h002; 
        10'b0110010111: data <= 9'h001; 
        10'b0110011000: data <= 9'h000; 
        10'b0110011001: data <= 9'h000; 
        10'b0110011010: data <= 9'h000; 
        10'b0110011011: data <= 9'h1ff; 
        10'b0110011100: data <= 9'h1ff; 
        10'b0110011101: data <= 9'h1ff; 
        10'b0110011110: data <= 9'h1ff; 
        10'b0110011111: data <= 9'h1ff; 
        10'b0110100000: data <= 9'h1ff; 
        10'b0110100001: data <= 9'h000; 
        10'b0110100010: data <= 9'h000; 
        10'b0110100011: data <= 9'h000; 
        10'b0110100100: data <= 9'h000; 
        10'b0110100101: data <= 9'h000; 
        10'b0110100110: data <= 9'h000; 
        10'b0110100111: data <= 9'h000; 
        10'b0110101000: data <= 9'h000; 
        10'b0110101001: data <= 9'h1ff; 
        10'b0110101010: data <= 9'h1fe; 
        10'b0110101011: data <= 9'h1fe; 
        10'b0110101100: data <= 9'h1fe; 
        10'b0110101101: data <= 9'h1ff; 
        10'b0110101110: data <= 9'h000; 
        10'b0110101111: data <= 9'h000; 
        10'b0110110000: data <= 9'h002; 
        10'b0110110001: data <= 9'h002; 
        10'b0110110010: data <= 9'h002; 
        10'b0110110011: data <= 9'h001; 
        10'b0110110100: data <= 9'h000; 
        10'b0110110101: data <= 9'h000; 
        10'b0110110110: data <= 9'h000; 
        10'b0110110111: data <= 9'h1fe; 
        10'b0110111000: data <= 9'h1fe; 
        10'b0110111001: data <= 9'h1fe; 
        10'b0110111010: data <= 9'h1ff; 
        10'b0110111011: data <= 9'h1ff; 
        10'b0110111100: data <= 9'h1ff; 
        10'b0110111101: data <= 9'h000; 
        10'b0110111110: data <= 9'h1ff; 
        10'b0110111111: data <= 9'h000; 
        10'b0111000000: data <= 9'h000; 
        10'b0111000001: data <= 9'h000; 
        10'b0111000010: data <= 9'h000; 
        10'b0111000011: data <= 9'h000; 
        10'b0111000100: data <= 9'h1ff; 
        10'b0111000101: data <= 9'h1ff; 
        10'b0111000110: data <= 9'h1fe; 
        10'b0111000111: data <= 9'h1ff; 
        10'b0111001000: data <= 9'h001; 
        10'b0111001001: data <= 9'h001; 
        10'b0111001010: data <= 9'h000; 
        10'b0111001011: data <= 9'h001; 
        10'b0111001100: data <= 9'h002; 
        10'b0111001101: data <= 9'h001; 
        10'b0111001110: data <= 9'h001; 
        10'b0111001111: data <= 9'h001; 
        10'b0111010000: data <= 9'h000; 
        10'b0111010001: data <= 9'h1ff; 
        10'b0111010010: data <= 9'h1ff; 
        10'b0111010011: data <= 9'h1fe; 
        10'b0111010100: data <= 9'h1fe; 
        10'b0111010101: data <= 9'h1fe; 
        10'b0111010110: data <= 9'h1fe; 
        10'b0111010111: data <= 9'h1ff; 
        10'b0111011000: data <= 9'h1ff; 
        10'b0111011001: data <= 9'h000; 
        10'b0111011010: data <= 9'h000; 
        10'b0111011011: data <= 9'h000; 
        10'b0111011100: data <= 9'h000; 
        10'b0111011101: data <= 9'h000; 
        10'b0111011110: data <= 9'h000; 
        10'b0111011111: data <= 9'h000; 
        10'b0111100000: data <= 9'h000; 
        10'b0111100001: data <= 9'h1ff; 
        10'b0111100010: data <= 9'h1fe; 
        10'b0111100011: data <= 9'h000; 
        10'b0111100100: data <= 9'h002; 
        10'b0111100101: data <= 9'h002; 
        10'b0111100110: data <= 9'h001; 
        10'b0111100111: data <= 9'h002; 
        10'b0111101000: data <= 9'h002; 
        10'b0111101001: data <= 9'h002; 
        10'b0111101010: data <= 9'h000; 
        10'b0111101011: data <= 9'h000; 
        10'b0111101100: data <= 9'h000; 
        10'b0111101101: data <= 9'h1ff; 
        10'b0111101110: data <= 9'h1fe; 
        10'b0111101111: data <= 9'h1ff; 
        10'b0111110000: data <= 9'h1ff; 
        10'b0111110001: data <= 9'h1ff; 
        10'b0111110010: data <= 9'h1ff; 
        10'b0111110011: data <= 9'h1ff; 
        10'b0111110100: data <= 9'h000; 
        10'b0111110101: data <= 9'h1ff; 
        10'b0111110110: data <= 9'h000; 
        10'b0111110111: data <= 9'h000; 
        10'b0111111000: data <= 9'h000; 
        10'b0111111001: data <= 9'h000; 
        10'b0111111010: data <= 9'h000; 
        10'b0111111011: data <= 9'h1ff; 
        10'b0111111100: data <= 9'h1ff; 
        10'b0111111101: data <= 9'h1ff; 
        10'b0111111110: data <= 9'h000; 
        10'b0111111111: data <= 9'h000; 
        10'b1000000000: data <= 9'h001; 
        10'b1000000001: data <= 9'h002; 
        10'b1000000010: data <= 9'h002; 
        10'b1000000011: data <= 9'h002; 
        10'b1000000100: data <= 9'h001; 
        10'b1000000101: data <= 9'h001; 
        10'b1000000110: data <= 9'h1ff; 
        10'b1000000111: data <= 9'h000; 
        10'b1000001000: data <= 9'h1ff; 
        10'b1000001001: data <= 9'h1fe; 
        10'b1000001010: data <= 9'h000; 
        10'b1000001011: data <= 9'h000; 
        10'b1000001100: data <= 9'h000; 
        10'b1000001101: data <= 9'h1ff; 
        10'b1000001110: data <= 9'h000; 
        10'b1000001111: data <= 9'h1ff; 
        10'b1000010000: data <= 9'h1ff; 
        10'b1000010001: data <= 9'h1ff; 
        10'b1000010010: data <= 9'h000; 
        10'b1000010011: data <= 9'h000; 
        10'b1000010100: data <= 9'h000; 
        10'b1000010101: data <= 9'h000; 
        10'b1000010110: data <= 9'h000; 
        10'b1000010111: data <= 9'h1ff; 
        10'b1000011000: data <= 9'h1ff; 
        10'b1000011001: data <= 9'h000; 
        10'b1000011010: data <= 9'h000; 
        10'b1000011011: data <= 9'h001; 
        10'b1000011100: data <= 9'h001; 
        10'b1000011101: data <= 9'h002; 
        10'b1000011110: data <= 9'h001; 
        10'b1000011111: data <= 9'h000; 
        10'b1000100000: data <= 9'h000; 
        10'b1000100001: data <= 9'h1ff; 
        10'b1000100010: data <= 9'h1ff; 
        10'b1000100011: data <= 9'h000; 
        10'b1000100100: data <= 9'h000; 
        10'b1000100101: data <= 9'h1ff; 
        10'b1000100110: data <= 9'h000; 
        10'b1000100111: data <= 9'h000; 
        10'b1000101000: data <= 9'h001; 
        10'b1000101001: data <= 9'h000; 
        10'b1000101010: data <= 9'h000; 
        10'b1000101011: data <= 9'h000; 
        10'b1000101100: data <= 9'h1ff; 
        10'b1000101101: data <= 9'h000; 
        10'b1000101110: data <= 9'h000; 
        10'b1000101111: data <= 9'h000; 
        10'b1000110000: data <= 9'h000; 
        10'b1000110001: data <= 9'h000; 
        10'b1000110010: data <= 9'h000; 
        10'b1000110011: data <= 9'h000; 
        10'b1000110100: data <= 9'h1ff; 
        10'b1000110101: data <= 9'h000; 
        10'b1000110110: data <= 9'h000; 
        10'b1000110111: data <= 9'h001; 
        10'b1000111000: data <= 9'h000; 
        10'b1000111001: data <= 9'h000; 
        10'b1000111010: data <= 9'h000; 
        10'b1000111011: data <= 9'h1ff; 
        10'b1000111100: data <= 9'h000; 
        10'b1000111101: data <= 9'h000; 
        10'b1000111110: data <= 9'h1ff; 
        10'b1000111111: data <= 9'h000; 
        10'b1001000000: data <= 9'h1ff; 
        10'b1001000001: data <= 9'h000; 
        10'b1001000010: data <= 9'h000; 
        10'b1001000011: data <= 9'h000; 
        10'b1001000100: data <= 9'h000; 
        10'b1001000101: data <= 9'h001; 
        10'b1001000110: data <= 9'h001; 
        10'b1001000111: data <= 9'h000; 
        10'b1001001000: data <= 9'h000; 
        10'b1001001001: data <= 9'h1ff; 
        10'b1001001010: data <= 9'h000; 
        10'b1001001011: data <= 9'h000; 
        10'b1001001100: data <= 9'h000; 
        10'b1001001101: data <= 9'h000; 
        10'b1001001110: data <= 9'h000; 
        10'b1001001111: data <= 9'h1ff; 
        10'b1001010000: data <= 9'h1ff; 
        10'b1001010001: data <= 9'h000; 
        10'b1001010010: data <= 9'h001; 
        10'b1001010011: data <= 9'h001; 
        10'b1001010100: data <= 9'h000; 
        10'b1001010101: data <= 9'h001; 
        10'b1001010110: data <= 9'h000; 
        10'b1001010111: data <= 9'h1ff; 
        10'b1001011000: data <= 9'h000; 
        10'b1001011001: data <= 9'h000; 
        10'b1001011010: data <= 9'h000; 
        10'b1001011011: data <= 9'h000; 
        10'b1001011100: data <= 9'h1ff; 
        10'b1001011101: data <= 9'h000; 
        10'b1001011110: data <= 9'h000; 
        10'b1001011111: data <= 9'h000; 
        10'b1001100000: data <= 9'h000; 
        10'b1001100001: data <= 9'h000; 
        10'b1001100010: data <= 9'h000; 
        10'b1001100011: data <= 9'h000; 
        10'b1001100100: data <= 9'h000; 
        10'b1001100101: data <= 9'h000; 
        10'b1001100110: data <= 9'h000; 
        10'b1001100111: data <= 9'h000; 
        10'b1001101000: data <= 9'h000; 
        10'b1001101001: data <= 9'h000; 
        10'b1001101010: data <= 9'h000; 
        10'b1001101011: data <= 9'h000; 
        10'b1001101100: data <= 9'h1ff; 
        10'b1001101101: data <= 9'h1ff; 
        10'b1001101110: data <= 9'h000; 
        10'b1001101111: data <= 9'h000; 
        10'b1001110000: data <= 9'h000; 
        10'b1001110001: data <= 9'h000; 
        10'b1001110010: data <= 9'h000; 
        10'b1001110011: data <= 9'h000; 
        10'b1001110100: data <= 9'h002; 
        10'b1001110101: data <= 9'h002; 
        10'b1001110110: data <= 9'h001; 
        10'b1001110111: data <= 9'h001; 
        10'b1001111000: data <= 9'h000; 
        10'b1001111001: data <= 9'h000; 
        10'b1001111010: data <= 9'h000; 
        10'b1001111011: data <= 9'h1ff; 
        10'b1001111100: data <= 9'h1ff; 
        10'b1001111101: data <= 9'h000; 
        10'b1001111110: data <= 9'h000; 
        10'b1001111111: data <= 9'h000; 
        10'b1010000000: data <= 9'h000; 
        10'b1010000001: data <= 9'h000; 
        10'b1010000010: data <= 9'h000; 
        10'b1010000011: data <= 9'h000; 
        10'b1010000100: data <= 9'h000; 
        10'b1010000101: data <= 9'h000; 
        10'b1010000110: data <= 9'h000; 
        10'b1010000111: data <= 9'h000; 
        10'b1010001000: data <= 9'h1ff; 
        10'b1010001001: data <= 9'h1fe; 
        10'b1010001010: data <= 9'h1fe; 
        10'b1010001011: data <= 9'h1ff; 
        10'b1010001100: data <= 9'h000; 
        10'b1010001101: data <= 9'h000; 
        10'b1010001110: data <= 9'h001; 
        10'b1010001111: data <= 9'h001; 
        10'b1010010000: data <= 9'h002; 
        10'b1010010001: data <= 9'h003; 
        10'b1010010010: data <= 9'h002; 
        10'b1010010011: data <= 9'h002; 
        10'b1010010100: data <= 9'h002; 
        10'b1010010101: data <= 9'h001; 
        10'b1010010110: data <= 9'h001; 
        10'b1010010111: data <= 9'h001; 
        10'b1010011000: data <= 9'h001; 
        10'b1010011001: data <= 9'h000; 
        10'b1010011010: data <= 9'h000; 
        10'b1010011011: data <= 9'h000; 
        10'b1010011100: data <= 9'h1ff; 
        10'b1010011101: data <= 9'h000; 
        10'b1010011110: data <= 9'h000; 
        10'b1010011111: data <= 9'h000; 
        10'b1010100000: data <= 9'h000; 
        10'b1010100001: data <= 9'h000; 
        10'b1010100010: data <= 9'h000; 
        10'b1010100011: data <= 9'h000; 
        10'b1010100100: data <= 9'h000; 
        10'b1010100101: data <= 9'h1fe; 
        10'b1010100110: data <= 9'h1fe; 
        10'b1010100111: data <= 9'h1fe; 
        10'b1010101000: data <= 9'h000; 
        10'b1010101001: data <= 9'h000; 
        10'b1010101010: data <= 9'h000; 
        10'b1010101011: data <= 9'h001; 
        10'b1010101100: data <= 9'h001; 
        10'b1010101101: data <= 9'h000; 
        10'b1010101110: data <= 9'h001; 
        10'b1010101111: data <= 9'h002; 
        10'b1010110000: data <= 9'h002; 
        10'b1010110001: data <= 9'h001; 
        10'b1010110010: data <= 9'h002; 
        10'b1010110011: data <= 9'h002; 
        10'b1010110100: data <= 9'h001; 
        10'b1010110101: data <= 9'h000; 
        10'b1010110110: data <= 9'h000; 
        10'b1010110111: data <= 9'h000; 
        10'b1010111000: data <= 9'h000; 
        10'b1010111001: data <= 9'h000; 
        10'b1010111010: data <= 9'h000; 
        10'b1010111011: data <= 9'h000; 
        10'b1010111100: data <= 9'h000; 
        10'b1010111101: data <= 9'h000; 
        10'b1010111110: data <= 9'h000; 
        10'b1010111111: data <= 9'h000; 
        10'b1011000000: data <= 9'h000; 
        10'b1011000001: data <= 9'h1ff; 
        10'b1011000010: data <= 9'h1ff; 
        10'b1011000011: data <= 9'h1ff; 
        10'b1011000100: data <= 9'h1ff; 
        10'b1011000101: data <= 9'h1ff; 
        10'b1011000110: data <= 9'h000; 
        10'b1011000111: data <= 9'h1ff; 
        10'b1011001000: data <= 9'h000; 
        10'b1011001001: data <= 9'h000; 
        10'b1011001010: data <= 9'h000; 
        10'b1011001011: data <= 9'h001; 
        10'b1011001100: data <= 9'h001; 
        10'b1011001101: data <= 9'h001; 
        10'b1011001110: data <= 9'h001; 
        10'b1011001111: data <= 9'h000; 
        10'b1011010000: data <= 9'h000; 
        10'b1011010001: data <= 9'h000; 
        10'b1011010010: data <= 9'h000; 
        10'b1011010011: data <= 9'h000; 
        10'b1011010100: data <= 9'h000; 
        10'b1011010101: data <= 9'h000; 
        10'b1011010110: data <= 9'h000; 
        10'b1011010111: data <= 9'h000; 
        10'b1011011000: data <= 9'h000; 
        10'b1011011001: data <= 9'h000; 
        10'b1011011010: data <= 9'h000; 
        10'b1011011011: data <= 9'h000; 
        10'b1011011100: data <= 9'h000; 
        10'b1011011101: data <= 9'h000; 
        10'b1011011110: data <= 9'h1ff; 
        10'b1011011111: data <= 9'h000; 
        10'b1011100000: data <= 9'h1ff; 
        10'b1011100001: data <= 9'h000; 
        10'b1011100010: data <= 9'h1ff; 
        10'b1011100011: data <= 9'h000; 
        10'b1011100100: data <= 9'h000; 
        10'b1011100101: data <= 9'h000; 
        10'b1011100110: data <= 9'h000; 
        10'b1011100111: data <= 9'h000; 
        10'b1011101000: data <= 9'h000; 
        10'b1011101001: data <= 9'h1ff; 
        10'b1011101010: data <= 9'h1ff; 
        10'b1011101011: data <= 9'h000; 
        10'b1011101100: data <= 9'h000; 
        10'b1011101101: data <= 9'h000; 
        10'b1011101110: data <= 9'h000; 
        10'b1011101111: data <= 9'h000; 
        10'b1011110000: data <= 9'h000; 
        10'b1011110001: data <= 9'h000; 
        10'b1011110010: data <= 9'h000; 
        10'b1011110011: data <= 9'h000; 
        10'b1011110100: data <= 9'h000; 
        10'b1011110101: data <= 9'h000; 
        10'b1011110110: data <= 9'h000; 
        10'b1011110111: data <= 9'h000; 
        10'b1011111000: data <= 9'h000; 
        10'b1011111001: data <= 9'h000; 
        10'b1011111010: data <= 9'h000; 
        10'b1011111011: data <= 9'h000; 
        10'b1011111100: data <= 9'h000; 
        10'b1011111101: data <= 9'h000; 
        10'b1011111110: data <= 9'h000; 
        10'b1011111111: data <= 9'h000; 
        10'b1100000000: data <= 9'h000; 
        10'b1100000001: data <= 9'h000; 
        10'b1100000010: data <= 9'h000; 
        10'b1100000011: data <= 9'h000; 
        10'b1100000100: data <= 9'h000; 
        10'b1100000101: data <= 9'h000; 
        10'b1100000110: data <= 9'h000; 
        10'b1100000111: data <= 9'h000; 
        10'b1100001000: data <= 9'h000; 
        10'b1100001001: data <= 9'h000; 
        10'b1100001010: data <= 9'h000; 
        10'b1100001011: data <= 9'h000; 
        10'b1100001100: data <= 9'h000; 
        10'b1100001101: data <= 9'h000; 
        10'b1100001110: data <= 9'h000; 
        10'b1100001111: data <= 9'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 4) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 10'h000; 
        10'b0000000001: data <= 10'h000; 
        10'b0000000010: data <= 10'h000; 
        10'b0000000011: data <= 10'h000; 
        10'b0000000100: data <= 10'h000; 
        10'b0000000101: data <= 10'h000; 
        10'b0000000110: data <= 10'h3ff; 
        10'b0000000111: data <= 10'h000; 
        10'b0000001000: data <= 10'h3ff; 
        10'b0000001001: data <= 10'h3ff; 
        10'b0000001010: data <= 10'h3ff; 
        10'b0000001011: data <= 10'h000; 
        10'b0000001100: data <= 10'h000; 
        10'b0000001101: data <= 10'h000; 
        10'b0000001110: data <= 10'h3ff; 
        10'b0000001111: data <= 10'h000; 
        10'b0000010000: data <= 10'h000; 
        10'b0000010001: data <= 10'h3ff; 
        10'b0000010010: data <= 10'h000; 
        10'b0000010011: data <= 10'h000; 
        10'b0000010100: data <= 10'h000; 
        10'b0000010101: data <= 10'h000; 
        10'b0000010110: data <= 10'h000; 
        10'b0000010111: data <= 10'h000; 
        10'b0000011000: data <= 10'h000; 
        10'b0000011001: data <= 10'h3ff; 
        10'b0000011010: data <= 10'h3ff; 
        10'b0000011011: data <= 10'h000; 
        10'b0000011100: data <= 10'h000; 
        10'b0000011101: data <= 10'h3ff; 
        10'b0000011110: data <= 10'h000; 
        10'b0000011111: data <= 10'h000; 
        10'b0000100000: data <= 10'h3ff; 
        10'b0000100001: data <= 10'h3ff; 
        10'b0000100010: data <= 10'h3ff; 
        10'b0000100011: data <= 10'h3ff; 
        10'b0000100100: data <= 10'h000; 
        10'b0000100101: data <= 10'h000; 
        10'b0000100110: data <= 10'h000; 
        10'b0000100111: data <= 10'h3ff; 
        10'b0000101000: data <= 10'h000; 
        10'b0000101001: data <= 10'h000; 
        10'b0000101010: data <= 10'h3ff; 
        10'b0000101011: data <= 10'h000; 
        10'b0000101100: data <= 10'h000; 
        10'b0000101101: data <= 10'h000; 
        10'b0000101110: data <= 10'h3ff; 
        10'b0000101111: data <= 10'h000; 
        10'b0000110000: data <= 10'h000; 
        10'b0000110001: data <= 10'h3ff; 
        10'b0000110010: data <= 10'h000; 
        10'b0000110011: data <= 10'h3ff; 
        10'b0000110100: data <= 10'h000; 
        10'b0000110101: data <= 10'h000; 
        10'b0000110110: data <= 10'h3ff; 
        10'b0000110111: data <= 10'h3ff; 
        10'b0000111000: data <= 10'h3ff; 
        10'b0000111001: data <= 10'h000; 
        10'b0000111010: data <= 10'h000; 
        10'b0000111011: data <= 10'h000; 
        10'b0000111100: data <= 10'h3ff; 
        10'b0000111101: data <= 10'h3ff; 
        10'b0000111110: data <= 10'h000; 
        10'b0000111111: data <= 10'h3ff; 
        10'b0001000000: data <= 10'h000; 
        10'b0001000001: data <= 10'h3ff; 
        10'b0001000010: data <= 10'h3ff; 
        10'b0001000011: data <= 10'h000; 
        10'b0001000100: data <= 10'h000; 
        10'b0001000101: data <= 10'h3ff; 
        10'b0001000110: data <= 10'h000; 
        10'b0001000111: data <= 10'h000; 
        10'b0001001000: data <= 10'h3ff; 
        10'b0001001001: data <= 10'h3ff; 
        10'b0001001010: data <= 10'h3ff; 
        10'b0001001011: data <= 10'h000; 
        10'b0001001100: data <= 10'h000; 
        10'b0001001101: data <= 10'h000; 
        10'b0001001110: data <= 10'h000; 
        10'b0001001111: data <= 10'h000; 
        10'b0001010000: data <= 10'h000; 
        10'b0001010001: data <= 10'h3ff; 
        10'b0001010010: data <= 10'h000; 
        10'b0001010011: data <= 10'h000; 
        10'b0001010100: data <= 10'h3ff; 
        10'b0001010101: data <= 10'h000; 
        10'b0001010110: data <= 10'h000; 
        10'b0001010111: data <= 10'h3ff; 
        10'b0001011000: data <= 10'h000; 
        10'b0001011001: data <= 10'h3ff; 
        10'b0001011010: data <= 10'h3ff; 
        10'b0001011011: data <= 10'h3ff; 
        10'b0001011100: data <= 10'h3ff; 
        10'b0001011101: data <= 10'h000; 
        10'b0001011110: data <= 10'h3ff; 
        10'b0001011111: data <= 10'h3ff; 
        10'b0001100000: data <= 10'h3ff; 
        10'b0001100001: data <= 10'h3fe; 
        10'b0001100010: data <= 10'h3ff; 
        10'b0001100011: data <= 10'h3ff; 
        10'b0001100100: data <= 10'h3ff; 
        10'b0001100101: data <= 10'h3ff; 
        10'b0001100110: data <= 10'h3ff; 
        10'b0001100111: data <= 10'h000; 
        10'b0001101000: data <= 10'h3ff; 
        10'b0001101001: data <= 10'h000; 
        10'b0001101010: data <= 10'h3ff; 
        10'b0001101011: data <= 10'h000; 
        10'b0001101100: data <= 10'h3ff; 
        10'b0001101101: data <= 10'h000; 
        10'b0001101110: data <= 10'h000; 
        10'b0001101111: data <= 10'h3ff; 
        10'b0001110000: data <= 10'h000; 
        10'b0001110001: data <= 10'h000; 
        10'b0001110010: data <= 10'h3ff; 
        10'b0001110011: data <= 10'h3ff; 
        10'b0001110100: data <= 10'h000; 
        10'b0001110101: data <= 10'h000; 
        10'b0001110110: data <= 10'h000; 
        10'b0001110111: data <= 10'h3ff; 
        10'b0001111000: data <= 10'h3ff; 
        10'b0001111001: data <= 10'h000; 
        10'b0001111010: data <= 10'h000; 
        10'b0001111011: data <= 10'h000; 
        10'b0001111100: data <= 10'h001; 
        10'b0001111101: data <= 10'h001; 
        10'b0001111110: data <= 10'h003; 
        10'b0001111111: data <= 10'h002; 
        10'b0010000000: data <= 10'h001; 
        10'b0010000001: data <= 10'h000; 
        10'b0010000010: data <= 10'h001; 
        10'b0010000011: data <= 10'h3ff; 
        10'b0010000100: data <= 10'h3ff; 
        10'b0010000101: data <= 10'h000; 
        10'b0010000110: data <= 10'h3ff; 
        10'b0010000111: data <= 10'h3ff; 
        10'b0010001000: data <= 10'h000; 
        10'b0010001001: data <= 10'h000; 
        10'b0010001010: data <= 10'h000; 
        10'b0010001011: data <= 10'h000; 
        10'b0010001100: data <= 10'h000; 
        10'b0010001101: data <= 10'h000; 
        10'b0010001110: data <= 10'h000; 
        10'b0010001111: data <= 10'h000; 
        10'b0010010000: data <= 10'h3ff; 
        10'b0010010001: data <= 10'h000; 
        10'b0010010010: data <= 10'h3ff; 
        10'b0010010011: data <= 10'h3fe; 
        10'b0010010100: data <= 10'h3ff; 
        10'b0010010101: data <= 10'h001; 
        10'b0010010110: data <= 10'h3ff; 
        10'b0010010111: data <= 10'h002; 
        10'b0010011000: data <= 10'h003; 
        10'b0010011001: data <= 10'h003; 
        10'b0010011010: data <= 10'h003; 
        10'b0010011011: data <= 10'h001; 
        10'b0010011100: data <= 10'h001; 
        10'b0010011101: data <= 10'h003; 
        10'b0010011110: data <= 10'h000; 
        10'b0010011111: data <= 10'h000; 
        10'b0010100000: data <= 10'h001; 
        10'b0010100001: data <= 10'h001; 
        10'b0010100010: data <= 10'h3fe; 
        10'b0010100011: data <= 10'h3ff; 
        10'b0010100100: data <= 10'h3ff; 
        10'b0010100101: data <= 10'h001; 
        10'b0010100110: data <= 10'h000; 
        10'b0010100111: data <= 10'h000; 
        10'b0010101000: data <= 10'h3ff; 
        10'b0010101001: data <= 10'h3ff; 
        10'b0010101010: data <= 10'h3ff; 
        10'b0010101011: data <= 10'h3ff; 
        10'b0010101100: data <= 10'h3ff; 
        10'b0010101101: data <= 10'h3ff; 
        10'b0010101110: data <= 10'h3fe; 
        10'b0010101111: data <= 10'h3fe; 
        10'b0010110000: data <= 10'h000; 
        10'b0010110001: data <= 10'h000; 
        10'b0010110010: data <= 10'h000; 
        10'b0010110011: data <= 10'h001; 
        10'b0010110100: data <= 10'h001; 
        10'b0010110101: data <= 10'h001; 
        10'b0010110110: data <= 10'h002; 
        10'b0010110111: data <= 10'h003; 
        10'b0010111000: data <= 10'h001; 
        10'b0010111001: data <= 10'h002; 
        10'b0010111010: data <= 10'h000; 
        10'b0010111011: data <= 10'h002; 
        10'b0010111100: data <= 10'h001; 
        10'b0010111101: data <= 10'h001; 
        10'b0010111110: data <= 10'h001; 
        10'b0010111111: data <= 10'h001; 
        10'b0011000000: data <= 10'h001; 
        10'b0011000001: data <= 10'h000; 
        10'b0011000010: data <= 10'h000; 
        10'b0011000011: data <= 10'h000; 
        10'b0011000100: data <= 10'h000; 
        10'b0011000101: data <= 10'h3ff; 
        10'b0011000110: data <= 10'h3ff; 
        10'b0011000111: data <= 10'h3ff; 
        10'b0011001000: data <= 10'h3ff; 
        10'b0011001001: data <= 10'h000; 
        10'b0011001010: data <= 10'h3ff; 
        10'b0011001011: data <= 10'h000; 
        10'b0011001100: data <= 10'h001; 
        10'b0011001101: data <= 10'h000; 
        10'b0011001110: data <= 10'h001; 
        10'b0011001111: data <= 10'h000; 
        10'b0011010000: data <= 10'h3ff; 
        10'b0011010001: data <= 10'h3ff; 
        10'b0011010010: data <= 10'h3fe; 
        10'b0011010011: data <= 10'h001; 
        10'b0011010100: data <= 10'h001; 
        10'b0011010101: data <= 10'h000; 
        10'b0011010110: data <= 10'h001; 
        10'b0011010111: data <= 10'h3ff; 
        10'b0011011000: data <= 10'h001; 
        10'b0011011001: data <= 10'h002; 
        10'b0011011010: data <= 10'h000; 
        10'b0011011011: data <= 10'h004; 
        10'b0011011100: data <= 10'h002; 
        10'b0011011101: data <= 10'h000; 
        10'b0011011110: data <= 10'h000; 
        10'b0011011111: data <= 10'h000; 
        10'b0011100000: data <= 10'h000; 
        10'b0011100001: data <= 10'h000; 
        10'b0011100010: data <= 10'h000; 
        10'b0011100011: data <= 10'h3ff; 
        10'b0011100100: data <= 10'h000; 
        10'b0011100101: data <= 10'h000; 
        10'b0011100110: data <= 10'h002; 
        10'b0011100111: data <= 10'h001; 
        10'b0011101000: data <= 10'h000; 
        10'b0011101001: data <= 10'h003; 
        10'b0011101010: data <= 10'h000; 
        10'b0011101011: data <= 10'h000; 
        10'b0011101100: data <= 10'h002; 
        10'b0011101101: data <= 10'h002; 
        10'b0011101110: data <= 10'h3fe; 
        10'b0011101111: data <= 10'h3fe; 
        10'b0011110000: data <= 10'h001; 
        10'b0011110001: data <= 10'h3ff; 
        10'b0011110010: data <= 10'h000; 
        10'b0011110011: data <= 10'h001; 
        10'b0011110100: data <= 10'h001; 
        10'b0011110101: data <= 10'h002; 
        10'b0011110110: data <= 10'h002; 
        10'b0011110111: data <= 10'h003; 
        10'b0011111000: data <= 10'h003; 
        10'b0011111001: data <= 10'h000; 
        10'b0011111010: data <= 10'h000; 
        10'b0011111011: data <= 10'h000; 
        10'b0011111100: data <= 10'h000; 
        10'b0011111101: data <= 10'h000; 
        10'b0011111110: data <= 10'h000; 
        10'b0011111111: data <= 10'h000; 
        10'b0100000000: data <= 10'h000; 
        10'b0100000001: data <= 10'h002; 
        10'b0100000010: data <= 10'h001; 
        10'b0100000011: data <= 10'h002; 
        10'b0100000100: data <= 10'h003; 
        10'b0100000101: data <= 10'h003; 
        10'b0100000110: data <= 10'h002; 
        10'b0100000111: data <= 10'h003; 
        10'b0100001000: data <= 10'h001; 
        10'b0100001001: data <= 10'h001; 
        10'b0100001010: data <= 10'h3fc; 
        10'b0100001011: data <= 10'h3fb; 
        10'b0100001100: data <= 10'h3fe; 
        10'b0100001101: data <= 10'h000; 
        10'b0100001110: data <= 10'h001; 
        10'b0100001111: data <= 10'h001; 
        10'b0100010000: data <= 10'h001; 
        10'b0100010001: data <= 10'h001; 
        10'b0100010010: data <= 10'h003; 
        10'b0100010011: data <= 10'h003; 
        10'b0100010100: data <= 10'h000; 
        10'b0100010101: data <= 10'h000; 
        10'b0100010110: data <= 10'h001; 
        10'b0100010111: data <= 10'h3ff; 
        10'b0100011000: data <= 10'h3ff; 
        10'b0100011001: data <= 10'h000; 
        10'b0100011010: data <= 10'h3ff; 
        10'b0100011011: data <= 10'h000; 
        10'b0100011100: data <= 10'h001; 
        10'b0100011101: data <= 10'h002; 
        10'b0100011110: data <= 10'h002; 
        10'b0100011111: data <= 10'h004; 
        10'b0100100000: data <= 10'h003; 
        10'b0100100001: data <= 10'h003; 
        10'b0100100010: data <= 10'h004; 
        10'b0100100011: data <= 10'h002; 
        10'b0100100100: data <= 10'h002; 
        10'b0100100101: data <= 10'h002; 
        10'b0100100110: data <= 10'h3ff; 
        10'b0100100111: data <= 10'h3fb; 
        10'b0100101000: data <= 10'h3fc; 
        10'b0100101001: data <= 10'h3ff; 
        10'b0100101010: data <= 10'h001; 
        10'b0100101011: data <= 10'h001; 
        10'b0100101100: data <= 10'h001; 
        10'b0100101101: data <= 10'h003; 
        10'b0100101110: data <= 10'h004; 
        10'b0100101111: data <= 10'h003; 
        10'b0100110000: data <= 10'h000; 
        10'b0100110001: data <= 10'h000; 
        10'b0100110010: data <= 10'h000; 
        10'b0100110011: data <= 10'h3ff; 
        10'b0100110100: data <= 10'h3ff; 
        10'b0100110101: data <= 10'h000; 
        10'b0100110110: data <= 10'h000; 
        10'b0100110111: data <= 10'h3ff; 
        10'b0100111000: data <= 10'h001; 
        10'b0100111001: data <= 10'h002; 
        10'b0100111010: data <= 10'h004; 
        10'b0100111011: data <= 10'h005; 
        10'b0100111100: data <= 10'h004; 
        10'b0100111101: data <= 10'h005; 
        10'b0100111110: data <= 10'h004; 
        10'b0100111111: data <= 10'h002; 
        10'b0101000000: data <= 10'h002; 
        10'b0101000001: data <= 10'h005; 
        10'b0101000010: data <= 10'h006; 
        10'b0101000011: data <= 10'h3ff; 
        10'b0101000100: data <= 10'h3fc; 
        10'b0101000101: data <= 10'h3ff; 
        10'b0101000110: data <= 10'h3ff; 
        10'b0101000111: data <= 10'h001; 
        10'b0101001000: data <= 10'h003; 
        10'b0101001001: data <= 10'h003; 
        10'b0101001010: data <= 10'h005; 
        10'b0101001011: data <= 10'h004; 
        10'b0101001100: data <= 10'h003; 
        10'b0101001101: data <= 10'h000; 
        10'b0101001110: data <= 10'h000; 
        10'b0101001111: data <= 10'h000; 
        10'b0101010000: data <= 10'h3ff; 
        10'b0101010001: data <= 10'h000; 
        10'b0101010010: data <= 10'h3ff; 
        10'b0101010011: data <= 10'h000; 
        10'b0101010100: data <= 10'h000; 
        10'b0101010101: data <= 10'h003; 
        10'b0101010110: data <= 10'h002; 
        10'b0101010111: data <= 10'h003; 
        10'b0101011000: data <= 10'h003; 
        10'b0101011001: data <= 10'h004; 
        10'b0101011010: data <= 10'h001; 
        10'b0101011011: data <= 10'h001; 
        10'b0101011100: data <= 10'h001; 
        10'b0101011101: data <= 10'h006; 
        10'b0101011110: data <= 10'h006; 
        10'b0101011111: data <= 10'h001; 
        10'b0101100000: data <= 10'h000; 
        10'b0101100001: data <= 10'h3ff; 
        10'b0101100010: data <= 10'h000; 
        10'b0101100011: data <= 10'h002; 
        10'b0101100100: data <= 10'h003; 
        10'b0101100101: data <= 10'h005; 
        10'b0101100110: data <= 10'h005; 
        10'b0101100111: data <= 10'h004; 
        10'b0101101000: data <= 10'h003; 
        10'b0101101001: data <= 10'h001; 
        10'b0101101010: data <= 10'h001; 
        10'b0101101011: data <= 10'h3ff; 
        10'b0101101100: data <= 10'h3ff; 
        10'b0101101101: data <= 10'h000; 
        10'b0101101110: data <= 10'h000; 
        10'b0101101111: data <= 10'h3ff; 
        10'b0101110000: data <= 10'h3ff; 
        10'b0101110001: data <= 10'h000; 
        10'b0101110010: data <= 10'h000; 
        10'b0101110011: data <= 10'h000; 
        10'b0101110100: data <= 10'h000; 
        10'b0101110101: data <= 10'h000; 
        10'b0101110110: data <= 10'h3ff; 
        10'b0101110111: data <= 10'h001; 
        10'b0101111000: data <= 10'h002; 
        10'b0101111001: data <= 10'h006; 
        10'b0101111010: data <= 10'h002; 
        10'b0101111011: data <= 10'h004; 
        10'b0101111100: data <= 10'h002; 
        10'b0101111101: data <= 10'h3ff; 
        10'b0101111110: data <= 10'h000; 
        10'b0101111111: data <= 10'h000; 
        10'b0110000000: data <= 10'h002; 
        10'b0110000001: data <= 10'h002; 
        10'b0110000010: data <= 10'h001; 
        10'b0110000011: data <= 10'h001; 
        10'b0110000100: data <= 10'h001; 
        10'b0110000101: data <= 10'h000; 
        10'b0110000110: data <= 10'h000; 
        10'b0110000111: data <= 10'h000; 
        10'b0110001000: data <= 10'h3ff; 
        10'b0110001001: data <= 10'h3ff; 
        10'b0110001010: data <= 10'h000; 
        10'b0110001011: data <= 10'h000; 
        10'b0110001100: data <= 10'h3ff; 
        10'b0110001101: data <= 10'h3fe; 
        10'b0110001110: data <= 10'h3fd; 
        10'b0110001111: data <= 10'h3fc; 
        10'b0110010000: data <= 10'h3fb; 
        10'b0110010001: data <= 10'h3fc; 
        10'b0110010010: data <= 10'h3ff; 
        10'b0110010011: data <= 10'h002; 
        10'b0110010100: data <= 10'h002; 
        10'b0110010101: data <= 10'h005; 
        10'b0110010110: data <= 10'h004; 
        10'b0110010111: data <= 10'h003; 
        10'b0110011000: data <= 10'h000; 
        10'b0110011001: data <= 10'h000; 
        10'b0110011010: data <= 10'h3ff; 
        10'b0110011011: data <= 10'h3fe; 
        10'b0110011100: data <= 10'h3fd; 
        10'b0110011101: data <= 10'h3fe; 
        10'b0110011110: data <= 10'h3fe; 
        10'b0110011111: data <= 10'h3fe; 
        10'b0110100000: data <= 10'h3ff; 
        10'b0110100001: data <= 10'h000; 
        10'b0110100010: data <= 10'h3ff; 
        10'b0110100011: data <= 10'h000; 
        10'b0110100100: data <= 10'h000; 
        10'b0110100101: data <= 10'h3ff; 
        10'b0110100110: data <= 10'h3ff; 
        10'b0110100111: data <= 10'h000; 
        10'b0110101000: data <= 10'h3ff; 
        10'b0110101001: data <= 10'h3fe; 
        10'b0110101010: data <= 10'h3fc; 
        10'b0110101011: data <= 10'h3fb; 
        10'b0110101100: data <= 10'h3fc; 
        10'b0110101101: data <= 10'h3ff; 
        10'b0110101110: data <= 10'h000; 
        10'b0110101111: data <= 10'h000; 
        10'b0110110000: data <= 10'h003; 
        10'b0110110001: data <= 10'h004; 
        10'b0110110010: data <= 10'h003; 
        10'b0110110011: data <= 10'h002; 
        10'b0110110100: data <= 10'h3ff; 
        10'b0110110101: data <= 10'h3ff; 
        10'b0110110110: data <= 10'h3ff; 
        10'b0110110111: data <= 10'h3fd; 
        10'b0110111000: data <= 10'h3fc; 
        10'b0110111001: data <= 10'h3fd; 
        10'b0110111010: data <= 10'h3fe; 
        10'b0110111011: data <= 10'h3fe; 
        10'b0110111100: data <= 10'h3fe; 
        10'b0110111101: data <= 10'h000; 
        10'b0110111110: data <= 10'h3ff; 
        10'b0110111111: data <= 10'h000; 
        10'b0111000000: data <= 10'h000; 
        10'b0111000001: data <= 10'h3ff; 
        10'b0111000010: data <= 10'h3ff; 
        10'b0111000011: data <= 10'h000; 
        10'b0111000100: data <= 10'h3ff; 
        10'b0111000101: data <= 10'h3fe; 
        10'b0111000110: data <= 10'h3fc; 
        10'b0111000111: data <= 10'h3fe; 
        10'b0111001000: data <= 10'h002; 
        10'b0111001001: data <= 10'h002; 
        10'b0111001010: data <= 10'h001; 
        10'b0111001011: data <= 10'h002; 
        10'b0111001100: data <= 10'h003; 
        10'b0111001101: data <= 10'h003; 
        10'b0111001110: data <= 10'h001; 
        10'b0111001111: data <= 10'h002; 
        10'b0111010000: data <= 10'h001; 
        10'b0111010001: data <= 10'h3ff; 
        10'b0111010010: data <= 10'h3fd; 
        10'b0111010011: data <= 10'h3fc; 
        10'b0111010100: data <= 10'h3fc; 
        10'b0111010101: data <= 10'h3fc; 
        10'b0111010110: data <= 10'h3fd; 
        10'b0111010111: data <= 10'h3ff; 
        10'b0111011000: data <= 10'h3ff; 
        10'b0111011001: data <= 10'h000; 
        10'b0111011010: data <= 10'h3ff; 
        10'b0111011011: data <= 10'h3ff; 
        10'b0111011100: data <= 10'h000; 
        10'b0111011101: data <= 10'h000; 
        10'b0111011110: data <= 10'h3ff; 
        10'b0111011111: data <= 10'h3ff; 
        10'b0111100000: data <= 10'h3ff; 
        10'b0111100001: data <= 10'h3fd; 
        10'b0111100010: data <= 10'h3fd; 
        10'b0111100011: data <= 10'h001; 
        10'b0111100100: data <= 10'h003; 
        10'b0111100101: data <= 10'h004; 
        10'b0111100110: data <= 10'h001; 
        10'b0111100111: data <= 10'h003; 
        10'b0111101000: data <= 10'h005; 
        10'b0111101001: data <= 10'h003; 
        10'b0111101010: data <= 10'h000; 
        10'b0111101011: data <= 10'h3ff; 
        10'b0111101100: data <= 10'h000; 
        10'b0111101101: data <= 10'h3fe; 
        10'b0111101110: data <= 10'h3fc; 
        10'b0111101111: data <= 10'h3fe; 
        10'b0111110000: data <= 10'h3fe; 
        10'b0111110001: data <= 10'h3fd; 
        10'b0111110010: data <= 10'h3fe; 
        10'b0111110011: data <= 10'h3ff; 
        10'b0111110100: data <= 10'h3ff; 
        10'b0111110101: data <= 10'h3ff; 
        10'b0111110110: data <= 10'h000; 
        10'b0111110111: data <= 10'h3ff; 
        10'b0111111000: data <= 10'h3ff; 
        10'b0111111001: data <= 10'h000; 
        10'b0111111010: data <= 10'h3ff; 
        10'b0111111011: data <= 10'h3ff; 
        10'b0111111100: data <= 10'h3fe; 
        10'b0111111101: data <= 10'h3fe; 
        10'b0111111110: data <= 10'h3ff; 
        10'b0111111111: data <= 10'h001; 
        10'b1000000000: data <= 10'h003; 
        10'b1000000001: data <= 10'h005; 
        10'b1000000010: data <= 10'h003; 
        10'b1000000011: data <= 10'h005; 
        10'b1000000100: data <= 10'h003; 
        10'b1000000101: data <= 10'h002; 
        10'b1000000110: data <= 10'h3fe; 
        10'b1000000111: data <= 10'h3ff; 
        10'b1000001000: data <= 10'h3ff; 
        10'b1000001001: data <= 10'h3fd; 
        10'b1000001010: data <= 10'h3ff; 
        10'b1000001011: data <= 10'h3ff; 
        10'b1000001100: data <= 10'h000; 
        10'b1000001101: data <= 10'h3fe; 
        10'b1000001110: data <= 10'h000; 
        10'b1000001111: data <= 10'h3ff; 
        10'b1000010000: data <= 10'h3fe; 
        10'b1000010001: data <= 10'h3ff; 
        10'b1000010010: data <= 10'h000; 
        10'b1000010011: data <= 10'h000; 
        10'b1000010100: data <= 10'h3ff; 
        10'b1000010101: data <= 10'h000; 
        10'b1000010110: data <= 10'h000; 
        10'b1000010111: data <= 10'h3ff; 
        10'b1000011000: data <= 10'h3fe; 
        10'b1000011001: data <= 10'h3ff; 
        10'b1000011010: data <= 10'h000; 
        10'b1000011011: data <= 10'h001; 
        10'b1000011100: data <= 10'h001; 
        10'b1000011101: data <= 10'h003; 
        10'b1000011110: data <= 10'h002; 
        10'b1000011111: data <= 10'h000; 
        10'b1000100000: data <= 10'h001; 
        10'b1000100001: data <= 10'h3fe; 
        10'b1000100010: data <= 10'h3fd; 
        10'b1000100011: data <= 10'h3ff; 
        10'b1000100100: data <= 10'h3ff; 
        10'b1000100101: data <= 10'h3ff; 
        10'b1000100110: data <= 10'h001; 
        10'b1000100111: data <= 10'h000; 
        10'b1000101000: data <= 10'h001; 
        10'b1000101001: data <= 10'h000; 
        10'b1000101010: data <= 10'h001; 
        10'b1000101011: data <= 10'h3ff; 
        10'b1000101100: data <= 10'h3fe; 
        10'b1000101101: data <= 10'h3ff; 
        10'b1000101110: data <= 10'h3ff; 
        10'b1000101111: data <= 10'h000; 
        10'b1000110000: data <= 10'h3ff; 
        10'b1000110001: data <= 10'h000; 
        10'b1000110010: data <= 10'h3ff; 
        10'b1000110011: data <= 10'h3ff; 
        10'b1000110100: data <= 10'h3fe; 
        10'b1000110101: data <= 10'h000; 
        10'b1000110110: data <= 10'h000; 
        10'b1000110111: data <= 10'h003; 
        10'b1000111000: data <= 10'h001; 
        10'b1000111001: data <= 10'h000; 
        10'b1000111010: data <= 10'h000; 
        10'b1000111011: data <= 10'h3fe; 
        10'b1000111100: data <= 10'h000; 
        10'b1000111101: data <= 10'h000; 
        10'b1000111110: data <= 10'h3fe; 
        10'b1000111111: data <= 10'h000; 
        10'b1001000000: data <= 10'h3fd; 
        10'b1001000001: data <= 10'h3ff; 
        10'b1001000010: data <= 10'h000; 
        10'b1001000011: data <= 10'h000; 
        10'b1001000100: data <= 10'h001; 
        10'b1001000101: data <= 10'h001; 
        10'b1001000110: data <= 10'h001; 
        10'b1001000111: data <= 10'h000; 
        10'b1001001000: data <= 10'h3ff; 
        10'b1001001001: data <= 10'h3ff; 
        10'b1001001010: data <= 10'h000; 
        10'b1001001011: data <= 10'h3ff; 
        10'b1001001100: data <= 10'h000; 
        10'b1001001101: data <= 10'h000; 
        10'b1001001110: data <= 10'h000; 
        10'b1001001111: data <= 10'h3fe; 
        10'b1001010000: data <= 10'h3fe; 
        10'b1001010001: data <= 10'h000; 
        10'b1001010010: data <= 10'h001; 
        10'b1001010011: data <= 10'h003; 
        10'b1001010100: data <= 10'h001; 
        10'b1001010101: data <= 10'h001; 
        10'b1001010110: data <= 10'h000; 
        10'b1001010111: data <= 10'h3fe; 
        10'b1001011000: data <= 10'h3ff; 
        10'b1001011001: data <= 10'h001; 
        10'b1001011010: data <= 10'h000; 
        10'b1001011011: data <= 10'h000; 
        10'b1001011100: data <= 10'h3fe; 
        10'b1001011101: data <= 10'h3ff; 
        10'b1001011110: data <= 10'h3ff; 
        10'b1001011111: data <= 10'h000; 
        10'b1001100000: data <= 10'h000; 
        10'b1001100001: data <= 10'h000; 
        10'b1001100010: data <= 10'h000; 
        10'b1001100011: data <= 10'h3ff; 
        10'b1001100100: data <= 10'h3ff; 
        10'b1001100101: data <= 10'h000; 
        10'b1001100110: data <= 10'h000; 
        10'b1001100111: data <= 10'h000; 
        10'b1001101000: data <= 10'h000; 
        10'b1001101001: data <= 10'h3ff; 
        10'b1001101010: data <= 10'h3ff; 
        10'b1001101011: data <= 10'h3ff; 
        10'b1001101100: data <= 10'h3fe; 
        10'b1001101101: data <= 10'h3fd; 
        10'b1001101110: data <= 10'h000; 
        10'b1001101111: data <= 10'h001; 
        10'b1001110000: data <= 10'h000; 
        10'b1001110001: data <= 10'h3ff; 
        10'b1001110010: data <= 10'h001; 
        10'b1001110011: data <= 10'h000; 
        10'b1001110100: data <= 10'h003; 
        10'b1001110101: data <= 10'h003; 
        10'b1001110110: data <= 10'h002; 
        10'b1001110111: data <= 10'h002; 
        10'b1001111000: data <= 10'h000; 
        10'b1001111001: data <= 10'h000; 
        10'b1001111010: data <= 10'h001; 
        10'b1001111011: data <= 10'h3ff; 
        10'b1001111100: data <= 10'h3ff; 
        10'b1001111101: data <= 10'h000; 
        10'b1001111110: data <= 10'h000; 
        10'b1001111111: data <= 10'h3ff; 
        10'b1010000000: data <= 10'h000; 
        10'b1010000001: data <= 10'h000; 
        10'b1010000010: data <= 10'h000; 
        10'b1010000011: data <= 10'h3ff; 
        10'b1010000100: data <= 10'h3ff; 
        10'b1010000101: data <= 10'h000; 
        10'b1010000110: data <= 10'h000; 
        10'b1010000111: data <= 10'h3ff; 
        10'b1010001000: data <= 10'h3fe; 
        10'b1010001001: data <= 10'h3fb; 
        10'b1010001010: data <= 10'h3fc; 
        10'b1010001011: data <= 10'h3fe; 
        10'b1010001100: data <= 10'h001; 
        10'b1010001101: data <= 10'h001; 
        10'b1010001110: data <= 10'h001; 
        10'b1010001111: data <= 10'h002; 
        10'b1010010000: data <= 10'h004; 
        10'b1010010001: data <= 10'h006; 
        10'b1010010010: data <= 10'h005; 
        10'b1010010011: data <= 10'h004; 
        10'b1010010100: data <= 10'h003; 
        10'b1010010101: data <= 10'h002; 
        10'b1010010110: data <= 10'h002; 
        10'b1010010111: data <= 10'h002; 
        10'b1010011000: data <= 10'h002; 
        10'b1010011001: data <= 10'h000; 
        10'b1010011010: data <= 10'h000; 
        10'b1010011011: data <= 10'h3ff; 
        10'b1010011100: data <= 10'h3ff; 
        10'b1010011101: data <= 10'h000; 
        10'b1010011110: data <= 10'h3ff; 
        10'b1010011111: data <= 10'h000; 
        10'b1010100000: data <= 10'h000; 
        10'b1010100001: data <= 10'h000; 
        10'b1010100010: data <= 10'h000; 
        10'b1010100011: data <= 10'h3ff; 
        10'b1010100100: data <= 10'h3ff; 
        10'b1010100101: data <= 10'h3fd; 
        10'b1010100110: data <= 10'h3fc; 
        10'b1010100111: data <= 10'h3fc; 
        10'b1010101000: data <= 10'h000; 
        10'b1010101001: data <= 10'h001; 
        10'b1010101010: data <= 10'h000; 
        10'b1010101011: data <= 10'h002; 
        10'b1010101100: data <= 10'h001; 
        10'b1010101101: data <= 10'h001; 
        10'b1010101110: data <= 10'h002; 
        10'b1010101111: data <= 10'h004; 
        10'b1010110000: data <= 10'h004; 
        10'b1010110001: data <= 10'h003; 
        10'b1010110010: data <= 10'h004; 
        10'b1010110011: data <= 10'h004; 
        10'b1010110100: data <= 10'h001; 
        10'b1010110101: data <= 10'h000; 
        10'b1010110110: data <= 10'h3ff; 
        10'b1010110111: data <= 10'h000; 
        10'b1010111000: data <= 10'h000; 
        10'b1010111001: data <= 10'h3ff; 
        10'b1010111010: data <= 10'h000; 
        10'b1010111011: data <= 10'h000; 
        10'b1010111100: data <= 10'h000; 
        10'b1010111101: data <= 10'h000; 
        10'b1010111110: data <= 10'h000; 
        10'b1010111111: data <= 10'h3ff; 
        10'b1011000000: data <= 10'h3ff; 
        10'b1011000001: data <= 10'h3ff; 
        10'b1011000010: data <= 10'h3fe; 
        10'b1011000011: data <= 10'h3fe; 
        10'b1011000100: data <= 10'h3fe; 
        10'b1011000101: data <= 10'h3fe; 
        10'b1011000110: data <= 10'h3ff; 
        10'b1011000111: data <= 10'h3fe; 
        10'b1011001000: data <= 10'h3ff; 
        10'b1011001001: data <= 10'h3ff; 
        10'b1011001010: data <= 10'h000; 
        10'b1011001011: data <= 10'h001; 
        10'b1011001100: data <= 10'h001; 
        10'b1011001101: data <= 10'h001; 
        10'b1011001110: data <= 10'h001; 
        10'b1011001111: data <= 10'h000; 
        10'b1011010000: data <= 10'h000; 
        10'b1011010001: data <= 10'h000; 
        10'b1011010010: data <= 10'h3ff; 
        10'b1011010011: data <= 10'h3ff; 
        10'b1011010100: data <= 10'h000; 
        10'b1011010101: data <= 10'h000; 
        10'b1011010110: data <= 10'h3ff; 
        10'b1011010111: data <= 10'h000; 
        10'b1011011000: data <= 10'h000; 
        10'b1011011001: data <= 10'h000; 
        10'b1011011010: data <= 10'h000; 
        10'b1011011011: data <= 10'h3ff; 
        10'b1011011100: data <= 10'h3ff; 
        10'b1011011101: data <= 10'h3ff; 
        10'b1011011110: data <= 10'h3ff; 
        10'b1011011111: data <= 10'h000; 
        10'b1011100000: data <= 10'h3ff; 
        10'b1011100001: data <= 10'h3ff; 
        10'b1011100010: data <= 10'h3ff; 
        10'b1011100011: data <= 10'h3ff; 
        10'b1011100100: data <= 10'h3ff; 
        10'b1011100101: data <= 10'h3ff; 
        10'b1011100110: data <= 10'h3ff; 
        10'b1011100111: data <= 10'h3ff; 
        10'b1011101000: data <= 10'h3ff; 
        10'b1011101001: data <= 10'h3ff; 
        10'b1011101010: data <= 10'h3ff; 
        10'b1011101011: data <= 10'h3ff; 
        10'b1011101100: data <= 10'h3ff; 
        10'b1011101101: data <= 10'h000; 
        10'b1011101110: data <= 10'h000; 
        10'b1011101111: data <= 10'h000; 
        10'b1011110000: data <= 10'h000; 
        10'b1011110001: data <= 10'h3ff; 
        10'b1011110010: data <= 10'h000; 
        10'b1011110011: data <= 10'h000; 
        10'b1011110100: data <= 10'h000; 
        10'b1011110101: data <= 10'h3ff; 
        10'b1011110110: data <= 10'h000; 
        10'b1011110111: data <= 10'h000; 
        10'b1011111000: data <= 10'h000; 
        10'b1011111001: data <= 10'h3ff; 
        10'b1011111010: data <= 10'h000; 
        10'b1011111011: data <= 10'h3ff; 
        10'b1011111100: data <= 10'h000; 
        10'b1011111101: data <= 10'h000; 
        10'b1011111110: data <= 10'h3ff; 
        10'b1011111111: data <= 10'h000; 
        10'b1100000000: data <= 10'h3ff; 
        10'b1100000001: data <= 10'h3ff; 
        10'b1100000010: data <= 10'h000; 
        10'b1100000011: data <= 10'h000; 
        10'b1100000100: data <= 10'h000; 
        10'b1100000101: data <= 10'h000; 
        10'b1100000110: data <= 10'h000; 
        10'b1100000111: data <= 10'h000; 
        10'b1100001000: data <= 10'h000; 
        10'b1100001001: data <= 10'h000; 
        10'b1100001010: data <= 10'h000; 
        10'b1100001011: data <= 10'h3ff; 
        10'b1100001100: data <= 10'h000; 
        10'b1100001101: data <= 10'h000; 
        10'b1100001110: data <= 10'h3ff; 
        10'b1100001111: data <= 10'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 5) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 11'h7ff; 
        10'b0000000001: data <= 11'h7ff; 
        10'b0000000010: data <= 11'h7ff; 
        10'b0000000011: data <= 11'h000; 
        10'b0000000100: data <= 11'h7ff; 
        10'b0000000101: data <= 11'h000; 
        10'b0000000110: data <= 11'h7fe; 
        10'b0000000111: data <= 11'h000; 
        10'b0000001000: data <= 11'h7ff; 
        10'b0000001001: data <= 11'h7ff; 
        10'b0000001010: data <= 11'h7ff; 
        10'b0000001011: data <= 11'h000; 
        10'b0000001100: data <= 11'h7ff; 
        10'b0000001101: data <= 11'h000; 
        10'b0000001110: data <= 11'h7fe; 
        10'b0000001111: data <= 11'h000; 
        10'b0000010000: data <= 11'h000; 
        10'b0000010001: data <= 11'h7fe; 
        10'b0000010010: data <= 11'h000; 
        10'b0000010011: data <= 11'h7ff; 
        10'b0000010100: data <= 11'h7ff; 
        10'b0000010101: data <= 11'h7ff; 
        10'b0000010110: data <= 11'h7ff; 
        10'b0000010111: data <= 11'h000; 
        10'b0000011000: data <= 11'h000; 
        10'b0000011001: data <= 11'h7ff; 
        10'b0000011010: data <= 11'h7ff; 
        10'b0000011011: data <= 11'h7ff; 
        10'b0000011100: data <= 11'h7ff; 
        10'b0000011101: data <= 11'h7fe; 
        10'b0000011110: data <= 11'h000; 
        10'b0000011111: data <= 11'h000; 
        10'b0000100000: data <= 11'h7fe; 
        10'b0000100001: data <= 11'h7fe; 
        10'b0000100010: data <= 11'h7fe; 
        10'b0000100011: data <= 11'h7fe; 
        10'b0000100100: data <= 11'h000; 
        10'b0000100101: data <= 11'h7ff; 
        10'b0000100110: data <= 11'h7ff; 
        10'b0000100111: data <= 11'h7fe; 
        10'b0000101000: data <= 11'h000; 
        10'b0000101001: data <= 11'h000; 
        10'b0000101010: data <= 11'h7ff; 
        10'b0000101011: data <= 11'h7ff; 
        10'b0000101100: data <= 11'h000; 
        10'b0000101101: data <= 11'h7ff; 
        10'b0000101110: data <= 11'h7ff; 
        10'b0000101111: data <= 11'h7ff; 
        10'b0000110000: data <= 11'h000; 
        10'b0000110001: data <= 11'h7fe; 
        10'b0000110010: data <= 11'h000; 
        10'b0000110011: data <= 11'h7ff; 
        10'b0000110100: data <= 11'h000; 
        10'b0000110101: data <= 11'h000; 
        10'b0000110110: data <= 11'h7ff; 
        10'b0000110111: data <= 11'h7ff; 
        10'b0000111000: data <= 11'h7fe; 
        10'b0000111001: data <= 11'h000; 
        10'b0000111010: data <= 11'h7ff; 
        10'b0000111011: data <= 11'h7ff; 
        10'b0000111100: data <= 11'h7ff; 
        10'b0000111101: data <= 11'h7fe; 
        10'b0000111110: data <= 11'h7ff; 
        10'b0000111111: data <= 11'h7fe; 
        10'b0001000000: data <= 11'h000; 
        10'b0001000001: data <= 11'h7fe; 
        10'b0001000010: data <= 11'h7fe; 
        10'b0001000011: data <= 11'h000; 
        10'b0001000100: data <= 11'h7ff; 
        10'b0001000101: data <= 11'h7fe; 
        10'b0001000110: data <= 11'h000; 
        10'b0001000111: data <= 11'h7ff; 
        10'b0001001000: data <= 11'h7fe; 
        10'b0001001001: data <= 11'h7ff; 
        10'b0001001010: data <= 11'h7ff; 
        10'b0001001011: data <= 11'h000; 
        10'b0001001100: data <= 11'h000; 
        10'b0001001101: data <= 11'h000; 
        10'b0001001110: data <= 11'h000; 
        10'b0001001111: data <= 11'h7ff; 
        10'b0001010000: data <= 11'h000; 
        10'b0001010001: data <= 11'h7ff; 
        10'b0001010010: data <= 11'h000; 
        10'b0001010011: data <= 11'h000; 
        10'b0001010100: data <= 11'h7ff; 
        10'b0001010101: data <= 11'h7ff; 
        10'b0001010110: data <= 11'h7ff; 
        10'b0001010111: data <= 11'h7fe; 
        10'b0001011000: data <= 11'h000; 
        10'b0001011001: data <= 11'h7fe; 
        10'b0001011010: data <= 11'h7fe; 
        10'b0001011011: data <= 11'h7ff; 
        10'b0001011100: data <= 11'h7fe; 
        10'b0001011101: data <= 11'h7ff; 
        10'b0001011110: data <= 11'h7ff; 
        10'b0001011111: data <= 11'h7fd; 
        10'b0001100000: data <= 11'h7fd; 
        10'b0001100001: data <= 11'h7fd; 
        10'b0001100010: data <= 11'h7fd; 
        10'b0001100011: data <= 11'h7fe; 
        10'b0001100100: data <= 11'h7fd; 
        10'b0001100101: data <= 11'h7fe; 
        10'b0001100110: data <= 11'h7fe; 
        10'b0001100111: data <= 11'h7ff; 
        10'b0001101000: data <= 11'h7fe; 
        10'b0001101001: data <= 11'h000; 
        10'b0001101010: data <= 11'h7ff; 
        10'b0001101011: data <= 11'h000; 
        10'b0001101100: data <= 11'h7ff; 
        10'b0001101101: data <= 11'h000; 
        10'b0001101110: data <= 11'h7ff; 
        10'b0001101111: data <= 11'h7fe; 
        10'b0001110000: data <= 11'h7ff; 
        10'b0001110001: data <= 11'h000; 
        10'b0001110010: data <= 11'h7ff; 
        10'b0001110011: data <= 11'h7fe; 
        10'b0001110100: data <= 11'h000; 
        10'b0001110101: data <= 11'h000; 
        10'b0001110110: data <= 11'h7ff; 
        10'b0001110111: data <= 11'h7fe; 
        10'b0001111000: data <= 11'h7fe; 
        10'b0001111001: data <= 11'h7ff; 
        10'b0001111010: data <= 11'h7ff; 
        10'b0001111011: data <= 11'h000; 
        10'b0001111100: data <= 11'h002; 
        10'b0001111101: data <= 11'h002; 
        10'b0001111110: data <= 11'h005; 
        10'b0001111111: data <= 11'h004; 
        10'b0010000000: data <= 11'h002; 
        10'b0010000001: data <= 11'h001; 
        10'b0010000010: data <= 11'h002; 
        10'b0010000011: data <= 11'h7ff; 
        10'b0010000100: data <= 11'h7fe; 
        10'b0010000101: data <= 11'h7ff; 
        10'b0010000110: data <= 11'h7fe; 
        10'b0010000111: data <= 11'h7fe; 
        10'b0010001000: data <= 11'h000; 
        10'b0010001001: data <= 11'h000; 
        10'b0010001010: data <= 11'h7ff; 
        10'b0010001011: data <= 11'h7ff; 
        10'b0010001100: data <= 11'h7ff; 
        10'b0010001101: data <= 11'h000; 
        10'b0010001110: data <= 11'h000; 
        10'b0010001111: data <= 11'h000; 
        10'b0010010000: data <= 11'h7ff; 
        10'b0010010001: data <= 11'h7ff; 
        10'b0010010010: data <= 11'h7ff; 
        10'b0010010011: data <= 11'h7fd; 
        10'b0010010100: data <= 11'h7ff; 
        10'b0010010101: data <= 11'h001; 
        10'b0010010110: data <= 11'h7fd; 
        10'b0010010111: data <= 11'h004; 
        10'b0010011000: data <= 11'h007; 
        10'b0010011001: data <= 11'h006; 
        10'b0010011010: data <= 11'h006; 
        10'b0010011011: data <= 11'h003; 
        10'b0010011100: data <= 11'h002; 
        10'b0010011101: data <= 11'h006; 
        10'b0010011110: data <= 11'h000; 
        10'b0010011111: data <= 11'h000; 
        10'b0010100000: data <= 11'h002; 
        10'b0010100001: data <= 11'h001; 
        10'b0010100010: data <= 11'h7fd; 
        10'b0010100011: data <= 11'h7fd; 
        10'b0010100100: data <= 11'h7fe; 
        10'b0010100101: data <= 11'h001; 
        10'b0010100110: data <= 11'h7ff; 
        10'b0010100111: data <= 11'h000; 
        10'b0010101000: data <= 11'h7ff; 
        10'b0010101001: data <= 11'h7ff; 
        10'b0010101010: data <= 11'h7fe; 
        10'b0010101011: data <= 11'h7fe; 
        10'b0010101100: data <= 11'h7fe; 
        10'b0010101101: data <= 11'h7fe; 
        10'b0010101110: data <= 11'h7fd; 
        10'b0010101111: data <= 11'h7fd; 
        10'b0010110000: data <= 11'h000; 
        10'b0010110001: data <= 11'h001; 
        10'b0010110010: data <= 11'h000; 
        10'b0010110011: data <= 11'h002; 
        10'b0010110100: data <= 11'h003; 
        10'b0010110101: data <= 11'h002; 
        10'b0010110110: data <= 11'h003; 
        10'b0010110111: data <= 11'h006; 
        10'b0010111000: data <= 11'h003; 
        10'b0010111001: data <= 11'h003; 
        10'b0010111010: data <= 11'h001; 
        10'b0010111011: data <= 11'h004; 
        10'b0010111100: data <= 11'h001; 
        10'b0010111101: data <= 11'h002; 
        10'b0010111110: data <= 11'h002; 
        10'b0010111111: data <= 11'h002; 
        10'b0011000000: data <= 11'h002; 
        10'b0011000001: data <= 11'h001; 
        10'b0011000010: data <= 11'h7ff; 
        10'b0011000011: data <= 11'h000; 
        10'b0011000100: data <= 11'h000; 
        10'b0011000101: data <= 11'h7ff; 
        10'b0011000110: data <= 11'h7fe; 
        10'b0011000111: data <= 11'h7ff; 
        10'b0011001000: data <= 11'h7fe; 
        10'b0011001001: data <= 11'h7ff; 
        10'b0011001010: data <= 11'h7fe; 
        10'b0011001011: data <= 11'h000; 
        10'b0011001100: data <= 11'h002; 
        10'b0011001101: data <= 11'h001; 
        10'b0011001110: data <= 11'h001; 
        10'b0011001111: data <= 11'h7ff; 
        10'b0011010000: data <= 11'h7fd; 
        10'b0011010001: data <= 11'h7fe; 
        10'b0011010010: data <= 11'h7fd; 
        10'b0011010011: data <= 11'h002; 
        10'b0011010100: data <= 11'h002; 
        10'b0011010101: data <= 11'h000; 
        10'b0011010110: data <= 11'h002; 
        10'b0011010111: data <= 11'h7fe; 
        10'b0011011000: data <= 11'h002; 
        10'b0011011001: data <= 11'h004; 
        10'b0011011010: data <= 11'h001; 
        10'b0011011011: data <= 11'h008; 
        10'b0011011100: data <= 11'h005; 
        10'b0011011101: data <= 11'h000; 
        10'b0011011110: data <= 11'h000; 
        10'b0011011111: data <= 11'h000; 
        10'b0011100000: data <= 11'h000; 
        10'b0011100001: data <= 11'h000; 
        10'b0011100010: data <= 11'h000; 
        10'b0011100011: data <= 11'h7ff; 
        10'b0011100100: data <= 11'h000; 
        10'b0011100101: data <= 11'h7ff; 
        10'b0011100110: data <= 11'h003; 
        10'b0011100111: data <= 11'h002; 
        10'b0011101000: data <= 11'h001; 
        10'b0011101001: data <= 11'h005; 
        10'b0011101010: data <= 11'h000; 
        10'b0011101011: data <= 11'h000; 
        10'b0011101100: data <= 11'h004; 
        10'b0011101101: data <= 11'h005; 
        10'b0011101110: data <= 11'h7fc; 
        10'b0011101111: data <= 11'h7fd; 
        10'b0011110000: data <= 11'h003; 
        10'b0011110001: data <= 11'h7fe; 
        10'b0011110010: data <= 11'h001; 
        10'b0011110011: data <= 11'h002; 
        10'b0011110100: data <= 11'h002; 
        10'b0011110101: data <= 11'h005; 
        10'b0011110110: data <= 11'h003; 
        10'b0011110111: data <= 11'h006; 
        10'b0011111000: data <= 11'h005; 
        10'b0011111001: data <= 11'h7ff; 
        10'b0011111010: data <= 11'h000; 
        10'b0011111011: data <= 11'h001; 
        10'b0011111100: data <= 11'h000; 
        10'b0011111101: data <= 11'h000; 
        10'b0011111110: data <= 11'h7ff; 
        10'b0011111111: data <= 11'h7ff; 
        10'b0100000000: data <= 11'h7ff; 
        10'b0100000001: data <= 11'h003; 
        10'b0100000010: data <= 11'h002; 
        10'b0100000011: data <= 11'h005; 
        10'b0100000100: data <= 11'h006; 
        10'b0100000101: data <= 11'h005; 
        10'b0100000110: data <= 11'h003; 
        10'b0100000111: data <= 11'h006; 
        10'b0100001000: data <= 11'h002; 
        10'b0100001001: data <= 11'h002; 
        10'b0100001010: data <= 11'h7f9; 
        10'b0100001011: data <= 11'h7f6; 
        10'b0100001100: data <= 11'h7fd; 
        10'b0100001101: data <= 11'h001; 
        10'b0100001110: data <= 11'h001; 
        10'b0100001111: data <= 11'h002; 
        10'b0100010000: data <= 11'h003; 
        10'b0100010001: data <= 11'h002; 
        10'b0100010010: data <= 11'h005; 
        10'b0100010011: data <= 11'h005; 
        10'b0100010100: data <= 11'h7ff; 
        10'b0100010101: data <= 11'h7ff; 
        10'b0100010110: data <= 11'h001; 
        10'b0100010111: data <= 11'h7fe; 
        10'b0100011000: data <= 11'h7ff; 
        10'b0100011001: data <= 11'h000; 
        10'b0100011010: data <= 11'h7ff; 
        10'b0100011011: data <= 11'h000; 
        10'b0100011100: data <= 11'h001; 
        10'b0100011101: data <= 11'h004; 
        10'b0100011110: data <= 11'h004; 
        10'b0100011111: data <= 11'h007; 
        10'b0100100000: data <= 11'h005; 
        10'b0100100001: data <= 11'h006; 
        10'b0100100010: data <= 11'h009; 
        10'b0100100011: data <= 11'h004; 
        10'b0100100100: data <= 11'h004; 
        10'b0100100101: data <= 11'h004; 
        10'b0100100110: data <= 11'h7ff; 
        10'b0100100111: data <= 11'h7f7; 
        10'b0100101000: data <= 11'h7f8; 
        10'b0100101001: data <= 11'h7fe; 
        10'b0100101010: data <= 11'h003; 
        10'b0100101011: data <= 11'h003; 
        10'b0100101100: data <= 11'h003; 
        10'b0100101101: data <= 11'h006; 
        10'b0100101110: data <= 11'h007; 
        10'b0100101111: data <= 11'h006; 
        10'b0100110000: data <= 11'h000; 
        10'b0100110001: data <= 11'h000; 
        10'b0100110010: data <= 11'h7ff; 
        10'b0100110011: data <= 11'h7ff; 
        10'b0100110100: data <= 11'h7ff; 
        10'b0100110101: data <= 11'h000; 
        10'b0100110110: data <= 11'h000; 
        10'b0100110111: data <= 11'h7fe; 
        10'b0100111000: data <= 11'h002; 
        10'b0100111001: data <= 11'h004; 
        10'b0100111010: data <= 11'h008; 
        10'b0100111011: data <= 11'h00b; 
        10'b0100111100: data <= 11'h008; 
        10'b0100111101: data <= 11'h00a; 
        10'b0100111110: data <= 11'h007; 
        10'b0100111111: data <= 11'h003; 
        10'b0101000000: data <= 11'h004; 
        10'b0101000001: data <= 11'h00a; 
        10'b0101000010: data <= 11'h00d; 
        10'b0101000011: data <= 11'h7fe; 
        10'b0101000100: data <= 11'h7f8; 
        10'b0101000101: data <= 11'h7fd; 
        10'b0101000110: data <= 11'h7fe; 
        10'b0101000111: data <= 11'h001; 
        10'b0101001000: data <= 11'h006; 
        10'b0101001001: data <= 11'h007; 
        10'b0101001010: data <= 11'h009; 
        10'b0101001011: data <= 11'h009; 
        10'b0101001100: data <= 11'h006; 
        10'b0101001101: data <= 11'h001; 
        10'b0101001110: data <= 11'h001; 
        10'b0101001111: data <= 11'h000; 
        10'b0101010000: data <= 11'h7ff; 
        10'b0101010001: data <= 11'h000; 
        10'b0101010010: data <= 11'h7ff; 
        10'b0101010011: data <= 11'h000; 
        10'b0101010100: data <= 11'h000; 
        10'b0101010101: data <= 11'h005; 
        10'b0101010110: data <= 11'h004; 
        10'b0101010111: data <= 11'h006; 
        10'b0101011000: data <= 11'h006; 
        10'b0101011001: data <= 11'h008; 
        10'b0101011010: data <= 11'h001; 
        10'b0101011011: data <= 11'h002; 
        10'b0101011100: data <= 11'h001; 
        10'b0101011101: data <= 11'h00d; 
        10'b0101011110: data <= 11'h00d; 
        10'b0101011111: data <= 11'h003; 
        10'b0101100000: data <= 11'h000; 
        10'b0101100001: data <= 11'h7ff; 
        10'b0101100010: data <= 11'h7ff; 
        10'b0101100011: data <= 11'h003; 
        10'b0101100100: data <= 11'h005; 
        10'b0101100101: data <= 11'h009; 
        10'b0101100110: data <= 11'h00b; 
        10'b0101100111: data <= 11'h009; 
        10'b0101101000: data <= 11'h006; 
        10'b0101101001: data <= 11'h002; 
        10'b0101101010: data <= 11'h001; 
        10'b0101101011: data <= 11'h7fe; 
        10'b0101101100: data <= 11'h7fe; 
        10'b0101101101: data <= 11'h7ff; 
        10'b0101101110: data <= 11'h000; 
        10'b0101101111: data <= 11'h7fe; 
        10'b0101110000: data <= 11'h7ff; 
        10'b0101110001: data <= 11'h000; 
        10'b0101110010: data <= 11'h7ff; 
        10'b0101110011: data <= 11'h7ff; 
        10'b0101110100: data <= 11'h001; 
        10'b0101110101: data <= 11'h7ff; 
        10'b0101110110: data <= 11'h7fd; 
        10'b0101110111: data <= 11'h001; 
        10'b0101111000: data <= 11'h005; 
        10'b0101111001: data <= 11'h00c; 
        10'b0101111010: data <= 11'h004; 
        10'b0101111011: data <= 11'h009; 
        10'b0101111100: data <= 11'h003; 
        10'b0101111101: data <= 11'h7fe; 
        10'b0101111110: data <= 11'h000; 
        10'b0101111111: data <= 11'h000; 
        10'b0110000000: data <= 11'h004; 
        10'b0110000001: data <= 11'h003; 
        10'b0110000010: data <= 11'h002; 
        10'b0110000011: data <= 11'h003; 
        10'b0110000100: data <= 11'h001; 
        10'b0110000101: data <= 11'h000; 
        10'b0110000110: data <= 11'h000; 
        10'b0110000111: data <= 11'h000; 
        10'b0110001000: data <= 11'h7ff; 
        10'b0110001001: data <= 11'h7fe; 
        10'b0110001010: data <= 11'h000; 
        10'b0110001011: data <= 11'h7ff; 
        10'b0110001100: data <= 11'h7fe; 
        10'b0110001101: data <= 11'h7fd; 
        10'b0110001110: data <= 11'h7fa; 
        10'b0110001111: data <= 11'h7f8; 
        10'b0110010000: data <= 11'h7f7; 
        10'b0110010001: data <= 11'h7f9; 
        10'b0110010010: data <= 11'h7ff; 
        10'b0110010011: data <= 11'h005; 
        10'b0110010100: data <= 11'h005; 
        10'b0110010101: data <= 11'h00a; 
        10'b0110010110: data <= 11'h008; 
        10'b0110010111: data <= 11'h005; 
        10'b0110011000: data <= 11'h7ff; 
        10'b0110011001: data <= 11'h001; 
        10'b0110011010: data <= 11'h7ff; 
        10'b0110011011: data <= 11'h7fd; 
        10'b0110011100: data <= 11'h7fb; 
        10'b0110011101: data <= 11'h7fb; 
        10'b0110011110: data <= 11'h7fc; 
        10'b0110011111: data <= 11'h7fb; 
        10'b0110100000: data <= 11'h7fe; 
        10'b0110100001: data <= 11'h000; 
        10'b0110100010: data <= 11'h7fe; 
        10'b0110100011: data <= 11'h000; 
        10'b0110100100: data <= 11'h000; 
        10'b0110100101: data <= 11'h7ff; 
        10'b0110100110: data <= 11'h7ff; 
        10'b0110100111: data <= 11'h7ff; 
        10'b0110101000: data <= 11'h7fe; 
        10'b0110101001: data <= 11'h7fd; 
        10'b0110101010: data <= 11'h7f8; 
        10'b0110101011: data <= 11'h7f7; 
        10'b0110101100: data <= 11'h7f7; 
        10'b0110101101: data <= 11'h7fe; 
        10'b0110101110: data <= 11'h000; 
        10'b0110101111: data <= 11'h000; 
        10'b0110110000: data <= 11'h007; 
        10'b0110110001: data <= 11'h008; 
        10'b0110110010: data <= 11'h007; 
        10'b0110110011: data <= 11'h004; 
        10'b0110110100: data <= 11'h7fe; 
        10'b0110110101: data <= 11'h7fe; 
        10'b0110110110: data <= 11'h7ff; 
        10'b0110110111: data <= 11'h7f9; 
        10'b0110111000: data <= 11'h7f7; 
        10'b0110111001: data <= 11'h7f9; 
        10'b0110111010: data <= 11'h7fc; 
        10'b0110111011: data <= 11'h7fc; 
        10'b0110111100: data <= 11'h7fd; 
        10'b0110111101: data <= 11'h7ff; 
        10'b0110111110: data <= 11'h7fe; 
        10'b0110111111: data <= 11'h000; 
        10'b0111000000: data <= 11'h7ff; 
        10'b0111000001: data <= 11'h7fe; 
        10'b0111000010: data <= 11'h7ff; 
        10'b0111000011: data <= 11'h7ff; 
        10'b0111000100: data <= 11'h7fd; 
        10'b0111000101: data <= 11'h7fb; 
        10'b0111000110: data <= 11'h7f8; 
        10'b0111000111: data <= 11'h7fb; 
        10'b0111001000: data <= 11'h003; 
        10'b0111001001: data <= 11'h003; 
        10'b0111001010: data <= 11'h001; 
        10'b0111001011: data <= 11'h003; 
        10'b0111001100: data <= 11'h006; 
        10'b0111001101: data <= 11'h006; 
        10'b0111001110: data <= 11'h002; 
        10'b0111001111: data <= 11'h003; 
        10'b0111010000: data <= 11'h001; 
        10'b0111010001: data <= 11'h7fd; 
        10'b0111010010: data <= 11'h7fa; 
        10'b0111010011: data <= 11'h7f8; 
        10'b0111010100: data <= 11'h7f8; 
        10'b0111010101: data <= 11'h7f8; 
        10'b0111010110: data <= 11'h7fa; 
        10'b0111010111: data <= 11'h7fe; 
        10'b0111011000: data <= 11'h7fd; 
        10'b0111011001: data <= 11'h7ff; 
        10'b0111011010: data <= 11'h7ff; 
        10'b0111011011: data <= 11'h7fe; 
        10'b0111011100: data <= 11'h000; 
        10'b0111011101: data <= 11'h000; 
        10'b0111011110: data <= 11'h7ff; 
        10'b0111011111: data <= 11'h7fe; 
        10'b0111100000: data <= 11'h7fe; 
        10'b0111100001: data <= 11'h7fb; 
        10'b0111100010: data <= 11'h7f9; 
        10'b0111100011: data <= 11'h001; 
        10'b0111100100: data <= 11'h007; 
        10'b0111100101: data <= 11'h008; 
        10'b0111100110: data <= 11'h003; 
        10'b0111100111: data <= 11'h006; 
        10'b0111101000: data <= 11'h00a; 
        10'b0111101001: data <= 11'h006; 
        10'b0111101010: data <= 11'h001; 
        10'b0111101011: data <= 11'h7fe; 
        10'b0111101100: data <= 11'h001; 
        10'b0111101101: data <= 11'h7fd; 
        10'b0111101110: data <= 11'h7f8; 
        10'b0111101111: data <= 11'h7fc; 
        10'b0111110000: data <= 11'h7fc; 
        10'b0111110001: data <= 11'h7fb; 
        10'b0111110010: data <= 11'h7fc; 
        10'b0111110011: data <= 11'h7fd; 
        10'b0111110100: data <= 11'h7ff; 
        10'b0111110101: data <= 11'h7fe; 
        10'b0111110110: data <= 11'h000; 
        10'b0111110111: data <= 11'h7ff; 
        10'b0111111000: data <= 11'h7ff; 
        10'b0111111001: data <= 11'h000; 
        10'b0111111010: data <= 11'h7fe; 
        10'b0111111011: data <= 11'h7fe; 
        10'b0111111100: data <= 11'h7fd; 
        10'b0111111101: data <= 11'h7fd; 
        10'b0111111110: data <= 11'h7fe; 
        10'b0111111111: data <= 11'h002; 
        10'b1000000000: data <= 11'h005; 
        10'b1000000001: data <= 11'h00a; 
        10'b1000000010: data <= 11'h007; 
        10'b1000000011: data <= 11'h009; 
        10'b1000000100: data <= 11'h006; 
        10'b1000000101: data <= 11'h003; 
        10'b1000000110: data <= 11'h7fc; 
        10'b1000000111: data <= 11'h7ff; 
        10'b1000001000: data <= 11'h7fe; 
        10'b1000001001: data <= 11'h7fa; 
        10'b1000001010: data <= 11'h7fe; 
        10'b1000001011: data <= 11'h7ff; 
        10'b1000001100: data <= 11'h000; 
        10'b1000001101: data <= 11'h7fd; 
        10'b1000001110: data <= 11'h7ff; 
        10'b1000001111: data <= 11'h7fd; 
        10'b1000010000: data <= 11'h7fc; 
        10'b1000010001: data <= 11'h7fe; 
        10'b1000010010: data <= 11'h000; 
        10'b1000010011: data <= 11'h000; 
        10'b1000010100: data <= 11'h7ff; 
        10'b1000010101: data <= 11'h7ff; 
        10'b1000010110: data <= 11'h000; 
        10'b1000010111: data <= 11'h7fd; 
        10'b1000011000: data <= 11'h7fd; 
        10'b1000011001: data <= 11'h7ff; 
        10'b1000011010: data <= 11'h001; 
        10'b1000011011: data <= 11'h003; 
        10'b1000011100: data <= 11'h003; 
        10'b1000011101: data <= 11'h007; 
        10'b1000011110: data <= 11'h003; 
        10'b1000011111: data <= 11'h000; 
        10'b1000100000: data <= 11'h002; 
        10'b1000100001: data <= 11'h7fc; 
        10'b1000100010: data <= 11'h7fb; 
        10'b1000100011: data <= 11'h7fe; 
        10'b1000100100: data <= 11'h7fe; 
        10'b1000100101: data <= 11'h7fe; 
        10'b1000100110: data <= 11'h002; 
        10'b1000100111: data <= 11'h000; 
        10'b1000101000: data <= 11'h002; 
        10'b1000101001: data <= 11'h000; 
        10'b1000101010: data <= 11'h001; 
        10'b1000101011: data <= 11'h7ff; 
        10'b1000101100: data <= 11'h7fd; 
        10'b1000101101: data <= 11'h7fe; 
        10'b1000101110: data <= 11'h7fe; 
        10'b1000101111: data <= 11'h000; 
        10'b1000110000: data <= 11'h7ff; 
        10'b1000110001: data <= 11'h000; 
        10'b1000110010: data <= 11'h7ff; 
        10'b1000110011: data <= 11'h7fe; 
        10'b1000110100: data <= 11'h7fc; 
        10'b1000110101: data <= 11'h7ff; 
        10'b1000110110: data <= 11'h001; 
        10'b1000110111: data <= 11'h006; 
        10'b1000111000: data <= 11'h002; 
        10'b1000111001: data <= 11'h7ff; 
        10'b1000111010: data <= 11'h000; 
        10'b1000111011: data <= 11'h7fb; 
        10'b1000111100: data <= 11'h000; 
        10'b1000111101: data <= 11'h000; 
        10'b1000111110: data <= 11'h7fb; 
        10'b1000111111: data <= 11'h7ff; 
        10'b1001000000: data <= 11'h7fb; 
        10'b1001000001: data <= 11'h7fe; 
        10'b1001000010: data <= 11'h001; 
        10'b1001000011: data <= 11'h001; 
        10'b1001000100: data <= 11'h002; 
        10'b1001000101: data <= 11'h003; 
        10'b1001000110: data <= 11'h003; 
        10'b1001000111: data <= 11'h7ff; 
        10'b1001001000: data <= 11'h7fe; 
        10'b1001001001: data <= 11'h7fe; 
        10'b1001001010: data <= 11'h7ff; 
        10'b1001001011: data <= 11'h7ff; 
        10'b1001001100: data <= 11'h000; 
        10'b1001001101: data <= 11'h7ff; 
        10'b1001001110: data <= 11'h000; 
        10'b1001001111: data <= 11'h7fd; 
        10'b1001010000: data <= 11'h7fb; 
        10'b1001010001: data <= 11'h000; 
        10'b1001010010: data <= 11'h002; 
        10'b1001010011: data <= 11'h005; 
        10'b1001010100: data <= 11'h001; 
        10'b1001010101: data <= 11'h002; 
        10'b1001010110: data <= 11'h000; 
        10'b1001010111: data <= 11'h7fd; 
        10'b1001011000: data <= 11'h7fe; 
        10'b1001011001: data <= 11'h001; 
        10'b1001011010: data <= 11'h000; 
        10'b1001011011: data <= 11'h7ff; 
        10'b1001011100: data <= 11'h7fc; 
        10'b1001011101: data <= 11'h7fe; 
        10'b1001011110: data <= 11'h7ff; 
        10'b1001011111: data <= 11'h000; 
        10'b1001100000: data <= 11'h000; 
        10'b1001100001: data <= 11'h001; 
        10'b1001100010: data <= 11'h001; 
        10'b1001100011: data <= 11'h7ff; 
        10'b1001100100: data <= 11'h7ff; 
        10'b1001100101: data <= 11'h000; 
        10'b1001100110: data <= 11'h000; 
        10'b1001100111: data <= 11'h7ff; 
        10'b1001101000: data <= 11'h000; 
        10'b1001101001: data <= 11'h7fe; 
        10'b1001101010: data <= 11'h7ff; 
        10'b1001101011: data <= 11'h7fe; 
        10'b1001101100: data <= 11'h7fc; 
        10'b1001101101: data <= 11'h7fa; 
        10'b1001101110: data <= 11'h001; 
        10'b1001101111: data <= 11'h001; 
        10'b1001110000: data <= 11'h000; 
        10'b1001110001: data <= 11'h7fe; 
        10'b1001110010: data <= 11'h001; 
        10'b1001110011: data <= 11'h000; 
        10'b1001110100: data <= 11'h007; 
        10'b1001110101: data <= 11'h007; 
        10'b1001110110: data <= 11'h005; 
        10'b1001110111: data <= 11'h004; 
        10'b1001111000: data <= 11'h000; 
        10'b1001111001: data <= 11'h000; 
        10'b1001111010: data <= 11'h002; 
        10'b1001111011: data <= 11'h7fe; 
        10'b1001111100: data <= 11'h7fe; 
        10'b1001111101: data <= 11'h001; 
        10'b1001111110: data <= 11'h000; 
        10'b1001111111: data <= 11'h7ff; 
        10'b1010000000: data <= 11'h000; 
        10'b1010000001: data <= 11'h000; 
        10'b1010000010: data <= 11'h000; 
        10'b1010000011: data <= 11'h7ff; 
        10'b1010000100: data <= 11'h7ff; 
        10'b1010000101: data <= 11'h000; 
        10'b1010000110: data <= 11'h7ff; 
        10'b1010000111: data <= 11'h7fe; 
        10'b1010001000: data <= 11'h7fc; 
        10'b1010001001: data <= 11'h7f7; 
        10'b1010001010: data <= 11'h7f9; 
        10'b1010001011: data <= 11'h7fc; 
        10'b1010001100: data <= 11'h001; 
        10'b1010001101: data <= 11'h001; 
        10'b1010001110: data <= 11'h003; 
        10'b1010001111: data <= 11'h004; 
        10'b1010010000: data <= 11'h008; 
        10'b1010010001: data <= 11'h00b; 
        10'b1010010010: data <= 11'h00a; 
        10'b1010010011: data <= 11'h008; 
        10'b1010010100: data <= 11'h006; 
        10'b1010010101: data <= 11'h004; 
        10'b1010010110: data <= 11'h004; 
        10'b1010010111: data <= 11'h004; 
        10'b1010011000: data <= 11'h003; 
        10'b1010011001: data <= 11'h001; 
        10'b1010011010: data <= 11'h000; 
        10'b1010011011: data <= 11'h7ff; 
        10'b1010011100: data <= 11'h7fe; 
        10'b1010011101: data <= 11'h000; 
        10'b1010011110: data <= 11'h7fe; 
        10'b1010011111: data <= 11'h000; 
        10'b1010100000: data <= 11'h000; 
        10'b1010100001: data <= 11'h000; 
        10'b1010100010: data <= 11'h000; 
        10'b1010100011: data <= 11'h7fe; 
        10'b1010100100: data <= 11'h7fe; 
        10'b1010100101: data <= 11'h7fa; 
        10'b1010100110: data <= 11'h7f8; 
        10'b1010100111: data <= 11'h7f9; 
        10'b1010101000: data <= 11'h000; 
        10'b1010101001: data <= 11'h002; 
        10'b1010101010: data <= 11'h7ff; 
        10'b1010101011: data <= 11'h003; 
        10'b1010101100: data <= 11'h002; 
        10'b1010101101: data <= 11'h001; 
        10'b1010101110: data <= 11'h004; 
        10'b1010101111: data <= 11'h008; 
        10'b1010110000: data <= 11'h009; 
        10'b1010110001: data <= 11'h006; 
        10'b1010110010: data <= 11'h008; 
        10'b1010110011: data <= 11'h008; 
        10'b1010110100: data <= 11'h002; 
        10'b1010110101: data <= 11'h000; 
        10'b1010110110: data <= 11'h7fe; 
        10'b1010110111: data <= 11'h000; 
        10'b1010111000: data <= 11'h7ff; 
        10'b1010111001: data <= 11'h7ff; 
        10'b1010111010: data <= 11'h000; 
        10'b1010111011: data <= 11'h000; 
        10'b1010111100: data <= 11'h000; 
        10'b1010111101: data <= 11'h000; 
        10'b1010111110: data <= 11'h000; 
        10'b1010111111: data <= 11'h7fe; 
        10'b1011000000: data <= 11'h7ff; 
        10'b1011000001: data <= 11'h7fe; 
        10'b1011000010: data <= 11'h7fd; 
        10'b1011000011: data <= 11'h7fc; 
        10'b1011000100: data <= 11'h7fc; 
        10'b1011000101: data <= 11'h7fc; 
        10'b1011000110: data <= 11'h7fe; 
        10'b1011000111: data <= 11'h7fd; 
        10'b1011001000: data <= 11'h7fe; 
        10'b1011001001: data <= 11'h7fe; 
        10'b1011001010: data <= 11'h000; 
        10'b1011001011: data <= 11'h003; 
        10'b1011001100: data <= 11'h002; 
        10'b1011001101: data <= 11'h003; 
        10'b1011001110: data <= 11'h003; 
        10'b1011001111: data <= 11'h000; 
        10'b1011010000: data <= 11'h7ff; 
        10'b1011010001: data <= 11'h000; 
        10'b1011010010: data <= 11'h7fe; 
        10'b1011010011: data <= 11'h7fe; 
        10'b1011010100: data <= 11'h000; 
        10'b1011010101: data <= 11'h7ff; 
        10'b1011010110: data <= 11'h7ff; 
        10'b1011010111: data <= 11'h7ff; 
        10'b1011011000: data <= 11'h000; 
        10'b1011011001: data <= 11'h000; 
        10'b1011011010: data <= 11'h7ff; 
        10'b1011011011: data <= 11'h7ff; 
        10'b1011011100: data <= 11'h7fe; 
        10'b1011011101: data <= 11'h7fe; 
        10'b1011011110: data <= 11'h7fe; 
        10'b1011011111: data <= 11'h7ff; 
        10'b1011100000: data <= 11'h7fe; 
        10'b1011100001: data <= 11'h7fe; 
        10'b1011100010: data <= 11'h7fe; 
        10'b1011100011: data <= 11'h7ff; 
        10'b1011100100: data <= 11'h7ff; 
        10'b1011100101: data <= 11'h7ff; 
        10'b1011100110: data <= 11'h7fe; 
        10'b1011100111: data <= 11'h7ff; 
        10'b1011101000: data <= 11'h7fe; 
        10'b1011101001: data <= 11'h7fe; 
        10'b1011101010: data <= 11'h7fe; 
        10'b1011101011: data <= 11'h7ff; 
        10'b1011101100: data <= 11'h7ff; 
        10'b1011101101: data <= 11'h000; 
        10'b1011101110: data <= 11'h7ff; 
        10'b1011101111: data <= 11'h000; 
        10'b1011110000: data <= 11'h000; 
        10'b1011110001: data <= 11'h7fe; 
        10'b1011110010: data <= 11'h7ff; 
        10'b1011110011: data <= 11'h7ff; 
        10'b1011110100: data <= 11'h000; 
        10'b1011110101: data <= 11'h7ff; 
        10'b1011110110: data <= 11'h7ff; 
        10'b1011110111: data <= 11'h7ff; 
        10'b1011111000: data <= 11'h000; 
        10'b1011111001: data <= 11'h7fe; 
        10'b1011111010: data <= 11'h000; 
        10'b1011111011: data <= 11'h7ff; 
        10'b1011111100: data <= 11'h000; 
        10'b1011111101: data <= 11'h7ff; 
        10'b1011111110: data <= 11'h7fe; 
        10'b1011111111: data <= 11'h000; 
        10'b1100000000: data <= 11'h7ff; 
        10'b1100000001: data <= 11'h7fe; 
        10'b1100000010: data <= 11'h7ff; 
        10'b1100000011: data <= 11'h000; 
        10'b1100000100: data <= 11'h7ff; 
        10'b1100000101: data <= 11'h000; 
        10'b1100000110: data <= 11'h000; 
        10'b1100000111: data <= 11'h000; 
        10'b1100001000: data <= 11'h000; 
        10'b1100001001: data <= 11'h7ff; 
        10'b1100001010: data <= 11'h000; 
        10'b1100001011: data <= 11'h7ff; 
        10'b1100001100: data <= 11'h7ff; 
        10'b1100001101: data <= 11'h000; 
        10'b1100001110: data <= 11'h7fe; 
        10'b1100001111: data <= 11'h7ff; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 6) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 12'hffe; 
        10'b0000000001: data <= 12'hfff; 
        10'b0000000010: data <= 12'hffe; 
        10'b0000000011: data <= 12'hfff; 
        10'b0000000100: data <= 12'hfff; 
        10'b0000000101: data <= 12'h000; 
        10'b0000000110: data <= 12'hffc; 
        10'b0000000111: data <= 12'hfff; 
        10'b0000001000: data <= 12'hffe; 
        10'b0000001001: data <= 12'hffe; 
        10'b0000001010: data <= 12'hffd; 
        10'b0000001011: data <= 12'h000; 
        10'b0000001100: data <= 12'hfff; 
        10'b0000001101: data <= 12'h000; 
        10'b0000001110: data <= 12'hffd; 
        10'b0000001111: data <= 12'h000; 
        10'b0000010000: data <= 12'hfff; 
        10'b0000010001: data <= 12'hffd; 
        10'b0000010010: data <= 12'h000; 
        10'b0000010011: data <= 12'hfff; 
        10'b0000010100: data <= 12'hffe; 
        10'b0000010101: data <= 12'hffe; 
        10'b0000010110: data <= 12'hffe; 
        10'b0000010111: data <= 12'h001; 
        10'b0000011000: data <= 12'h000; 
        10'b0000011001: data <= 12'hffe; 
        10'b0000011010: data <= 12'hffd; 
        10'b0000011011: data <= 12'hffe; 
        10'b0000011100: data <= 12'hffe; 
        10'b0000011101: data <= 12'hffc; 
        10'b0000011110: data <= 12'h001; 
        10'b0000011111: data <= 12'h000; 
        10'b0000100000: data <= 12'hffd; 
        10'b0000100001: data <= 12'hffd; 
        10'b0000100010: data <= 12'hffc; 
        10'b0000100011: data <= 12'hffd; 
        10'b0000100100: data <= 12'h000; 
        10'b0000100101: data <= 12'hfff; 
        10'b0000100110: data <= 12'hfff; 
        10'b0000100111: data <= 12'hffc; 
        10'b0000101000: data <= 12'h000; 
        10'b0000101001: data <= 12'hfff; 
        10'b0000101010: data <= 12'hffe; 
        10'b0000101011: data <= 12'hffe; 
        10'b0000101100: data <= 12'hfff; 
        10'b0000101101: data <= 12'hfff; 
        10'b0000101110: data <= 12'hffd; 
        10'b0000101111: data <= 12'hfff; 
        10'b0000110000: data <= 12'h000; 
        10'b0000110001: data <= 12'hffd; 
        10'b0000110010: data <= 12'hfff; 
        10'b0000110011: data <= 12'hffd; 
        10'b0000110100: data <= 12'h000; 
        10'b0000110101: data <= 12'h001; 
        10'b0000110110: data <= 12'hffe; 
        10'b0000110111: data <= 12'hffd; 
        10'b0000111000: data <= 12'hffd; 
        10'b0000111001: data <= 12'h000; 
        10'b0000111010: data <= 12'hfff; 
        10'b0000111011: data <= 12'hffe; 
        10'b0000111100: data <= 12'hffd; 
        10'b0000111101: data <= 12'hffc; 
        10'b0000111110: data <= 12'hfff; 
        10'b0000111111: data <= 12'hffc; 
        10'b0001000000: data <= 12'h001; 
        10'b0001000001: data <= 12'hffc; 
        10'b0001000010: data <= 12'hffc; 
        10'b0001000011: data <= 12'hfff; 
        10'b0001000100: data <= 12'hfff; 
        10'b0001000101: data <= 12'hffc; 
        10'b0001000110: data <= 12'hfff; 
        10'b0001000111: data <= 12'hfff; 
        10'b0001001000: data <= 12'hffc; 
        10'b0001001001: data <= 12'hffe; 
        10'b0001001010: data <= 12'hffe; 
        10'b0001001011: data <= 12'hfff; 
        10'b0001001100: data <= 12'h000; 
        10'b0001001101: data <= 12'h000; 
        10'b0001001110: data <= 12'hfff; 
        10'b0001001111: data <= 12'hffe; 
        10'b0001010000: data <= 12'h000; 
        10'b0001010001: data <= 12'hffe; 
        10'b0001010010: data <= 12'hfff; 
        10'b0001010011: data <= 12'h000; 
        10'b0001010100: data <= 12'hffd; 
        10'b0001010101: data <= 12'hffe; 
        10'b0001010110: data <= 12'hffe; 
        10'b0001010111: data <= 12'hffd; 
        10'b0001011000: data <= 12'h001; 
        10'b0001011001: data <= 12'hffd; 
        10'b0001011010: data <= 12'hffd; 
        10'b0001011011: data <= 12'hffe; 
        10'b0001011100: data <= 12'hffc; 
        10'b0001011101: data <= 12'hfff; 
        10'b0001011110: data <= 12'hffd; 
        10'b0001011111: data <= 12'hffb; 
        10'b0001100000: data <= 12'hffa; 
        10'b0001100001: data <= 12'hff9; 
        10'b0001100010: data <= 12'hffa; 
        10'b0001100011: data <= 12'hffd; 
        10'b0001100100: data <= 12'hffa; 
        10'b0001100101: data <= 12'hffc; 
        10'b0001100110: data <= 12'hffd; 
        10'b0001100111: data <= 12'hffe; 
        10'b0001101000: data <= 12'hffc; 
        10'b0001101001: data <= 12'h000; 
        10'b0001101010: data <= 12'hffe; 
        10'b0001101011: data <= 12'h000; 
        10'b0001101100: data <= 12'hffe; 
        10'b0001101101: data <= 12'hfff; 
        10'b0001101110: data <= 12'hfff; 
        10'b0001101111: data <= 12'hffd; 
        10'b0001110000: data <= 12'hfff; 
        10'b0001110001: data <= 12'h000; 
        10'b0001110010: data <= 12'hffe; 
        10'b0001110011: data <= 12'hffd; 
        10'b0001110100: data <= 12'h000; 
        10'b0001110101: data <= 12'h000; 
        10'b0001110110: data <= 12'hfff; 
        10'b0001110111: data <= 12'hffd; 
        10'b0001111000: data <= 12'hffd; 
        10'b0001111001: data <= 12'hffe; 
        10'b0001111010: data <= 12'hffe; 
        10'b0001111011: data <= 12'hfff; 
        10'b0001111100: data <= 12'h005; 
        10'b0001111101: data <= 12'h003; 
        10'b0001111110: data <= 12'h00b; 
        10'b0001111111: data <= 12'h008; 
        10'b0010000000: data <= 12'h004; 
        10'b0010000001: data <= 12'h002; 
        10'b0010000010: data <= 12'h003; 
        10'b0010000011: data <= 12'hffd; 
        10'b0010000100: data <= 12'hffd; 
        10'b0010000101: data <= 12'hffe; 
        10'b0010000110: data <= 12'hffb; 
        10'b0010000111: data <= 12'hffc; 
        10'b0010001000: data <= 12'h000; 
        10'b0010001001: data <= 12'h000; 
        10'b0010001010: data <= 12'hffe; 
        10'b0010001011: data <= 12'hfff; 
        10'b0010001100: data <= 12'hfff; 
        10'b0010001101: data <= 12'hfff; 
        10'b0010001110: data <= 12'h000; 
        10'b0010001111: data <= 12'h000; 
        10'b0010010000: data <= 12'hffd; 
        10'b0010010001: data <= 12'hffe; 
        10'b0010010010: data <= 12'hffe; 
        10'b0010010011: data <= 12'hff9; 
        10'b0010010100: data <= 12'hffd; 
        10'b0010010101: data <= 12'h002; 
        10'b0010010110: data <= 12'hffa; 
        10'b0010010111: data <= 12'h007; 
        10'b0010011000: data <= 12'h00e; 
        10'b0010011001: data <= 12'h00c; 
        10'b0010011010: data <= 12'h00c; 
        10'b0010011011: data <= 12'h006; 
        10'b0010011100: data <= 12'h005; 
        10'b0010011101: data <= 12'h00b; 
        10'b0010011110: data <= 12'h001; 
        10'b0010011111: data <= 12'hfff; 
        10'b0010100000: data <= 12'h004; 
        10'b0010100001: data <= 12'h002; 
        10'b0010100010: data <= 12'hff9; 
        10'b0010100011: data <= 12'hffa; 
        10'b0010100100: data <= 12'hffc; 
        10'b0010100101: data <= 12'h003; 
        10'b0010100110: data <= 12'hfff; 
        10'b0010100111: data <= 12'h001; 
        10'b0010101000: data <= 12'hffd; 
        10'b0010101001: data <= 12'hffd; 
        10'b0010101010: data <= 12'hffc; 
        10'b0010101011: data <= 12'hffc; 
        10'b0010101100: data <= 12'hffc; 
        10'b0010101101: data <= 12'hffc; 
        10'b0010101110: data <= 12'hffa; 
        10'b0010101111: data <= 12'hffa; 
        10'b0010110000: data <= 12'h000; 
        10'b0010110001: data <= 12'h002; 
        10'b0010110010: data <= 12'h000; 
        10'b0010110011: data <= 12'h004; 
        10'b0010110100: data <= 12'h006; 
        10'b0010110101: data <= 12'h005; 
        10'b0010110110: data <= 12'h006; 
        10'b0010110111: data <= 12'h00c; 
        10'b0010111000: data <= 12'h006; 
        10'b0010111001: data <= 12'h007; 
        10'b0010111010: data <= 12'h001; 
        10'b0010111011: data <= 12'h008; 
        10'b0010111100: data <= 12'h003; 
        10'b0010111101: data <= 12'h004; 
        10'b0010111110: data <= 12'h005; 
        10'b0010111111: data <= 12'h004; 
        10'b0011000000: data <= 12'h004; 
        10'b0011000001: data <= 12'h002; 
        10'b0011000010: data <= 12'hfff; 
        10'b0011000011: data <= 12'h000; 
        10'b0011000100: data <= 12'h001; 
        10'b0011000101: data <= 12'hffd; 
        10'b0011000110: data <= 12'hffd; 
        10'b0011000111: data <= 12'hffe; 
        10'b0011001000: data <= 12'hffc; 
        10'b0011001001: data <= 12'hffe; 
        10'b0011001010: data <= 12'hffc; 
        10'b0011001011: data <= 12'h000; 
        10'b0011001100: data <= 12'h004; 
        10'b0011001101: data <= 12'h002; 
        10'b0011001110: data <= 12'h002; 
        10'b0011001111: data <= 12'hfff; 
        10'b0011010000: data <= 12'hffb; 
        10'b0011010001: data <= 12'hffc; 
        10'b0011010010: data <= 12'hffa; 
        10'b0011010011: data <= 12'h004; 
        10'b0011010100: data <= 12'h005; 
        10'b0011010101: data <= 12'h000; 
        10'b0011010110: data <= 12'h003; 
        10'b0011010111: data <= 12'hffd; 
        10'b0011011000: data <= 12'h005; 
        10'b0011011001: data <= 12'h007; 
        10'b0011011010: data <= 12'h001; 
        10'b0011011011: data <= 12'h00f; 
        10'b0011011100: data <= 12'h009; 
        10'b0011011101: data <= 12'h000; 
        10'b0011011110: data <= 12'h000; 
        10'b0011011111: data <= 12'hfff; 
        10'b0011100000: data <= 12'hfff; 
        10'b0011100001: data <= 12'h000; 
        10'b0011100010: data <= 12'hfff; 
        10'b0011100011: data <= 12'hffd; 
        10'b0011100100: data <= 12'hfff; 
        10'b0011100101: data <= 12'hfff; 
        10'b0011100110: data <= 12'h006; 
        10'b0011100111: data <= 12'h004; 
        10'b0011101000: data <= 12'h001; 
        10'b0011101001: data <= 12'h00b; 
        10'b0011101010: data <= 12'h001; 
        10'b0011101011: data <= 12'h000; 
        10'b0011101100: data <= 12'h007; 
        10'b0011101101: data <= 12'h009; 
        10'b0011101110: data <= 12'hff9; 
        10'b0011101111: data <= 12'hffa; 
        10'b0011110000: data <= 12'h005; 
        10'b0011110001: data <= 12'hffc; 
        10'b0011110010: data <= 12'h002; 
        10'b0011110011: data <= 12'h005; 
        10'b0011110100: data <= 12'h003; 
        10'b0011110101: data <= 12'h00a; 
        10'b0011110110: data <= 12'h007; 
        10'b0011110111: data <= 12'h00b; 
        10'b0011111000: data <= 12'h00a; 
        10'b0011111001: data <= 12'hfff; 
        10'b0011111010: data <= 12'hfff; 
        10'b0011111011: data <= 12'h001; 
        10'b0011111100: data <= 12'h000; 
        10'b0011111101: data <= 12'h000; 
        10'b0011111110: data <= 12'hffe; 
        10'b0011111111: data <= 12'hffe; 
        10'b0100000000: data <= 12'hfff; 
        10'b0100000001: data <= 12'h006; 
        10'b0100000010: data <= 12'h005; 
        10'b0100000011: data <= 12'h00a; 
        10'b0100000100: data <= 12'h00d; 
        10'b0100000101: data <= 12'h00b; 
        10'b0100000110: data <= 12'h007; 
        10'b0100000111: data <= 12'h00c; 
        10'b0100001000: data <= 12'h003; 
        10'b0100001001: data <= 12'h004; 
        10'b0100001010: data <= 12'hff2; 
        10'b0100001011: data <= 12'hfec; 
        10'b0100001100: data <= 12'hff9; 
        10'b0100001101: data <= 12'h001; 
        10'b0100001110: data <= 12'h002; 
        10'b0100001111: data <= 12'h004; 
        10'b0100010000: data <= 12'h005; 
        10'b0100010001: data <= 12'h004; 
        10'b0100010010: data <= 12'h00a; 
        10'b0100010011: data <= 12'h00b; 
        10'b0100010100: data <= 12'hffe; 
        10'b0100010101: data <= 12'hfff; 
        10'b0100010110: data <= 12'h002; 
        10'b0100010111: data <= 12'hffd; 
        10'b0100011000: data <= 12'hffd; 
        10'b0100011001: data <= 12'h000; 
        10'b0100011010: data <= 12'hffd; 
        10'b0100011011: data <= 12'h000; 
        10'b0100011100: data <= 12'h002; 
        10'b0100011101: data <= 12'h008; 
        10'b0100011110: data <= 12'h008; 
        10'b0100011111: data <= 12'h00e; 
        10'b0100100000: data <= 12'h00a; 
        10'b0100100001: data <= 12'h00c; 
        10'b0100100010: data <= 12'h012; 
        10'b0100100011: data <= 12'h009; 
        10'b0100100100: data <= 12'h009; 
        10'b0100100101: data <= 12'h007; 
        10'b0100100110: data <= 12'hffe; 
        10'b0100100111: data <= 12'hfed; 
        10'b0100101000: data <= 12'hff1; 
        10'b0100101001: data <= 12'hffb; 
        10'b0100101010: data <= 12'h005; 
        10'b0100101011: data <= 12'h005; 
        10'b0100101100: data <= 12'h005; 
        10'b0100101101: data <= 12'h00d; 
        10'b0100101110: data <= 12'h00e; 
        10'b0100101111: data <= 12'h00b; 
        10'b0100110000: data <= 12'h000; 
        10'b0100110001: data <= 12'hfff; 
        10'b0100110010: data <= 12'hfff; 
        10'b0100110011: data <= 12'hffe; 
        10'b0100110100: data <= 12'hffd; 
        10'b0100110101: data <= 12'h001; 
        10'b0100110110: data <= 12'h000; 
        10'b0100110111: data <= 12'hffc; 
        10'b0100111000: data <= 12'h004; 
        10'b0100111001: data <= 12'h009; 
        10'b0100111010: data <= 12'h010; 
        10'b0100111011: data <= 12'h015; 
        10'b0100111100: data <= 12'h011; 
        10'b0100111101: data <= 12'h015; 
        10'b0100111110: data <= 12'h00e; 
        10'b0100111111: data <= 12'h007; 
        10'b0101000000: data <= 12'h009; 
        10'b0101000001: data <= 12'h015; 
        10'b0101000010: data <= 12'h019; 
        10'b0101000011: data <= 12'hffd; 
        10'b0101000100: data <= 12'hff1; 
        10'b0101000101: data <= 12'hffb; 
        10'b0101000110: data <= 12'hffb; 
        10'b0101000111: data <= 12'h002; 
        10'b0101001000: data <= 12'h00b; 
        10'b0101001001: data <= 12'h00e; 
        10'b0101001010: data <= 12'h012; 
        10'b0101001011: data <= 12'h011; 
        10'b0101001100: data <= 12'h00c; 
        10'b0101001101: data <= 12'h002; 
        10'b0101001110: data <= 12'h001; 
        10'b0101001111: data <= 12'hfff; 
        10'b0101010000: data <= 12'hffe; 
        10'b0101010001: data <= 12'hfff; 
        10'b0101010010: data <= 12'hffe; 
        10'b0101010011: data <= 12'hfff; 
        10'b0101010100: data <= 12'hfff; 
        10'b0101010101: data <= 12'h00a; 
        10'b0101010110: data <= 12'h008; 
        10'b0101010111: data <= 12'h00d; 
        10'b0101011000: data <= 12'h00c; 
        10'b0101011001: data <= 12'h00f; 
        10'b0101011010: data <= 12'h003; 
        10'b0101011011: data <= 12'h004; 
        10'b0101011100: data <= 12'h002; 
        10'b0101011101: data <= 12'h019; 
        10'b0101011110: data <= 12'h019; 
        10'b0101011111: data <= 12'h006; 
        10'b0101100000: data <= 12'h001; 
        10'b0101100001: data <= 12'hffe; 
        10'b0101100010: data <= 12'hffe; 
        10'b0101100011: data <= 12'h006; 
        10'b0101100100: data <= 12'h00b; 
        10'b0101100101: data <= 12'h013; 
        10'b0101100110: data <= 12'h016; 
        10'b0101100111: data <= 12'h012; 
        10'b0101101000: data <= 12'h00b; 
        10'b0101101001: data <= 12'h005; 
        10'b0101101010: data <= 12'h002; 
        10'b0101101011: data <= 12'hffd; 
        10'b0101101100: data <= 12'hffc; 
        10'b0101101101: data <= 12'hfff; 
        10'b0101101110: data <= 12'h001; 
        10'b0101101111: data <= 12'hffd; 
        10'b0101110000: data <= 12'hffe; 
        10'b0101110001: data <= 12'h000; 
        10'b0101110010: data <= 12'hffe; 
        10'b0101110011: data <= 12'hffe; 
        10'b0101110100: data <= 12'h001; 
        10'b0101110101: data <= 12'hffe; 
        10'b0101110110: data <= 12'hffa; 
        10'b0101110111: data <= 12'h002; 
        10'b0101111000: data <= 12'h009; 
        10'b0101111001: data <= 12'h018; 
        10'b0101111010: data <= 12'h007; 
        10'b0101111011: data <= 12'h011; 
        10'b0101111100: data <= 12'h007; 
        10'b0101111101: data <= 12'hffc; 
        10'b0101111110: data <= 12'h000; 
        10'b0101111111: data <= 12'h001; 
        10'b0110000000: data <= 12'h008; 
        10'b0110000001: data <= 12'h007; 
        10'b0110000010: data <= 12'h004; 
        10'b0110000011: data <= 12'h006; 
        10'b0110000100: data <= 12'h003; 
        10'b0110000101: data <= 12'h001; 
        10'b0110000110: data <= 12'h001; 
        10'b0110000111: data <= 12'hfff; 
        10'b0110001000: data <= 12'hffe; 
        10'b0110001001: data <= 12'hffc; 
        10'b0110001010: data <= 12'h000; 
        10'b0110001011: data <= 12'hfff; 
        10'b0110001100: data <= 12'hffd; 
        10'b0110001101: data <= 12'hff9; 
        10'b0110001110: data <= 12'hff4; 
        10'b0110001111: data <= 12'hff0; 
        10'b0110010000: data <= 12'hfed; 
        10'b0110010001: data <= 12'hff1; 
        10'b0110010010: data <= 12'hffe; 
        10'b0110010011: data <= 12'h009; 
        10'b0110010100: data <= 12'h009; 
        10'b0110010101: data <= 12'h013; 
        10'b0110010110: data <= 12'h00f; 
        10'b0110010111: data <= 12'h00a; 
        10'b0110011000: data <= 12'hfff; 
        10'b0110011001: data <= 12'h001; 
        10'b0110011010: data <= 12'hffd; 
        10'b0110011011: data <= 12'hffa; 
        10'b0110011100: data <= 12'hff6; 
        10'b0110011101: data <= 12'hff7; 
        10'b0110011110: data <= 12'hff8; 
        10'b0110011111: data <= 12'hff7; 
        10'b0110100000: data <= 12'hffc; 
        10'b0110100001: data <= 12'hfff; 
        10'b0110100010: data <= 12'hffc; 
        10'b0110100011: data <= 12'h000; 
        10'b0110100100: data <= 12'h000; 
        10'b0110100101: data <= 12'hffe; 
        10'b0110100110: data <= 12'hffd; 
        10'b0110100111: data <= 12'hfff; 
        10'b0110101000: data <= 12'hffd; 
        10'b0110101001: data <= 12'hff9; 
        10'b0110101010: data <= 12'hff1; 
        10'b0110101011: data <= 12'hfed; 
        10'b0110101100: data <= 12'hfef; 
        10'b0110101101: data <= 12'hffc; 
        10'b0110101110: data <= 12'h001; 
        10'b0110101111: data <= 12'h000; 
        10'b0110110000: data <= 12'h00d; 
        10'b0110110001: data <= 12'h010; 
        10'b0110110010: data <= 12'h00e; 
        10'b0110110011: data <= 12'h008; 
        10'b0110110100: data <= 12'hffc; 
        10'b0110110101: data <= 12'hffd; 
        10'b0110110110: data <= 12'hffe; 
        10'b0110110111: data <= 12'hff2; 
        10'b0110111000: data <= 12'hfef; 
        10'b0110111001: data <= 12'hff3; 
        10'b0110111010: data <= 12'hff8; 
        10'b0110111011: data <= 12'hff8; 
        10'b0110111100: data <= 12'hffa; 
        10'b0110111101: data <= 12'hfff; 
        10'b0110111110: data <= 12'hffc; 
        10'b0110111111: data <= 12'h000; 
        10'b0111000000: data <= 12'hffe; 
        10'b0111000001: data <= 12'hffd; 
        10'b0111000010: data <= 12'hffe; 
        10'b0111000011: data <= 12'hfff; 
        10'b0111000100: data <= 12'hffa; 
        10'b0111000101: data <= 12'hff6; 
        10'b0111000110: data <= 12'hff0; 
        10'b0111000111: data <= 12'hff7; 
        10'b0111001000: data <= 12'h006; 
        10'b0111001001: data <= 12'h007; 
        10'b0111001010: data <= 12'h003; 
        10'b0111001011: data <= 12'h006; 
        10'b0111001100: data <= 12'h00d; 
        10'b0111001101: data <= 12'h00b; 
        10'b0111001110: data <= 12'h004; 
        10'b0111001111: data <= 12'h007; 
        10'b0111010000: data <= 12'h002; 
        10'b0111010001: data <= 12'hffb; 
        10'b0111010010: data <= 12'hff5; 
        10'b0111010011: data <= 12'hff0; 
        10'b0111010100: data <= 12'hff0; 
        10'b0111010101: data <= 12'hff0; 
        10'b0111010110: data <= 12'hff3; 
        10'b0111010111: data <= 12'hffc; 
        10'b0111011000: data <= 12'hffa; 
        10'b0111011001: data <= 12'hffe; 
        10'b0111011010: data <= 12'hffe; 
        10'b0111011011: data <= 12'hffc; 
        10'b0111011100: data <= 12'h001; 
        10'b0111011101: data <= 12'h001; 
        10'b0111011110: data <= 12'hffd; 
        10'b0111011111: data <= 12'hffd; 
        10'b0111100000: data <= 12'hffc; 
        10'b0111100001: data <= 12'hff6; 
        10'b0111100010: data <= 12'hff2; 
        10'b0111100011: data <= 12'h002; 
        10'b0111100100: data <= 12'h00d; 
        10'b0111100101: data <= 12'h010; 
        10'b0111100110: data <= 12'h005; 
        10'b0111100111: data <= 12'h00c; 
        10'b0111101000: data <= 12'h014; 
        10'b0111101001: data <= 12'h00c; 
        10'b0111101010: data <= 12'h001; 
        10'b0111101011: data <= 12'hffd; 
        10'b0111101100: data <= 12'h001; 
        10'b0111101101: data <= 12'hffa; 
        10'b0111101110: data <= 12'hff0; 
        10'b0111101111: data <= 12'hff8; 
        10'b0111110000: data <= 12'hff8; 
        10'b0111110001: data <= 12'hff5; 
        10'b0111110010: data <= 12'hff8; 
        10'b0111110011: data <= 12'hffb; 
        10'b0111110100: data <= 12'hffd; 
        10'b0111110101: data <= 12'hffc; 
        10'b0111110110: data <= 12'hfff; 
        10'b0111110111: data <= 12'hffe; 
        10'b0111111000: data <= 12'hffe; 
        10'b0111111001: data <= 12'h000; 
        10'b0111111010: data <= 12'hffc; 
        10'b0111111011: data <= 12'hffb; 
        10'b0111111100: data <= 12'hffa; 
        10'b0111111101: data <= 12'hffa; 
        10'b0111111110: data <= 12'hffc; 
        10'b0111111111: data <= 12'h004; 
        10'b1000000000: data <= 12'h00b; 
        10'b1000000001: data <= 12'h013; 
        10'b1000000010: data <= 12'h00d; 
        10'b1000000011: data <= 12'h012; 
        10'b1000000100: data <= 12'h00c; 
        10'b1000000101: data <= 12'h007; 
        10'b1000000110: data <= 12'hff8; 
        10'b1000000111: data <= 12'hffe; 
        10'b1000001000: data <= 12'hffb; 
        10'b1000001001: data <= 12'hff3; 
        10'b1000001010: data <= 12'hffd; 
        10'b1000001011: data <= 12'hffe; 
        10'b1000001100: data <= 12'h001; 
        10'b1000001101: data <= 12'hff9; 
        10'b1000001110: data <= 12'hfff; 
        10'b1000001111: data <= 12'hffa; 
        10'b1000010000: data <= 12'hff8; 
        10'b1000010001: data <= 12'hffc; 
        10'b1000010010: data <= 12'hfff; 
        10'b1000010011: data <= 12'h001; 
        10'b1000010100: data <= 12'hffe; 
        10'b1000010101: data <= 12'hfff; 
        10'b1000010110: data <= 12'hfff; 
        10'b1000010111: data <= 12'hffb; 
        10'b1000011000: data <= 12'hff9; 
        10'b1000011001: data <= 12'hffd; 
        10'b1000011010: data <= 12'h002; 
        10'b1000011011: data <= 12'h005; 
        10'b1000011100: data <= 12'h005; 
        10'b1000011101: data <= 12'h00d; 
        10'b1000011110: data <= 12'h007; 
        10'b1000011111: data <= 12'hfff; 
        10'b1000100000: data <= 12'h003; 
        10'b1000100001: data <= 12'hff7; 
        10'b1000100010: data <= 12'hff6; 
        10'b1000100011: data <= 12'hffc; 
        10'b1000100100: data <= 12'hffd; 
        10'b1000100101: data <= 12'hffc; 
        10'b1000100110: data <= 12'h003; 
        10'b1000100111: data <= 12'h001; 
        10'b1000101000: data <= 12'h004; 
        10'b1000101001: data <= 12'h000; 
        10'b1000101010: data <= 12'h003; 
        10'b1000101011: data <= 12'hffe; 
        10'b1000101100: data <= 12'hffa; 
        10'b1000101101: data <= 12'hffc; 
        10'b1000101110: data <= 12'hffd; 
        10'b1000101111: data <= 12'h000; 
        10'b1000110000: data <= 12'hffd; 
        10'b1000110001: data <= 12'hfff; 
        10'b1000110010: data <= 12'hffd; 
        10'b1000110011: data <= 12'hffc; 
        10'b1000110100: data <= 12'hff8; 
        10'b1000110101: data <= 12'hfff; 
        10'b1000110110: data <= 12'h001; 
        10'b1000110111: data <= 12'h00b; 
        10'b1000111000: data <= 12'h003; 
        10'b1000111001: data <= 12'hfff; 
        10'b1000111010: data <= 12'h000; 
        10'b1000111011: data <= 12'hff6; 
        10'b1000111100: data <= 12'h001; 
        10'b1000111101: data <= 12'h000; 
        10'b1000111110: data <= 12'hff7; 
        10'b1000111111: data <= 12'hffe; 
        10'b1001000000: data <= 12'hff5; 
        10'b1001000001: data <= 12'hffd; 
        10'b1001000010: data <= 12'h002; 
        10'b1001000011: data <= 12'h001; 
        10'b1001000100: data <= 12'h003; 
        10'b1001000101: data <= 12'h006; 
        10'b1001000110: data <= 12'h006; 
        10'b1001000111: data <= 12'hfff; 
        10'b1001001000: data <= 12'hffc; 
        10'b1001001001: data <= 12'hffb; 
        10'b1001001010: data <= 12'hfff; 
        10'b1001001011: data <= 12'hffd; 
        10'b1001001100: data <= 12'h000; 
        10'b1001001101: data <= 12'hffe; 
        10'b1001001110: data <= 12'h001; 
        10'b1001001111: data <= 12'hffa; 
        10'b1001010000: data <= 12'hff7; 
        10'b1001010001: data <= 12'hfff; 
        10'b1001010010: data <= 12'h005; 
        10'b1001010011: data <= 12'h00a; 
        10'b1001010100: data <= 12'h002; 
        10'b1001010101: data <= 12'h004; 
        10'b1001010110: data <= 12'hfff; 
        10'b1001010111: data <= 12'hff9; 
        10'b1001011000: data <= 12'hffc; 
        10'b1001011001: data <= 12'h002; 
        10'b1001011010: data <= 12'h000; 
        10'b1001011011: data <= 12'hfff; 
        10'b1001011100: data <= 12'hff8; 
        10'b1001011101: data <= 12'hffd; 
        10'b1001011110: data <= 12'hffe; 
        10'b1001011111: data <= 12'h000; 
        10'b1001100000: data <= 12'h000; 
        10'b1001100001: data <= 12'h002; 
        10'b1001100010: data <= 12'h002; 
        10'b1001100011: data <= 12'hffe; 
        10'b1001100100: data <= 12'hffd; 
        10'b1001100101: data <= 12'h000; 
        10'b1001100110: data <= 12'hfff; 
        10'b1001100111: data <= 12'hffe; 
        10'b1001101000: data <= 12'hfff; 
        10'b1001101001: data <= 12'hffc; 
        10'b1001101010: data <= 12'hffe; 
        10'b1001101011: data <= 12'hffc; 
        10'b1001101100: data <= 12'hff9; 
        10'b1001101101: data <= 12'hff5; 
        10'b1001101110: data <= 12'h001; 
        10'b1001101111: data <= 12'h003; 
        10'b1001110000: data <= 12'hfff; 
        10'b1001110001: data <= 12'hffc; 
        10'b1001110010: data <= 12'h002; 
        10'b1001110011: data <= 12'h001; 
        10'b1001110100: data <= 12'h00d; 
        10'b1001110101: data <= 12'h00e; 
        10'b1001110110: data <= 12'h00a; 
        10'b1001110111: data <= 12'h008; 
        10'b1001111000: data <= 12'hfff; 
        10'b1001111001: data <= 12'hfff; 
        10'b1001111010: data <= 12'h003; 
        10'b1001111011: data <= 12'hffc; 
        10'b1001111100: data <= 12'hffc; 
        10'b1001111101: data <= 12'h002; 
        10'b1001111110: data <= 12'hfff; 
        10'b1001111111: data <= 12'hffd; 
        10'b1010000000: data <= 12'hfff; 
        10'b1010000001: data <= 12'hfff; 
        10'b1010000010: data <= 12'hfff; 
        10'b1010000011: data <= 12'hffd; 
        10'b1010000100: data <= 12'hffd; 
        10'b1010000101: data <= 12'h000; 
        10'b1010000110: data <= 12'hfff; 
        10'b1010000111: data <= 12'hffc; 
        10'b1010001000: data <= 12'hff8; 
        10'b1010001001: data <= 12'hfed; 
        10'b1010001010: data <= 12'hff1; 
        10'b1010001011: data <= 12'hff9; 
        10'b1010001100: data <= 12'h003; 
        10'b1010001101: data <= 12'h002; 
        10'b1010001110: data <= 12'h005; 
        10'b1010001111: data <= 12'h007; 
        10'b1010010000: data <= 12'h010; 
        10'b1010010001: data <= 12'h017; 
        10'b1010010010: data <= 12'h013; 
        10'b1010010011: data <= 12'h00f; 
        10'b1010010100: data <= 12'h00c; 
        10'b1010010101: data <= 12'h009; 
        10'b1010010110: data <= 12'h007; 
        10'b1010010111: data <= 12'h009; 
        10'b1010011000: data <= 12'h007; 
        10'b1010011001: data <= 12'h002; 
        10'b1010011010: data <= 12'hfff; 
        10'b1010011011: data <= 12'hffe; 
        10'b1010011100: data <= 12'hffc; 
        10'b1010011101: data <= 12'h000; 
        10'b1010011110: data <= 12'hffc; 
        10'b1010011111: data <= 12'hfff; 
        10'b1010100000: data <= 12'h000; 
        10'b1010100001: data <= 12'hfff; 
        10'b1010100010: data <= 12'h001; 
        10'b1010100011: data <= 12'hffd; 
        10'b1010100100: data <= 12'hffd; 
        10'b1010100101: data <= 12'hff4; 
        10'b1010100110: data <= 12'hfef; 
        10'b1010100111: data <= 12'hff2; 
        10'b1010101000: data <= 12'hfff; 
        10'b1010101001: data <= 12'h003; 
        10'b1010101010: data <= 12'hfff; 
        10'b1010101011: data <= 12'h006; 
        10'b1010101100: data <= 12'h004; 
        10'b1010101101: data <= 12'h003; 
        10'b1010101110: data <= 12'h007; 
        10'b1010101111: data <= 12'h010; 
        10'b1010110000: data <= 12'h011; 
        10'b1010110001: data <= 12'h00b; 
        10'b1010110010: data <= 12'h010; 
        10'b1010110011: data <= 12'h00f; 
        10'b1010110100: data <= 12'h005; 
        10'b1010110101: data <= 12'h000; 
        10'b1010110110: data <= 12'hffd; 
        10'b1010110111: data <= 12'h000; 
        10'b1010111000: data <= 12'hfff; 
        10'b1010111001: data <= 12'hffe; 
        10'b1010111010: data <= 12'h001; 
        10'b1010111011: data <= 12'hfff; 
        10'b1010111100: data <= 12'h001; 
        10'b1010111101: data <= 12'hfff; 
        10'b1010111110: data <= 12'h000; 
        10'b1010111111: data <= 12'hffd; 
        10'b1011000000: data <= 12'hffe; 
        10'b1011000001: data <= 12'hffb; 
        10'b1011000010: data <= 12'hffa; 
        10'b1011000011: data <= 12'hff8; 
        10'b1011000100: data <= 12'hff7; 
        10'b1011000101: data <= 12'hff7; 
        10'b1011000110: data <= 12'hffd; 
        10'b1011000111: data <= 12'hffa; 
        10'b1011001000: data <= 12'hffc; 
        10'b1011001001: data <= 12'hffc; 
        10'b1011001010: data <= 12'h000; 
        10'b1011001011: data <= 12'h006; 
        10'b1011001100: data <= 12'h004; 
        10'b1011001101: data <= 12'h005; 
        10'b1011001110: data <= 12'h006; 
        10'b1011001111: data <= 12'h001; 
        10'b1011010000: data <= 12'hfff; 
        10'b1011010001: data <= 12'h000; 
        10'b1011010010: data <= 12'hffc; 
        10'b1011010011: data <= 12'hffc; 
        10'b1011010100: data <= 12'h000; 
        10'b1011010101: data <= 12'hfff; 
        10'b1011010110: data <= 12'hffe; 
        10'b1011010111: data <= 12'hfff; 
        10'b1011011000: data <= 12'hfff; 
        10'b1011011001: data <= 12'h000; 
        10'b1011011010: data <= 12'hffe; 
        10'b1011011011: data <= 12'hffd; 
        10'b1011011100: data <= 12'hffc; 
        10'b1011011101: data <= 12'hffd; 
        10'b1011011110: data <= 12'hffb; 
        10'b1011011111: data <= 12'hfff; 
        10'b1011100000: data <= 12'hffc; 
        10'b1011100001: data <= 12'hffc; 
        10'b1011100010: data <= 12'hffb; 
        10'b1011100011: data <= 12'hffd; 
        10'b1011100100: data <= 12'hffd; 
        10'b1011100101: data <= 12'hffe; 
        10'b1011100110: data <= 12'hffc; 
        10'b1011100111: data <= 12'hffd; 
        10'b1011101000: data <= 12'hffd; 
        10'b1011101001: data <= 12'hffc; 
        10'b1011101010: data <= 12'hffb; 
        10'b1011101011: data <= 12'hffd; 
        10'b1011101100: data <= 12'hffe; 
        10'b1011101101: data <= 12'hfff; 
        10'b1011101110: data <= 12'hffe; 
        10'b1011101111: data <= 12'h001; 
        10'b1011110000: data <= 12'h001; 
        10'b1011110001: data <= 12'hffd; 
        10'b1011110010: data <= 12'hfff; 
        10'b1011110011: data <= 12'hfff; 
        10'b1011110100: data <= 12'hfff; 
        10'b1011110101: data <= 12'hffd; 
        10'b1011110110: data <= 12'hffe; 
        10'b1011110111: data <= 12'hfff; 
        10'b1011111000: data <= 12'hfff; 
        10'b1011111001: data <= 12'hffc; 
        10'b1011111010: data <= 12'h000; 
        10'b1011111011: data <= 12'hffe; 
        10'b1011111100: data <= 12'h001; 
        10'b1011111101: data <= 12'hffe; 
        10'b1011111110: data <= 12'hffd; 
        10'b1011111111: data <= 12'h000; 
        10'b1100000000: data <= 12'hffd; 
        10'b1100000001: data <= 12'hffd; 
        10'b1100000010: data <= 12'hffe; 
        10'b1100000011: data <= 12'hfff; 
        10'b1100000100: data <= 12'hfff; 
        10'b1100000101: data <= 12'h000; 
        10'b1100000110: data <= 12'h000; 
        10'b1100000111: data <= 12'h001; 
        10'b1100001000: data <= 12'hfff; 
        10'b1100001001: data <= 12'hfff; 
        10'b1100001010: data <= 12'hfff; 
        10'b1100001011: data <= 12'hffd; 
        10'b1100001100: data <= 12'hfff; 
        10'b1100001101: data <= 12'h001; 
        10'b1100001110: data <= 12'hffd; 
        10'b1100001111: data <= 12'hfff; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 7) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 13'h1ffc; 
        10'b0000000001: data <= 13'h1ffd; 
        10'b0000000010: data <= 13'h1ffd; 
        10'b0000000011: data <= 13'h1ffe; 
        10'b0000000100: data <= 13'h1ffe; 
        10'b0000000101: data <= 13'h0001; 
        10'b0000000110: data <= 13'h1ff9; 
        10'b0000000111: data <= 13'h1ffe; 
        10'b0000001000: data <= 13'h1ffb; 
        10'b0000001001: data <= 13'h1ffc; 
        10'b0000001010: data <= 13'h1ffa; 
        10'b0000001011: data <= 13'h0001; 
        10'b0000001100: data <= 13'h1ffe; 
        10'b0000001101: data <= 13'h0000; 
        10'b0000001110: data <= 13'h1ffa; 
        10'b0000001111: data <= 13'h0000; 
        10'b0000010000: data <= 13'h1ffe; 
        10'b0000010001: data <= 13'h1ff9; 
        10'b0000010010: data <= 13'h0001; 
        10'b0000010011: data <= 13'h1ffd; 
        10'b0000010100: data <= 13'h1ffd; 
        10'b0000010101: data <= 13'h1ffc; 
        10'b0000010110: data <= 13'h1ffd; 
        10'b0000010111: data <= 13'h0001; 
        10'b0000011000: data <= 13'h0000; 
        10'b0000011001: data <= 13'h1ffc; 
        10'b0000011010: data <= 13'h1ffb; 
        10'b0000011011: data <= 13'h1ffd; 
        10'b0000011100: data <= 13'h1ffd; 
        10'b0000011101: data <= 13'h1ff9; 
        10'b0000011110: data <= 13'h0001; 
        10'b0000011111: data <= 13'h0000; 
        10'b0000100000: data <= 13'h1ff9; 
        10'b0000100001: data <= 13'h1ffa; 
        10'b0000100010: data <= 13'h1ff9; 
        10'b0000100011: data <= 13'h1ffa; 
        10'b0000100100: data <= 13'h0001; 
        10'b0000100101: data <= 13'h1ffd; 
        10'b0000100110: data <= 13'h1ffd; 
        10'b0000100111: data <= 13'h1ff9; 
        10'b0000101000: data <= 13'h0001; 
        10'b0000101001: data <= 13'h1fff; 
        10'b0000101010: data <= 13'h1ffb; 
        10'b0000101011: data <= 13'h1ffc; 
        10'b0000101100: data <= 13'h1fff; 
        10'b0000101101: data <= 13'h1ffe; 
        10'b0000101110: data <= 13'h1ffa; 
        10'b0000101111: data <= 13'h1ffe; 
        10'b0000110000: data <= 13'h0001; 
        10'b0000110001: data <= 13'h1ff9; 
        10'b0000110010: data <= 13'h1fff; 
        10'b0000110011: data <= 13'h1ffa; 
        10'b0000110100: data <= 13'h1fff; 
        10'b0000110101: data <= 13'h0002; 
        10'b0000110110: data <= 13'h1ffb; 
        10'b0000110111: data <= 13'h1ffa; 
        10'b0000111000: data <= 13'h1ffa; 
        10'b0000111001: data <= 13'h0000; 
        10'b0000111010: data <= 13'h1ffe; 
        10'b0000111011: data <= 13'h1ffd; 
        10'b0000111100: data <= 13'h1ffa; 
        10'b0000111101: data <= 13'h1ff9; 
        10'b0000111110: data <= 13'h1ffe; 
        10'b0000111111: data <= 13'h1ff9; 
        10'b0001000000: data <= 13'h0001; 
        10'b0001000001: data <= 13'h1ff9; 
        10'b0001000010: data <= 13'h1ff9; 
        10'b0001000011: data <= 13'h1fff; 
        10'b0001000100: data <= 13'h1ffe; 
        10'b0001000101: data <= 13'h1ff8; 
        10'b0001000110: data <= 13'h1ffe; 
        10'b0001000111: data <= 13'h1ffe; 
        10'b0001001000: data <= 13'h1ff8; 
        10'b0001001001: data <= 13'h1ffb; 
        10'b0001001010: data <= 13'h1ffb; 
        10'b0001001011: data <= 13'h1fff; 
        10'b0001001100: data <= 13'h0000; 
        10'b0001001101: data <= 13'h0000; 
        10'b0001001110: data <= 13'h1ffe; 
        10'b0001001111: data <= 13'h1ffd; 
        10'b0001010000: data <= 13'h0001; 
        10'b0001010001: data <= 13'h1ffb; 
        10'b0001010010: data <= 13'h1fff; 
        10'b0001010011: data <= 13'h0001; 
        10'b0001010100: data <= 13'h1ffb; 
        10'b0001010101: data <= 13'h1ffd; 
        10'b0001010110: data <= 13'h1ffd; 
        10'b0001010111: data <= 13'h1ffa; 
        10'b0001011000: data <= 13'h0001; 
        10'b0001011001: data <= 13'h1ffa; 
        10'b0001011010: data <= 13'h1ff9; 
        10'b0001011011: data <= 13'h1ffc; 
        10'b0001011100: data <= 13'h1ff9; 
        10'b0001011101: data <= 13'h1ffd; 
        10'b0001011110: data <= 13'h1ffb; 
        10'b0001011111: data <= 13'h1ff6; 
        10'b0001100000: data <= 13'h1ff5; 
        10'b0001100001: data <= 13'h1ff2; 
        10'b0001100010: data <= 13'h1ff5; 
        10'b0001100011: data <= 13'h1ff9; 
        10'b0001100100: data <= 13'h1ff5; 
        10'b0001100101: data <= 13'h1ff7; 
        10'b0001100110: data <= 13'h1ffa; 
        10'b0001100111: data <= 13'h1ffc; 
        10'b0001101000: data <= 13'h1ff7; 
        10'b0001101001: data <= 13'h0001; 
        10'b0001101010: data <= 13'h1ffc; 
        10'b0001101011: data <= 13'h0000; 
        10'b0001101100: data <= 13'h1ffb; 
        10'b0001101101: data <= 13'h1ffe; 
        10'b0001101110: data <= 13'h1ffe; 
        10'b0001101111: data <= 13'h1ff9; 
        10'b0001110000: data <= 13'h1ffd; 
        10'b0001110001: data <= 13'h1fff; 
        10'b0001110010: data <= 13'h1ffc; 
        10'b0001110011: data <= 13'h1ff9; 
        10'b0001110100: data <= 13'h0000; 
        10'b0001110101: data <= 13'h1fff; 
        10'b0001110110: data <= 13'h1ffd; 
        10'b0001110111: data <= 13'h1ffa; 
        10'b0001111000: data <= 13'h1ffa; 
        10'b0001111001: data <= 13'h1ffc; 
        10'b0001111010: data <= 13'h1ffd; 
        10'b0001111011: data <= 13'h1ffe; 
        10'b0001111100: data <= 13'h000a; 
        10'b0001111101: data <= 13'h0006; 
        10'b0001111110: data <= 13'h0015; 
        10'b0001111111: data <= 13'h0010; 
        10'b0010000000: data <= 13'h0007; 
        10'b0010000001: data <= 13'h0004; 
        10'b0010000010: data <= 13'h0006; 
        10'b0010000011: data <= 13'h1ffb; 
        10'b0010000100: data <= 13'h1ff9; 
        10'b0010000101: data <= 13'h1ffd; 
        10'b0010000110: data <= 13'h1ff6; 
        10'b0010000111: data <= 13'h1ff9; 
        10'b0010001000: data <= 13'h0000; 
        10'b0010001001: data <= 13'h0000; 
        10'b0010001010: data <= 13'h1ffc; 
        10'b0010001011: data <= 13'h1ffd; 
        10'b0010001100: data <= 13'h1ffd; 
        10'b0010001101: data <= 13'h1fff; 
        10'b0010001110: data <= 13'h1fff; 
        10'b0010001111: data <= 13'h0000; 
        10'b0010010000: data <= 13'h1ffa; 
        10'b0010010001: data <= 13'h1ffd; 
        10'b0010010010: data <= 13'h1ffb; 
        10'b0010010011: data <= 13'h1ff3; 
        10'b0010010100: data <= 13'h1ffb; 
        10'b0010010101: data <= 13'h0005; 
        10'b0010010110: data <= 13'h1ff5; 
        10'b0010010111: data <= 13'h000f; 
        10'b0010011000: data <= 13'h001c; 
        10'b0010011001: data <= 13'h0017; 
        10'b0010011010: data <= 13'h0018; 
        10'b0010011011: data <= 13'h000c; 
        10'b0010011100: data <= 13'h0009; 
        10'b0010011101: data <= 13'h0016; 
        10'b0010011110: data <= 13'h0001; 
        10'b0010011111: data <= 13'h1fff; 
        10'b0010100000: data <= 13'h0008; 
        10'b0010100001: data <= 13'h0004; 
        10'b0010100010: data <= 13'h1ff2; 
        10'b0010100011: data <= 13'h1ff5; 
        10'b0010100100: data <= 13'h1ff8; 
        10'b0010100101: data <= 13'h0006; 
        10'b0010100110: data <= 13'h1ffe; 
        10'b0010100111: data <= 13'h0001; 
        10'b0010101000: data <= 13'h1ffb; 
        10'b0010101001: data <= 13'h1ffa; 
        10'b0010101010: data <= 13'h1ff9; 
        10'b0010101011: data <= 13'h1ff9; 
        10'b0010101100: data <= 13'h1ff8; 
        10'b0010101101: data <= 13'h1ff8; 
        10'b0010101110: data <= 13'h1ff3; 
        10'b0010101111: data <= 13'h1ff3; 
        10'b0010110000: data <= 13'h0001; 
        10'b0010110001: data <= 13'h0004; 
        10'b0010110010: data <= 13'h1fff; 
        10'b0010110011: data <= 13'h0007; 
        10'b0010110100: data <= 13'h000b; 
        10'b0010110101: data <= 13'h0009; 
        10'b0010110110: data <= 13'h000d; 
        10'b0010110111: data <= 13'h0018; 
        10'b0010111000: data <= 13'h000c; 
        10'b0010111001: data <= 13'h000e; 
        10'b0010111010: data <= 13'h0003; 
        10'b0010111011: data <= 13'h0010; 
        10'b0010111100: data <= 13'h0006; 
        10'b0010111101: data <= 13'h0007; 
        10'b0010111110: data <= 13'h0009; 
        10'b0010111111: data <= 13'h0008; 
        10'b0011000000: data <= 13'h0007; 
        10'b0011000001: data <= 13'h0003; 
        10'b0011000010: data <= 13'h1ffd; 
        10'b0011000011: data <= 13'h1fff; 
        10'b0011000100: data <= 13'h0001; 
        10'b0011000101: data <= 13'h1ffb; 
        10'b0011000110: data <= 13'h1ffa; 
        10'b0011000111: data <= 13'h1ffb; 
        10'b0011001000: data <= 13'h1ff8; 
        10'b0011001001: data <= 13'h1ffd; 
        10'b0011001010: data <= 13'h1ff7; 
        10'b0011001011: data <= 13'h1fff; 
        10'b0011001100: data <= 13'h0009; 
        10'b0011001101: data <= 13'h0004; 
        10'b0011001110: data <= 13'h0004; 
        10'b0011001111: data <= 13'h1ffd; 
        10'b0011010000: data <= 13'h1ff5; 
        10'b0011010001: data <= 13'h1ff8; 
        10'b0011010010: data <= 13'h1ff4; 
        10'b0011010011: data <= 13'h0007; 
        10'b0011010100: data <= 13'h0009; 
        10'b0011010101: data <= 13'h1fff; 
        10'b0011010110: data <= 13'h0006; 
        10'b0011010111: data <= 13'h1ff9; 
        10'b0011011000: data <= 13'h0009; 
        10'b0011011001: data <= 13'h000e; 
        10'b0011011010: data <= 13'h0003; 
        10'b0011011011: data <= 13'h001e; 
        10'b0011011100: data <= 13'h0012; 
        10'b0011011101: data <= 13'h1fff; 
        10'b0011011110: data <= 13'h0000; 
        10'b0011011111: data <= 13'h1fff; 
        10'b0011100000: data <= 13'h1fff; 
        10'b0011100001: data <= 13'h0000; 
        10'b0011100010: data <= 13'h1fff; 
        10'b0011100011: data <= 13'h1ffa; 
        10'b0011100100: data <= 13'h1ffe; 
        10'b0011100101: data <= 13'h1ffd; 
        10'b0011100110: data <= 13'h000c; 
        10'b0011100111: data <= 13'h0008; 
        10'b0011101000: data <= 13'h0003; 
        10'b0011101001: data <= 13'h0016; 
        10'b0011101010: data <= 13'h0001; 
        10'b0011101011: data <= 13'h0001; 
        10'b0011101100: data <= 13'h000e; 
        10'b0011101101: data <= 13'h0013; 
        10'b0011101110: data <= 13'h1ff1; 
        10'b0011101111: data <= 13'h1ff3; 
        10'b0011110000: data <= 13'h000a; 
        10'b0011110001: data <= 13'h1ff9; 
        10'b0011110010: data <= 13'h0003; 
        10'b0011110011: data <= 13'h000a; 
        10'b0011110100: data <= 13'h0006; 
        10'b0011110101: data <= 13'h0014; 
        10'b0011110110: data <= 13'h000d; 
        10'b0011110111: data <= 13'h0017; 
        10'b0011111000: data <= 13'h0015; 
        10'b0011111001: data <= 13'h1ffe; 
        10'b0011111010: data <= 13'h1ffe; 
        10'b0011111011: data <= 13'h0002; 
        10'b0011111100: data <= 13'h0000; 
        10'b0011111101: data <= 13'h0000; 
        10'b0011111110: data <= 13'h1ffd; 
        10'b0011111111: data <= 13'h1ffc; 
        10'b0100000000: data <= 13'h1ffe; 
        10'b0100000001: data <= 13'h000d; 
        10'b0100000010: data <= 13'h0009; 
        10'b0100000011: data <= 13'h0013; 
        10'b0100000100: data <= 13'h001a; 
        10'b0100000101: data <= 13'h0016; 
        10'b0100000110: data <= 13'h000e; 
        10'b0100000111: data <= 13'h0018; 
        10'b0100001000: data <= 13'h0007; 
        10'b0100001001: data <= 13'h0007; 
        10'b0100001010: data <= 13'h1fe4; 
        10'b0100001011: data <= 13'h1fd9; 
        10'b0100001100: data <= 13'h1ff2; 
        10'b0100001101: data <= 13'h0002; 
        10'b0100001110: data <= 13'h0004; 
        10'b0100001111: data <= 13'h0008; 
        10'b0100010000: data <= 13'h000a; 
        10'b0100010001: data <= 13'h0009; 
        10'b0100010010: data <= 13'h0015; 
        10'b0100010011: data <= 13'h0015; 
        10'b0100010100: data <= 13'h1ffd; 
        10'b0100010101: data <= 13'h1ffd; 
        10'b0100010110: data <= 13'h0005; 
        10'b0100010111: data <= 13'h1ff9; 
        10'b0100011000: data <= 13'h1ffb; 
        10'b0100011001: data <= 13'h0000; 
        10'b0100011010: data <= 13'h1ffa; 
        10'b0100011011: data <= 13'h0001; 
        10'b0100011100: data <= 13'h0005; 
        10'b0100011101: data <= 13'h000f; 
        10'b0100011110: data <= 13'h000f; 
        10'b0100011111: data <= 13'h001c; 
        10'b0100100000: data <= 13'h0015; 
        10'b0100100001: data <= 13'h0018; 
        10'b0100100010: data <= 13'h0024; 
        10'b0100100011: data <= 13'h0011; 
        10'b0100100100: data <= 13'h0012; 
        10'b0100100101: data <= 13'h000f; 
        10'b0100100110: data <= 13'h1ffb; 
        10'b0100100111: data <= 13'h1fda; 
        10'b0100101000: data <= 13'h1fe1; 
        10'b0100101001: data <= 13'h1ff7; 
        10'b0100101010: data <= 13'h000b; 
        10'b0100101011: data <= 13'h000b; 
        10'b0100101100: data <= 13'h000b; 
        10'b0100101101: data <= 13'h0019; 
        10'b0100101110: data <= 13'h001c; 
        10'b0100101111: data <= 13'h0017; 
        10'b0100110000: data <= 13'h0000; 
        10'b0100110001: data <= 13'h1ffe; 
        10'b0100110010: data <= 13'h1ffd; 
        10'b0100110011: data <= 13'h1ffb; 
        10'b0100110100: data <= 13'h1ffa; 
        10'b0100110101: data <= 13'h0001; 
        10'b0100110110: data <= 13'h0000; 
        10'b0100110111: data <= 13'h1ff7; 
        10'b0100111000: data <= 13'h0007; 
        10'b0100111001: data <= 13'h0011; 
        10'b0100111010: data <= 13'h0021; 
        10'b0100111011: data <= 13'h002a; 
        10'b0100111100: data <= 13'h0021; 
        10'b0100111101: data <= 13'h002a; 
        10'b0100111110: data <= 13'h001d; 
        10'b0100111111: data <= 13'h000e; 
        10'b0101000000: data <= 13'h0011; 
        10'b0101000001: data <= 13'h002a; 
        10'b0101000010: data <= 13'h0033; 
        10'b0101000011: data <= 13'h1ffa; 
        10'b0101000100: data <= 13'h1fe2; 
        10'b0101000101: data <= 13'h1ff6; 
        10'b0101000110: data <= 13'h1ff6; 
        10'b0101000111: data <= 13'h0004; 
        10'b0101001000: data <= 13'h0017; 
        10'b0101001001: data <= 13'h001c; 
        10'b0101001010: data <= 13'h0025; 
        10'b0101001011: data <= 13'h0023; 
        10'b0101001100: data <= 13'h0018; 
        10'b0101001101: data <= 13'h0004; 
        10'b0101001110: data <= 13'h0002; 
        10'b0101001111: data <= 13'h1ffe; 
        10'b0101010000: data <= 13'h1ffb; 
        10'b0101010001: data <= 13'h1ffe; 
        10'b0101010010: data <= 13'h1ffc; 
        10'b0101010011: data <= 13'h1ffe; 
        10'b0101010100: data <= 13'h1ffe; 
        10'b0101010101: data <= 13'h0014; 
        10'b0101010110: data <= 13'h0011; 
        10'b0101010111: data <= 13'h001a; 
        10'b0101011000: data <= 13'h0018; 
        10'b0101011001: data <= 13'h001f; 
        10'b0101011010: data <= 13'h0005; 
        10'b0101011011: data <= 13'h0007; 
        10'b0101011100: data <= 13'h0004; 
        10'b0101011101: data <= 13'h0032; 
        10'b0101011110: data <= 13'h0033; 
        10'b0101011111: data <= 13'h000b; 
        10'b0101100000: data <= 13'h0002; 
        10'b0101100001: data <= 13'h1ffc; 
        10'b0101100010: data <= 13'h1ffc; 
        10'b0101100011: data <= 13'h000d; 
        10'b0101100100: data <= 13'h0016; 
        10'b0101100101: data <= 13'h0025; 
        10'b0101100110: data <= 13'h002b; 
        10'b0101100111: data <= 13'h0024; 
        10'b0101101000: data <= 13'h0017; 
        10'b0101101001: data <= 13'h0009; 
        10'b0101101010: data <= 13'h0004; 
        10'b0101101011: data <= 13'h1ffa; 
        10'b0101101100: data <= 13'h1ff9; 
        10'b0101101101: data <= 13'h1ffd; 
        10'b0101101110: data <= 13'h0001; 
        10'b0101101111: data <= 13'h1ffa; 
        10'b0101110000: data <= 13'h1ffb; 
        10'b0101110001: data <= 13'h0000; 
        10'b0101110010: data <= 13'h1ffd; 
        10'b0101110011: data <= 13'h1ffd; 
        10'b0101110100: data <= 13'h0003; 
        10'b0101110101: data <= 13'h1ffc; 
        10'b0101110110: data <= 13'h1ff5; 
        10'b0101110111: data <= 13'h0004; 
        10'b0101111000: data <= 13'h0013; 
        10'b0101111001: data <= 13'h002f; 
        10'b0101111010: data <= 13'h000e; 
        10'b0101111011: data <= 13'h0023; 
        10'b0101111100: data <= 13'h000e; 
        10'b0101111101: data <= 13'h1ff7; 
        10'b0101111110: data <= 13'h0001; 
        10'b0101111111: data <= 13'h0001; 
        10'b0110000000: data <= 13'h000f; 
        10'b0110000001: data <= 13'h000e; 
        10'b0110000010: data <= 13'h0008; 
        10'b0110000011: data <= 13'h000b; 
        10'b0110000100: data <= 13'h0006; 
        10'b0110000101: data <= 13'h0001; 
        10'b0110000110: data <= 13'h0001; 
        10'b0110000111: data <= 13'h1fff; 
        10'b0110001000: data <= 13'h1ffc; 
        10'b0110001001: data <= 13'h1ff9; 
        10'b0110001010: data <= 13'h1fff; 
        10'b0110001011: data <= 13'h1ffd; 
        10'b0110001100: data <= 13'h1ffa; 
        10'b0110001101: data <= 13'h1ff2; 
        10'b0110001110: data <= 13'h1fe8; 
        10'b0110001111: data <= 13'h1fe1; 
        10'b0110010000: data <= 13'h1fdb; 
        10'b0110010001: data <= 13'h1fe2; 
        10'b0110010010: data <= 13'h1ffc; 
        10'b0110010011: data <= 13'h0013; 
        10'b0110010100: data <= 13'h0012; 
        10'b0110010101: data <= 13'h0027; 
        10'b0110010110: data <= 13'h001f; 
        10'b0110010111: data <= 13'h0015; 
        10'b0110011000: data <= 13'h1ffd; 
        10'b0110011001: data <= 13'h0003; 
        10'b0110011010: data <= 13'h1ffb; 
        10'b0110011011: data <= 13'h1ff3; 
        10'b0110011100: data <= 13'h1fec; 
        10'b0110011101: data <= 13'h1fee; 
        10'b0110011110: data <= 13'h1ff0; 
        10'b0110011111: data <= 13'h1fed; 
        10'b0110100000: data <= 13'h1ff8; 
        10'b0110100001: data <= 13'h1fff; 
        10'b0110100010: data <= 13'h1ff8; 
        10'b0110100011: data <= 13'h0000; 
        10'b0110100100: data <= 13'h0001; 
        10'b0110100101: data <= 13'h1ffb; 
        10'b0110100110: data <= 13'h1ffb; 
        10'b0110100111: data <= 13'h1ffe; 
        10'b0110101000: data <= 13'h1ff9; 
        10'b0110101001: data <= 13'h1ff2; 
        10'b0110101010: data <= 13'h1fe1; 
        10'b0110101011: data <= 13'h1fdb; 
        10'b0110101100: data <= 13'h1fde; 
        10'b0110101101: data <= 13'h1ff8; 
        10'b0110101110: data <= 13'h0001; 
        10'b0110101111: data <= 13'h0001; 
        10'b0110110000: data <= 13'h001a; 
        10'b0110110001: data <= 13'h001f; 
        10'b0110110010: data <= 13'h001b; 
        10'b0110110011: data <= 13'h0010; 
        10'b0110110100: data <= 13'h1ff8; 
        10'b0110110101: data <= 13'h1ff9; 
        10'b0110110110: data <= 13'h1ffb; 
        10'b0110110111: data <= 13'h1fe4; 
        10'b0110111000: data <= 13'h1fde; 
        10'b0110111001: data <= 13'h1fe6; 
        10'b0110111010: data <= 13'h1fef; 
        10'b0110111011: data <= 13'h1ff0; 
        10'b0110111100: data <= 13'h1ff4; 
        10'b0110111101: data <= 13'h1ffe; 
        10'b0110111110: data <= 13'h1ff8; 
        10'b0110111111: data <= 13'h0001; 
        10'b0111000000: data <= 13'h1ffc; 
        10'b0111000001: data <= 13'h1ff9; 
        10'b0111000010: data <= 13'h1ffb; 
        10'b0111000011: data <= 13'h1ffe; 
        10'b0111000100: data <= 13'h1ff5; 
        10'b0111000101: data <= 13'h1fec; 
        10'b0111000110: data <= 13'h1fe0; 
        10'b0111000111: data <= 13'h1fed; 
        10'b0111001000: data <= 13'h000d; 
        10'b0111001001: data <= 13'h000e; 
        10'b0111001010: data <= 13'h0006; 
        10'b0111001011: data <= 13'h000d; 
        10'b0111001100: data <= 13'h0019; 
        10'b0111001101: data <= 13'h0016; 
        10'b0111001110: data <= 13'h0008; 
        10'b0111001111: data <= 13'h000d; 
        10'b0111010000: data <= 13'h0005; 
        10'b0111010001: data <= 13'h1ff6; 
        10'b0111010010: data <= 13'h1fea; 
        10'b0111010011: data <= 13'h1fe0; 
        10'b0111010100: data <= 13'h1fe0; 
        10'b0111010101: data <= 13'h1fe0; 
        10'b0111010110: data <= 13'h1fe6; 
        10'b0111010111: data <= 13'h1ff7; 
        10'b0111011000: data <= 13'h1ff5; 
        10'b0111011001: data <= 13'h1ffc; 
        10'b0111011010: data <= 13'h1ffc; 
        10'b0111011011: data <= 13'h1ff9; 
        10'b0111011100: data <= 13'h0002; 
        10'b0111011101: data <= 13'h0001; 
        10'b0111011110: data <= 13'h1ffb; 
        10'b0111011111: data <= 13'h1ff9; 
        10'b0111100000: data <= 13'h1ff9; 
        10'b0111100001: data <= 13'h1fec; 
        10'b0111100010: data <= 13'h1fe4; 
        10'b0111100011: data <= 13'h0005; 
        10'b0111100100: data <= 13'h001a; 
        10'b0111100101: data <= 13'h0020; 
        10'b0111100110: data <= 13'h000a; 
        10'b0111100111: data <= 13'h0018; 
        10'b0111101000: data <= 13'h0028; 
        10'b0111101001: data <= 13'h0018; 
        10'b0111101010: data <= 13'h0002; 
        10'b0111101011: data <= 13'h1ffa; 
        10'b0111101100: data <= 13'h0003; 
        10'b0111101101: data <= 13'h1ff4; 
        10'b0111101110: data <= 13'h1fdf; 
        10'b0111101111: data <= 13'h1ff0; 
        10'b0111110000: data <= 13'h1ff1; 
        10'b0111110001: data <= 13'h1fea; 
        10'b0111110010: data <= 13'h1ff0; 
        10'b0111110011: data <= 13'h1ff6; 
        10'b0111110100: data <= 13'h1ffa; 
        10'b0111110101: data <= 13'h1ff8; 
        10'b0111110110: data <= 13'h1fff; 
        10'b0111110111: data <= 13'h1ffc; 
        10'b0111111000: data <= 13'h1ffb; 
        10'b0111111001: data <= 13'h0000; 
        10'b0111111010: data <= 13'h1ff9; 
        10'b0111111011: data <= 13'h1ff7; 
        10'b0111111100: data <= 13'h1ff4; 
        10'b0111111101: data <= 13'h1ff3; 
        10'b0111111110: data <= 13'h1ff8; 
        10'b0111111111: data <= 13'h0008; 
        10'b1000000000: data <= 13'h0015; 
        10'b1000000001: data <= 13'h0027; 
        10'b1000000010: data <= 13'h001b; 
        10'b1000000011: data <= 13'h0025; 
        10'b1000000100: data <= 13'h0018; 
        10'b1000000101: data <= 13'h000e; 
        10'b1000000110: data <= 13'h1fef; 
        10'b1000000111: data <= 13'h1ffc; 
        10'b1000001000: data <= 13'h1ff7; 
        10'b1000001001: data <= 13'h1fe7; 
        10'b1000001010: data <= 13'h1ffa; 
        10'b1000001011: data <= 13'h1ffb; 
        10'b1000001100: data <= 13'h0002; 
        10'b1000001101: data <= 13'h1ff2; 
        10'b1000001110: data <= 13'h1ffe; 
        10'b1000001111: data <= 13'h1ff4; 
        10'b1000010000: data <= 13'h1ff0; 
        10'b1000010001: data <= 13'h1ff8; 
        10'b1000010010: data <= 13'h1fff; 
        10'b1000010011: data <= 13'h0001; 
        10'b1000010100: data <= 13'h1ffb; 
        10'b1000010101: data <= 13'h1ffe; 
        10'b1000010110: data <= 13'h1ffe; 
        10'b1000010111: data <= 13'h1ff5; 
        10'b1000011000: data <= 13'h1ff2; 
        10'b1000011001: data <= 13'h1ffa; 
        10'b1000011010: data <= 13'h0004; 
        10'b1000011011: data <= 13'h000a; 
        10'b1000011100: data <= 13'h000b; 
        10'b1000011101: data <= 13'h001a; 
        10'b1000011110: data <= 13'h000d; 
        10'b1000011111: data <= 13'h1ffe; 
        10'b1000100000: data <= 13'h0006; 
        10'b1000100001: data <= 13'h1fee; 
        10'b1000100010: data <= 13'h1fec; 
        10'b1000100011: data <= 13'h1ff8; 
        10'b1000100100: data <= 13'h1ffa; 
        10'b1000100101: data <= 13'h1ff8; 
        10'b1000100110: data <= 13'h0006; 
        10'b1000100111: data <= 13'h0002; 
        10'b1000101000: data <= 13'h0008; 
        10'b1000101001: data <= 13'h0001; 
        10'b1000101010: data <= 13'h0005; 
        10'b1000101011: data <= 13'h1ffb; 
        10'b1000101100: data <= 13'h1ff4; 
        10'b1000101101: data <= 13'h1ff9; 
        10'b1000101110: data <= 13'h1ffa; 
        10'b1000101111: data <= 13'h0001; 
        10'b1000110000: data <= 13'h1ffa; 
        10'b1000110001: data <= 13'h1fff; 
        10'b1000110010: data <= 13'h1ffb; 
        10'b1000110011: data <= 13'h1ff8; 
        10'b1000110100: data <= 13'h1ff0; 
        10'b1000110101: data <= 13'h1ffd; 
        10'b1000110110: data <= 13'h0003; 
        10'b1000110111: data <= 13'h0017; 
        10'b1000111000: data <= 13'h0007; 
        10'b1000111001: data <= 13'h1ffd; 
        10'b1000111010: data <= 13'h0000; 
        10'b1000111011: data <= 13'h1fed; 
        10'b1000111100: data <= 13'h0001; 
        10'b1000111101: data <= 13'h1fff; 
        10'b1000111110: data <= 13'h1fee; 
        10'b1000111111: data <= 13'h1ffd; 
        10'b1001000000: data <= 13'h1feb; 
        10'b1001000001: data <= 13'h1ff9; 
        10'b1001000010: data <= 13'h0004; 
        10'b1001000011: data <= 13'h0002; 
        10'b1001000100: data <= 13'h0007; 
        10'b1001000101: data <= 13'h000b; 
        10'b1001000110: data <= 13'h000b; 
        10'b1001000111: data <= 13'h1ffd; 
        10'b1001001000: data <= 13'h1ff9; 
        10'b1001001001: data <= 13'h1ff6; 
        10'b1001001010: data <= 13'h1ffd; 
        10'b1001001011: data <= 13'h1ffa; 
        10'b1001001100: data <= 13'h0001; 
        10'b1001001101: data <= 13'h1ffd; 
        10'b1001001110: data <= 13'h0001; 
        10'b1001001111: data <= 13'h1ff3; 
        10'b1001010000: data <= 13'h1fed; 
        10'b1001010001: data <= 13'h1ffe; 
        10'b1001010010: data <= 13'h000a; 
        10'b1001010011: data <= 13'h0015; 
        10'b1001010100: data <= 13'h0004; 
        10'b1001010101: data <= 13'h0009; 
        10'b1001010110: data <= 13'h1ffe; 
        10'b1001010111: data <= 13'h1ff2; 
        10'b1001011000: data <= 13'h1ff8; 
        10'b1001011001: data <= 13'h0005; 
        10'b1001011010: data <= 13'h0000; 
        10'b1001011011: data <= 13'h1ffe; 
        10'b1001011100: data <= 13'h1ff0; 
        10'b1001011101: data <= 13'h1ff9; 
        10'b1001011110: data <= 13'h1ffb; 
        10'b1001011111: data <= 13'h1fff; 
        10'b1001100000: data <= 13'h0000; 
        10'b1001100001: data <= 13'h0004; 
        10'b1001100010: data <= 13'h0003; 
        10'b1001100011: data <= 13'h1ffb; 
        10'b1001100100: data <= 13'h1ffa; 
        10'b1001100101: data <= 13'h0000; 
        10'b1001100110: data <= 13'h1fff; 
        10'b1001100111: data <= 13'h1ffc; 
        10'b1001101000: data <= 13'h1ffe; 
        10'b1001101001: data <= 13'h1ff9; 
        10'b1001101010: data <= 13'h1ffb; 
        10'b1001101011: data <= 13'h1ff8; 
        10'b1001101100: data <= 13'h1ff1; 
        10'b1001101101: data <= 13'h1fea; 
        10'b1001101110: data <= 13'h0003; 
        10'b1001101111: data <= 13'h0006; 
        10'b1001110000: data <= 13'h1fff; 
        10'b1001110001: data <= 13'h1ff9; 
        10'b1001110010: data <= 13'h0004; 
        10'b1001110011: data <= 13'h0002; 
        10'b1001110100: data <= 13'h001a; 
        10'b1001110101: data <= 13'h001c; 
        10'b1001110110: data <= 13'h0014; 
        10'b1001110111: data <= 13'h000f; 
        10'b1001111000: data <= 13'h1fff; 
        10'b1001111001: data <= 13'h1fff; 
        10'b1001111010: data <= 13'h0007; 
        10'b1001111011: data <= 13'h1ff8; 
        10'b1001111100: data <= 13'h1ff7; 
        10'b1001111101: data <= 13'h0004; 
        10'b1001111110: data <= 13'h1ffe; 
        10'b1001111111: data <= 13'h1ffa; 
        10'b1010000000: data <= 13'h1fff; 
        10'b1010000001: data <= 13'h1fff; 
        10'b1010000010: data <= 13'h1ffe; 
        10'b1010000011: data <= 13'h1ffb; 
        10'b1010000100: data <= 13'h1ffa; 
        10'b1010000101: data <= 13'h1fff; 
        10'b1010000110: data <= 13'h1ffd; 
        10'b1010000111: data <= 13'h1ff9; 
        10'b1010001000: data <= 13'h1ff0; 
        10'b1010001001: data <= 13'h1fdb; 
        10'b1010001010: data <= 13'h1fe3; 
        10'b1010001011: data <= 13'h1ff1; 
        10'b1010001100: data <= 13'h0005; 
        10'b1010001101: data <= 13'h0005; 
        10'b1010001110: data <= 13'h000b; 
        10'b1010001111: data <= 13'h000e; 
        10'b1010010000: data <= 13'h001f; 
        10'b1010010001: data <= 13'h002d; 
        10'b1010010010: data <= 13'h0026; 
        10'b1010010011: data <= 13'h001f; 
        10'b1010010100: data <= 13'h0019; 
        10'b1010010101: data <= 13'h0012; 
        10'b1010010110: data <= 13'h000e; 
        10'b1010010111: data <= 13'h0012; 
        10'b1010011000: data <= 13'h000d; 
        10'b1010011001: data <= 13'h0003; 
        10'b1010011010: data <= 13'h1ffe; 
        10'b1010011011: data <= 13'h1ffc; 
        10'b1010011100: data <= 13'h1ff8; 
        10'b1010011101: data <= 13'h1fff; 
        10'b1010011110: data <= 13'h1ff9; 
        10'b1010011111: data <= 13'h1fff; 
        10'b1010100000: data <= 13'h1fff; 
        10'b1010100001: data <= 13'h1fff; 
        10'b1010100010: data <= 13'h0001; 
        10'b1010100011: data <= 13'h1ffa; 
        10'b1010100100: data <= 13'h1ffa; 
        10'b1010100101: data <= 13'h1fe8; 
        10'b1010100110: data <= 13'h1fde; 
        10'b1010100111: data <= 13'h1fe3; 
        10'b1010101000: data <= 13'h1ffe; 
        10'b1010101001: data <= 13'h0007; 
        10'b1010101010: data <= 13'h1ffd; 
        10'b1010101011: data <= 13'h000c; 
        10'b1010101100: data <= 13'h0009; 
        10'b1010101101: data <= 13'h0006; 
        10'b1010101110: data <= 13'h000f; 
        10'b1010101111: data <= 13'h0020; 
        10'b1010110000: data <= 13'h0022; 
        10'b1010110001: data <= 13'h0017; 
        10'b1010110010: data <= 13'h0020; 
        10'b1010110011: data <= 13'h001e; 
        10'b1010110100: data <= 13'h000a; 
        10'b1010110101: data <= 13'h0001; 
        10'b1010110110: data <= 13'h1ff9; 
        10'b1010110111: data <= 13'h0001; 
        10'b1010111000: data <= 13'h1ffd; 
        10'b1010111001: data <= 13'h1ffb; 
        10'b1010111010: data <= 13'h0001; 
        10'b1010111011: data <= 13'h1ffe; 
        10'b1010111100: data <= 13'h0001; 
        10'b1010111101: data <= 13'h1fff; 
        10'b1010111110: data <= 13'h0001; 
        10'b1010111111: data <= 13'h1ffa; 
        10'b1011000000: data <= 13'h1ffb; 
        10'b1011000001: data <= 13'h1ff7; 
        10'b1011000010: data <= 13'h1ff3; 
        10'b1011000011: data <= 13'h1ff0; 
        10'b1011000100: data <= 13'h1fee; 
        10'b1011000101: data <= 13'h1fee; 
        10'b1011000110: data <= 13'h1ff9; 
        10'b1011000111: data <= 13'h1ff3; 
        10'b1011001000: data <= 13'h1ff9; 
        10'b1011001001: data <= 13'h1ff8; 
        10'b1011001010: data <= 13'h1fff; 
        10'b1011001011: data <= 13'h000b; 
        10'b1011001100: data <= 13'h0008; 
        10'b1011001101: data <= 13'h000a; 
        10'b1011001110: data <= 13'h000c; 
        10'b1011001111: data <= 13'h0002; 
        10'b1011010000: data <= 13'h1ffe; 
        10'b1011010001: data <= 13'h0000; 
        10'b1011010010: data <= 13'h1ff8; 
        10'b1011010011: data <= 13'h1ff9; 
        10'b1011010100: data <= 13'h1fff; 
        10'b1011010101: data <= 13'h1ffe; 
        10'b1011010110: data <= 13'h1ffb; 
        10'b1011010111: data <= 13'h1ffe; 
        10'b1011011000: data <= 13'h1fff; 
        10'b1011011001: data <= 13'h0000; 
        10'b1011011010: data <= 13'h1ffc; 
        10'b1011011011: data <= 13'h1ffb; 
        10'b1011011100: data <= 13'h1ff8; 
        10'b1011011101: data <= 13'h1ffa; 
        10'b1011011110: data <= 13'h1ff6; 
        10'b1011011111: data <= 13'h1ffd; 
        10'b1011100000: data <= 13'h1ff7; 
        10'b1011100001: data <= 13'h1ff8; 
        10'b1011100010: data <= 13'h1ff7; 
        10'b1011100011: data <= 13'h1ffb; 
        10'b1011100100: data <= 13'h1ffa; 
        10'b1011100101: data <= 13'h1ffb; 
        10'b1011100110: data <= 13'h1ff9; 
        10'b1011100111: data <= 13'h1ffb; 
        10'b1011101000: data <= 13'h1ffa; 
        10'b1011101001: data <= 13'h1ff8; 
        10'b1011101010: data <= 13'h1ff7; 
        10'b1011101011: data <= 13'h1ffa; 
        10'b1011101100: data <= 13'h1ffc; 
        10'b1011101101: data <= 13'h1fff; 
        10'b1011101110: data <= 13'h1ffc; 
        10'b1011101111: data <= 13'h0002; 
        10'b1011110000: data <= 13'h0002; 
        10'b1011110001: data <= 13'h1ff9; 
        10'b1011110010: data <= 13'h1ffe; 
        10'b1011110011: data <= 13'h1ffd; 
        10'b1011110100: data <= 13'h1ffe; 
        10'b1011110101: data <= 13'h1ffb; 
        10'b1011110110: data <= 13'h1ffd; 
        10'b1011110111: data <= 13'h1ffe; 
        10'b1011111000: data <= 13'h1ffe; 
        10'b1011111001: data <= 13'h1ff9; 
        10'b1011111010: data <= 13'h0000; 
        10'b1011111011: data <= 13'h1ffb; 
        10'b1011111100: data <= 13'h0001; 
        10'b1011111101: data <= 13'h1ffc; 
        10'b1011111110: data <= 13'h1ffa; 
        10'b1011111111: data <= 13'h1fff; 
        10'b1100000000: data <= 13'h1ffb; 
        10'b1100000001: data <= 13'h1ffa; 
        10'b1100000010: data <= 13'h1ffc; 
        10'b1100000011: data <= 13'h1ffe; 
        10'b1100000100: data <= 13'h1ffe; 
        10'b1100000101: data <= 13'h0000; 
        10'b1100000110: data <= 13'h0001; 
        10'b1100000111: data <= 13'h0001; 
        10'b1100001000: data <= 13'h1fff; 
        10'b1100001001: data <= 13'h1ffe; 
        10'b1100001010: data <= 13'h1fff; 
        10'b1100001011: data <= 13'h1ffa; 
        10'b1100001100: data <= 13'h1ffd; 
        10'b1100001101: data <= 13'h0001; 
        10'b1100001110: data <= 13'h1ff9; 
        10'b1100001111: data <= 13'h1ffd; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 8) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 14'h3ff9; 
        10'b0000000001: data <= 14'h3ffa; 
        10'b0000000010: data <= 14'h3ff9; 
        10'b0000000011: data <= 14'h3ffd; 
        10'b0000000100: data <= 14'h3ffc; 
        10'b0000000101: data <= 14'h0001; 
        10'b0000000110: data <= 14'h3ff1; 
        10'b0000000111: data <= 14'h3ffd; 
        10'b0000001000: data <= 14'h3ff6; 
        10'b0000001001: data <= 14'h3ff8; 
        10'b0000001010: data <= 14'h3ff4; 
        10'b0000001011: data <= 14'h0001; 
        10'b0000001100: data <= 14'h3ffb; 
        10'b0000001101: data <= 14'h3fff; 
        10'b0000001110: data <= 14'h3ff4; 
        10'b0000001111: data <= 14'h3fff; 
        10'b0000010000: data <= 14'h3ffc; 
        10'b0000010001: data <= 14'h3ff3; 
        10'b0000010010: data <= 14'h0001; 
        10'b0000010011: data <= 14'h3ffa; 
        10'b0000010100: data <= 14'h3ff9; 
        10'b0000010101: data <= 14'h3ff9; 
        10'b0000010110: data <= 14'h3ffa; 
        10'b0000010111: data <= 14'h0003; 
        10'b0000011000: data <= 14'h0000; 
        10'b0000011001: data <= 14'h3ff8; 
        10'b0000011010: data <= 14'h3ff6; 
        10'b0000011011: data <= 14'h3ff9; 
        10'b0000011100: data <= 14'h3ff9; 
        10'b0000011101: data <= 14'h3ff1; 
        10'b0000011110: data <= 14'h0002; 
        10'b0000011111: data <= 14'h0000; 
        10'b0000100000: data <= 14'h3ff3; 
        10'b0000100001: data <= 14'h3ff3; 
        10'b0000100010: data <= 14'h3ff2; 
        10'b0000100011: data <= 14'h3ff3; 
        10'b0000100100: data <= 14'h0002; 
        10'b0000100101: data <= 14'h3ffb; 
        10'b0000100110: data <= 14'h3ffa; 
        10'b0000100111: data <= 14'h3ff1; 
        10'b0000101000: data <= 14'h0002; 
        10'b0000101001: data <= 14'h3ffe; 
        10'b0000101010: data <= 14'h3ff6; 
        10'b0000101011: data <= 14'h3ff8; 
        10'b0000101100: data <= 14'h3ffe; 
        10'b0000101101: data <= 14'h3ffb; 
        10'b0000101110: data <= 14'h3ff5; 
        10'b0000101111: data <= 14'h3ffc; 
        10'b0000110000: data <= 14'h0001; 
        10'b0000110001: data <= 14'h3ff2; 
        10'b0000110010: data <= 14'h3ffe; 
        10'b0000110011: data <= 14'h3ff5; 
        10'b0000110100: data <= 14'h3fff; 
        10'b0000110101: data <= 14'h0003; 
        10'b0000110110: data <= 14'h3ff6; 
        10'b0000110111: data <= 14'h3ff5; 
        10'b0000111000: data <= 14'h3ff4; 
        10'b0000111001: data <= 14'h0000; 
        10'b0000111010: data <= 14'h3ffb; 
        10'b0000111011: data <= 14'h3ffa; 
        10'b0000111100: data <= 14'h3ff4; 
        10'b0000111101: data <= 14'h3ff2; 
        10'b0000111110: data <= 14'h3ffb; 
        10'b0000111111: data <= 14'h3ff1; 
        10'b0001000000: data <= 14'h0003; 
        10'b0001000001: data <= 14'h3ff1; 
        10'b0001000010: data <= 14'h3ff2; 
        10'b0001000011: data <= 14'h3ffd; 
        10'b0001000100: data <= 14'h3ffb; 
        10'b0001000101: data <= 14'h3ff1; 
        10'b0001000110: data <= 14'h3ffd; 
        10'b0001000111: data <= 14'h3ffc; 
        10'b0001001000: data <= 14'h3ff0; 
        10'b0001001001: data <= 14'h3ff7; 
        10'b0001001010: data <= 14'h3ff7; 
        10'b0001001011: data <= 14'h3ffe; 
        10'b0001001100: data <= 14'h0000; 
        10'b0001001101: data <= 14'h3fff; 
        10'b0001001110: data <= 14'h3ffc; 
        10'b0001001111: data <= 14'h3ff9; 
        10'b0001010000: data <= 14'h0001; 
        10'b0001010001: data <= 14'h3ff6; 
        10'b0001010010: data <= 14'h3ffe; 
        10'b0001010011: data <= 14'h0002; 
        10'b0001010100: data <= 14'h3ff5; 
        10'b0001010101: data <= 14'h3ffa; 
        10'b0001010110: data <= 14'h3ffa; 
        10'b0001010111: data <= 14'h3ff3; 
        10'b0001011000: data <= 14'h0003; 
        10'b0001011001: data <= 14'h3ff4; 
        10'b0001011010: data <= 14'h3ff2; 
        10'b0001011011: data <= 14'h3ff8; 
        10'b0001011100: data <= 14'h3ff2; 
        10'b0001011101: data <= 14'h3ffb; 
        10'b0001011110: data <= 14'h3ff5; 
        10'b0001011111: data <= 14'h3fec; 
        10'b0001100000: data <= 14'h3fea; 
        10'b0001100001: data <= 14'h3fe5; 
        10'b0001100010: data <= 14'h3fe9; 
        10'b0001100011: data <= 14'h3ff3; 
        10'b0001100100: data <= 14'h3fe9; 
        10'b0001100101: data <= 14'h3fee; 
        10'b0001100110: data <= 14'h3ff4; 
        10'b0001100111: data <= 14'h3ff9; 
        10'b0001101000: data <= 14'h3fef; 
        10'b0001101001: data <= 14'h0001; 
        10'b0001101010: data <= 14'h3ff7; 
        10'b0001101011: data <= 14'h3fff; 
        10'b0001101100: data <= 14'h3ff6; 
        10'b0001101101: data <= 14'h3ffd; 
        10'b0001101110: data <= 14'h3ffb; 
        10'b0001101111: data <= 14'h3ff3; 
        10'b0001110000: data <= 14'h3ffa; 
        10'b0001110001: data <= 14'h3ffe; 
        10'b0001110010: data <= 14'h3ff8; 
        10'b0001110011: data <= 14'h3ff3; 
        10'b0001110100: data <= 14'h3fff; 
        10'b0001110101: data <= 14'h3fff; 
        10'b0001110110: data <= 14'h3ffa; 
        10'b0001110111: data <= 14'h3ff4; 
        10'b0001111000: data <= 14'h3ff4; 
        10'b0001111001: data <= 14'h3ff9; 
        10'b0001111010: data <= 14'h3ffa; 
        10'b0001111011: data <= 14'h3ffd; 
        10'b0001111100: data <= 14'h0013; 
        10'b0001111101: data <= 14'h000d; 
        10'b0001111110: data <= 14'h002a; 
        10'b0001111111: data <= 14'h0020; 
        10'b0010000000: data <= 14'h000f; 
        10'b0010000001: data <= 14'h0008; 
        10'b0010000010: data <= 14'h000c; 
        10'b0010000011: data <= 14'h3ff5; 
        10'b0010000100: data <= 14'h3ff3; 
        10'b0010000101: data <= 14'h3ff9; 
        10'b0010000110: data <= 14'h3fec; 
        10'b0010000111: data <= 14'h3ff2; 
        10'b0010001000: data <= 14'h0000; 
        10'b0010001001: data <= 14'h0001; 
        10'b0010001010: data <= 14'h3ff8; 
        10'b0010001011: data <= 14'h3ffa; 
        10'b0010001100: data <= 14'h3ffa; 
        10'b0010001101: data <= 14'h3ffd; 
        10'b0010001110: data <= 14'h3ffe; 
        10'b0010001111: data <= 14'h3fff; 
        10'b0010010000: data <= 14'h3ff4; 
        10'b0010010001: data <= 14'h3ff9; 
        10'b0010010010: data <= 14'h3ff6; 
        10'b0010010011: data <= 14'h3fe5; 
        10'b0010010100: data <= 14'h3ff5; 
        10'b0010010101: data <= 14'h000a; 
        10'b0010010110: data <= 14'h3fea; 
        10'b0010010111: data <= 14'h001e; 
        10'b0010011000: data <= 14'h0038; 
        10'b0010011001: data <= 14'h002e; 
        10'b0010011010: data <= 14'h0030; 
        10'b0010011011: data <= 14'h0017; 
        10'b0010011100: data <= 14'h0013; 
        10'b0010011101: data <= 14'h002d; 
        10'b0010011110: data <= 14'h0002; 
        10'b0010011111: data <= 14'h3ffe; 
        10'b0010100000: data <= 14'h0010; 
        10'b0010100001: data <= 14'h0008; 
        10'b0010100010: data <= 14'h3fe5; 
        10'b0010100011: data <= 14'h3fe9; 
        10'b0010100100: data <= 14'h3ff0; 
        10'b0010100101: data <= 14'h000c; 
        10'b0010100110: data <= 14'h3ffb; 
        10'b0010100111: data <= 14'h0002; 
        10'b0010101000: data <= 14'h3ff5; 
        10'b0010101001: data <= 14'h3ff4; 
        10'b0010101010: data <= 14'h3ff2; 
        10'b0010101011: data <= 14'h3ff2; 
        10'b0010101100: data <= 14'h3ff0; 
        10'b0010101101: data <= 14'h3ff0; 
        10'b0010101110: data <= 14'h3fe7; 
        10'b0010101111: data <= 14'h3fe6; 
        10'b0010110000: data <= 14'h0002; 
        10'b0010110001: data <= 14'h0008; 
        10'b0010110010: data <= 14'h3ffe; 
        10'b0010110011: data <= 14'h000e; 
        10'b0010110100: data <= 14'h0017; 
        10'b0010110101: data <= 14'h0012; 
        10'b0010110110: data <= 14'h001a; 
        10'b0010110111: data <= 14'h0030; 
        10'b0010111000: data <= 14'h0017; 
        10'b0010111001: data <= 14'h001b; 
        10'b0010111010: data <= 14'h0006; 
        10'b0010111011: data <= 14'h001f; 
        10'b0010111100: data <= 14'h000c; 
        10'b0010111101: data <= 14'h000f; 
        10'b0010111110: data <= 14'h0012; 
        10'b0010111111: data <= 14'h0011; 
        10'b0011000000: data <= 14'h000e; 
        10'b0011000001: data <= 14'h0006; 
        10'b0011000010: data <= 14'h3ffa; 
        10'b0011000011: data <= 14'h3fff; 
        10'b0011000100: data <= 14'h0002; 
        10'b0011000101: data <= 14'h3ff5; 
        10'b0011000110: data <= 14'h3ff3; 
        10'b0011000111: data <= 14'h3ff6; 
        10'b0011001000: data <= 14'h3fef; 
        10'b0011001001: data <= 14'h3ffa; 
        10'b0011001010: data <= 14'h3fef; 
        10'b0011001011: data <= 14'h3fff; 
        10'b0011001100: data <= 14'h0011; 
        10'b0011001101: data <= 14'h0007; 
        10'b0011001110: data <= 14'h0009; 
        10'b0011001111: data <= 14'h3ffb; 
        10'b0011010000: data <= 14'h3fea; 
        10'b0011010001: data <= 14'h3ff0; 
        10'b0011010010: data <= 14'h3fe8; 
        10'b0011010011: data <= 14'h000f; 
        10'b0011010100: data <= 14'h0012; 
        10'b0011010101: data <= 14'h3fff; 
        10'b0011010110: data <= 14'h000c; 
        10'b0011010111: data <= 14'h3ff2; 
        10'b0011011000: data <= 14'h0013; 
        10'b0011011001: data <= 14'h001d; 
        10'b0011011010: data <= 14'h0005; 
        10'b0011011011: data <= 14'h003c; 
        10'b0011011100: data <= 14'h0025; 
        10'b0011011101: data <= 14'h3fff; 
        10'b0011011110: data <= 14'h0001; 
        10'b0011011111: data <= 14'h3ffd; 
        10'b0011100000: data <= 14'h3ffd; 
        10'b0011100001: data <= 14'h0001; 
        10'b0011100010: data <= 14'h3ffd; 
        10'b0011100011: data <= 14'h3ff4; 
        10'b0011100100: data <= 14'h3ffd; 
        10'b0011100101: data <= 14'h3ffa; 
        10'b0011100110: data <= 14'h0019; 
        10'b0011100111: data <= 14'h000f; 
        10'b0011101000: data <= 14'h0006; 
        10'b0011101001: data <= 14'h002b; 
        10'b0011101010: data <= 14'h0002; 
        10'b0011101011: data <= 14'h0001; 
        10'b0011101100: data <= 14'h001d; 
        10'b0011101101: data <= 14'h0025; 
        10'b0011101110: data <= 14'h3fe3; 
        10'b0011101111: data <= 14'h3fe7; 
        10'b0011110000: data <= 14'h0014; 
        10'b0011110001: data <= 14'h3ff2; 
        10'b0011110010: data <= 14'h0007; 
        10'b0011110011: data <= 14'h0014; 
        10'b0011110100: data <= 14'h000d; 
        10'b0011110101: data <= 14'h0028; 
        10'b0011110110: data <= 14'h001b; 
        10'b0011110111: data <= 14'h002d; 
        10'b0011111000: data <= 14'h0029; 
        10'b0011111001: data <= 14'h3ffb; 
        10'b0011111010: data <= 14'h3ffc; 
        10'b0011111011: data <= 14'h0004; 
        10'b0011111100: data <= 14'h0000; 
        10'b0011111101: data <= 14'h0001; 
        10'b0011111110: data <= 14'h3ffa; 
        10'b0011111111: data <= 14'h3ff8; 
        10'b0100000000: data <= 14'h3ffc; 
        10'b0100000001: data <= 14'h0019; 
        10'b0100000010: data <= 14'h0013; 
        10'b0100000011: data <= 14'h0027; 
        10'b0100000100: data <= 14'h0034; 
        10'b0100000101: data <= 14'h002c; 
        10'b0100000110: data <= 14'h001c; 
        10'b0100000111: data <= 14'h0031; 
        10'b0100001000: data <= 14'h000d; 
        10'b0100001001: data <= 14'h000e; 
        10'b0100001010: data <= 14'h3fc7; 
        10'b0100001011: data <= 14'h3fb1; 
        10'b0100001100: data <= 14'h3fe4; 
        10'b0100001101: data <= 14'h0004; 
        10'b0100001110: data <= 14'h0009; 
        10'b0100001111: data <= 14'h000f; 
        10'b0100010000: data <= 14'h0014; 
        10'b0100010001: data <= 14'h0011; 
        10'b0100010010: data <= 14'h002a; 
        10'b0100010011: data <= 14'h002b; 
        10'b0100010100: data <= 14'h3ff9; 
        10'b0100010101: data <= 14'h3ffa; 
        10'b0100010110: data <= 14'h000a; 
        10'b0100010111: data <= 14'h3ff3; 
        10'b0100011000: data <= 14'h3ff6; 
        10'b0100011001: data <= 14'h0000; 
        10'b0100011010: data <= 14'h3ff5; 
        10'b0100011011: data <= 14'h0001; 
        10'b0100011100: data <= 14'h000a; 
        10'b0100011101: data <= 14'h001f; 
        10'b0100011110: data <= 14'h001f; 
        10'b0100011111: data <= 14'h0038; 
        10'b0100100000: data <= 14'h002a; 
        10'b0100100001: data <= 14'h0031; 
        10'b0100100010: data <= 14'h0047; 
        10'b0100100011: data <= 14'h0022; 
        10'b0100100100: data <= 14'h0024; 
        10'b0100100101: data <= 14'h001d; 
        10'b0100100110: data <= 14'h3ff7; 
        10'b0100100111: data <= 14'h3fb5; 
        10'b0100101000: data <= 14'h3fc2; 
        10'b0100101001: data <= 14'h3fed; 
        10'b0100101010: data <= 14'h0015; 
        10'b0100101011: data <= 14'h0015; 
        10'b0100101100: data <= 14'h0016; 
        10'b0100101101: data <= 14'h0033; 
        10'b0100101110: data <= 14'h0038; 
        10'b0100101111: data <= 14'h002e; 
        10'b0100110000: data <= 14'h0001; 
        10'b0100110001: data <= 14'h3ffd; 
        10'b0100110010: data <= 14'h3ffa; 
        10'b0100110011: data <= 14'h3ff6; 
        10'b0100110100: data <= 14'h3ff5; 
        10'b0100110101: data <= 14'h0003; 
        10'b0100110110: data <= 14'h3fff; 
        10'b0100110111: data <= 14'h3fef; 
        10'b0100111000: data <= 14'h000f; 
        10'b0100111001: data <= 14'h0022; 
        10'b0100111010: data <= 14'h0041; 
        10'b0100111011: data <= 14'h0054; 
        10'b0100111100: data <= 14'h0042; 
        10'b0100111101: data <= 14'h0054; 
        10'b0100111110: data <= 14'h0039; 
        10'b0100111111: data <= 14'h001b; 
        10'b0101000000: data <= 14'h0023; 
        10'b0101000001: data <= 14'h0053; 
        10'b0101000010: data <= 14'h0066; 
        10'b0101000011: data <= 14'h3ff3; 
        10'b0101000100: data <= 14'h3fc3; 
        10'b0101000101: data <= 14'h3feb; 
        10'b0101000110: data <= 14'h3fec; 
        10'b0101000111: data <= 14'h0008; 
        10'b0101001000: data <= 14'h002e; 
        10'b0101001001: data <= 14'h0037; 
        10'b0101001010: data <= 14'h0049; 
        10'b0101001011: data <= 14'h0045; 
        10'b0101001100: data <= 14'h0030; 
        10'b0101001101: data <= 14'h0008; 
        10'b0101001110: data <= 14'h0004; 
        10'b0101001111: data <= 14'h3ffc; 
        10'b0101010000: data <= 14'h3ff6; 
        10'b0101010001: data <= 14'h3ffd; 
        10'b0101010010: data <= 14'h3ff8; 
        10'b0101010011: data <= 14'h3ffc; 
        10'b0101010100: data <= 14'h3ffd; 
        10'b0101010101: data <= 14'h0029; 
        10'b0101010110: data <= 14'h0022; 
        10'b0101010111: data <= 14'h0034; 
        10'b0101011000: data <= 14'h0031; 
        10'b0101011001: data <= 14'h003d; 
        10'b0101011010: data <= 14'h000a; 
        10'b0101011011: data <= 14'h000f; 
        10'b0101011100: data <= 14'h0008; 
        10'b0101011101: data <= 14'h0065; 
        10'b0101011110: data <= 14'h0065; 
        10'b0101011111: data <= 14'h0017; 
        10'b0101100000: data <= 14'h0004; 
        10'b0101100001: data <= 14'h3ff7; 
        10'b0101100010: data <= 14'h3ff9; 
        10'b0101100011: data <= 14'h0019; 
        10'b0101100100: data <= 14'h002b; 
        10'b0101100101: data <= 14'h004a; 
        10'b0101100110: data <= 14'h0056; 
        10'b0101100111: data <= 14'h0048; 
        10'b0101101000: data <= 14'h002d; 
        10'b0101101001: data <= 14'h0012; 
        10'b0101101010: data <= 14'h0009; 
        10'b0101101011: data <= 14'h3ff3; 
        10'b0101101100: data <= 14'h3ff2; 
        10'b0101101101: data <= 14'h3ffb; 
        10'b0101101110: data <= 14'h0003; 
        10'b0101101111: data <= 14'h3ff4; 
        10'b0101110000: data <= 14'h3ff7; 
        10'b0101110001: data <= 14'h0000; 
        10'b0101110010: data <= 14'h3ff9; 
        10'b0101110011: data <= 14'h3ffa; 
        10'b0101110100: data <= 14'h0006; 
        10'b0101110101: data <= 14'h3ff9; 
        10'b0101110110: data <= 14'h3fea; 
        10'b0101110111: data <= 14'h0008; 
        10'b0101111000: data <= 14'h0025; 
        10'b0101111001: data <= 14'h005e; 
        10'b0101111010: data <= 14'h001c; 
        10'b0101111011: data <= 14'h0045; 
        10'b0101111100: data <= 14'h001c; 
        10'b0101111101: data <= 14'h3fee; 
        10'b0101111110: data <= 14'h0002; 
        10'b0101111111: data <= 14'h0002; 
        10'b0110000000: data <= 14'h001f; 
        10'b0110000001: data <= 14'h001c; 
        10'b0110000010: data <= 14'h0010; 
        10'b0110000011: data <= 14'h0017; 
        10'b0110000100: data <= 14'h000c; 
        10'b0110000101: data <= 14'h0003; 
        10'b0110000110: data <= 14'h0003; 
        10'b0110000111: data <= 14'h3ffe; 
        10'b0110001000: data <= 14'h3ff7; 
        10'b0110001001: data <= 14'h3ff2; 
        10'b0110001010: data <= 14'h3ffe; 
        10'b0110001011: data <= 14'h3ffa; 
        10'b0110001100: data <= 14'h3ff3; 
        10'b0110001101: data <= 14'h3fe5; 
        10'b0110001110: data <= 14'h3fcf; 
        10'b0110001111: data <= 14'h3fc1; 
        10'b0110010000: data <= 14'h3fb6; 
        10'b0110010001: data <= 14'h3fc5; 
        10'b0110010010: data <= 14'h3ff8; 
        10'b0110010011: data <= 14'h0026; 
        10'b0110010100: data <= 14'h0025; 
        10'b0110010101: data <= 14'h004d; 
        10'b0110010110: data <= 14'h003e; 
        10'b0110010111: data <= 14'h002a; 
        10'b0110011000: data <= 14'h3ffb; 
        10'b0110011001: data <= 14'h0005; 
        10'b0110011010: data <= 14'h3ff5; 
        10'b0110011011: data <= 14'h3fe7; 
        10'b0110011100: data <= 14'h3fd7; 
        10'b0110011101: data <= 14'h3fdb; 
        10'b0110011110: data <= 14'h3fe0; 
        10'b0110011111: data <= 14'h3fdb; 
        10'b0110100000: data <= 14'h3fef; 
        10'b0110100001: data <= 14'h3ffe; 
        10'b0110100010: data <= 14'h3ff1; 
        10'b0110100011: data <= 14'h0000; 
        10'b0110100100: data <= 14'h0001; 
        10'b0110100101: data <= 14'h3ff7; 
        10'b0110100110: data <= 14'h3ff5; 
        10'b0110100111: data <= 14'h3ffc; 
        10'b0110101000: data <= 14'h3ff2; 
        10'b0110101001: data <= 14'h3fe5; 
        10'b0110101010: data <= 14'h3fc3; 
        10'b0110101011: data <= 14'h3fb5; 
        10'b0110101100: data <= 14'h3fbc; 
        10'b0110101101: data <= 14'h3fef; 
        10'b0110101110: data <= 14'h0003; 
        10'b0110101111: data <= 14'h0002; 
        10'b0110110000: data <= 14'h0035; 
        10'b0110110001: data <= 14'h003e; 
        10'b0110110010: data <= 14'h0037; 
        10'b0110110011: data <= 14'h001f; 
        10'b0110110100: data <= 14'h3ff0; 
        10'b0110110101: data <= 14'h3ff2; 
        10'b0110110110: data <= 14'h3ff6; 
        10'b0110110111: data <= 14'h3fc9; 
        10'b0110111000: data <= 14'h3fbb; 
        10'b0110111001: data <= 14'h3fcb; 
        10'b0110111010: data <= 14'h3fdf; 
        10'b0110111011: data <= 14'h3fe0; 
        10'b0110111100: data <= 14'h3fe8; 
        10'b0110111101: data <= 14'h3ffc; 
        10'b0110111110: data <= 14'h3fef; 
        10'b0110111111: data <= 14'h0001; 
        10'b0111000000: data <= 14'h3ff9; 
        10'b0111000001: data <= 14'h3ff2; 
        10'b0111000010: data <= 14'h3ff7; 
        10'b0111000011: data <= 14'h3ffb; 
        10'b0111000100: data <= 14'h3fea; 
        10'b0111000101: data <= 14'h3fd9; 
        10'b0111000110: data <= 14'h3fc1; 
        10'b0111000111: data <= 14'h3fdb; 
        10'b0111001000: data <= 14'h0019; 
        10'b0111001001: data <= 14'h001c; 
        10'b0111001010: data <= 14'h000b; 
        10'b0111001011: data <= 14'h001a; 
        10'b0111001100: data <= 14'h0033; 
        10'b0111001101: data <= 14'h002d; 
        10'b0111001110: data <= 14'h0010; 
        10'b0111001111: data <= 14'h001b; 
        10'b0111010000: data <= 14'h0009; 
        10'b0111010001: data <= 14'h3feb; 
        10'b0111010010: data <= 14'h3fd3; 
        10'b0111010011: data <= 14'h3fc0; 
        10'b0111010100: data <= 14'h3fc0; 
        10'b0111010101: data <= 14'h3fbf; 
        10'b0111010110: data <= 14'h3fcc; 
        10'b0111010111: data <= 14'h3fef; 
        10'b0111011000: data <= 14'h3fe9; 
        10'b0111011001: data <= 14'h3ff8; 
        10'b0111011010: data <= 14'h3ff8; 
        10'b0111011011: data <= 14'h3ff2; 
        10'b0111011100: data <= 14'h0003; 
        10'b0111011101: data <= 14'h0002; 
        10'b0111011110: data <= 14'h3ff5; 
        10'b0111011111: data <= 14'h3ff3; 
        10'b0111100000: data <= 14'h3ff1; 
        10'b0111100001: data <= 14'h3fd7; 
        10'b0111100010: data <= 14'h3fc8; 
        10'b0111100011: data <= 14'h000a; 
        10'b0111100100: data <= 14'h0034; 
        10'b0111100101: data <= 14'h0040; 
        10'b0111100110: data <= 14'h0015; 
        10'b0111100111: data <= 14'h0031; 
        10'b0111101000: data <= 14'h004f; 
        10'b0111101001: data <= 14'h0030; 
        10'b0111101010: data <= 14'h0004; 
        10'b0111101011: data <= 14'h3ff3; 
        10'b0111101100: data <= 14'h0006; 
        10'b0111101101: data <= 14'h3fe7; 
        10'b0111101110: data <= 14'h3fbf; 
        10'b0111101111: data <= 14'h3fe1; 
        10'b0111110000: data <= 14'h3fe1; 
        10'b0111110001: data <= 14'h3fd5; 
        10'b0111110010: data <= 14'h3fe0; 
        10'b0111110011: data <= 14'h3fec; 
        10'b0111110100: data <= 14'h3ff4; 
        10'b0111110101: data <= 14'h3fef; 
        10'b0111110110: data <= 14'h3ffd; 
        10'b0111110111: data <= 14'h3ff7; 
        10'b0111111000: data <= 14'h3ff6; 
        10'b0111111001: data <= 14'h0001; 
        10'b0111111010: data <= 14'h3ff2; 
        10'b0111111011: data <= 14'h3fee; 
        10'b0111111100: data <= 14'h3fe7; 
        10'b0111111101: data <= 14'h3fe6; 
        10'b0111111110: data <= 14'h3ff0; 
        10'b0111111111: data <= 14'h000f; 
        10'b1000000000: data <= 14'h002b; 
        10'b1000000001: data <= 14'h004d; 
        10'b1000000010: data <= 14'h0036; 
        10'b1000000011: data <= 14'h004a; 
        10'b1000000100: data <= 14'h0030; 
        10'b1000000101: data <= 14'h001c; 
        10'b1000000110: data <= 14'h3fdf; 
        10'b1000000111: data <= 14'h3ff7; 
        10'b1000001000: data <= 14'h3fed; 
        10'b1000001001: data <= 14'h3fce; 
        10'b1000001010: data <= 14'h3ff4; 
        10'b1000001011: data <= 14'h3ff7; 
        10'b1000001100: data <= 14'h0004; 
        10'b1000001101: data <= 14'h3fe4; 
        10'b1000001110: data <= 14'h3ffc; 
        10'b1000001111: data <= 14'h3fe9; 
        10'b1000010000: data <= 14'h3fe0; 
        10'b1000010001: data <= 14'h3ff0; 
        10'b1000010010: data <= 14'h3ffd; 
        10'b1000010011: data <= 14'h0002; 
        10'b1000010100: data <= 14'h3ff6; 
        10'b1000010101: data <= 14'h3ffb; 
        10'b1000010110: data <= 14'h3ffc; 
        10'b1000010111: data <= 14'h3fea; 
        10'b1000011000: data <= 14'h3fe4; 
        10'b1000011001: data <= 14'h3ff5; 
        10'b1000011010: data <= 14'h0007; 
        10'b1000011011: data <= 14'h0014; 
        10'b1000011100: data <= 14'h0015; 
        10'b1000011101: data <= 14'h0034; 
        10'b1000011110: data <= 14'h001b; 
        10'b1000011111: data <= 14'h3ffc; 
        10'b1000100000: data <= 14'h000d; 
        10'b1000100001: data <= 14'h3fdd; 
        10'b1000100010: data <= 14'h3fd7; 
        10'b1000100011: data <= 14'h3ff0; 
        10'b1000100100: data <= 14'h3ff3; 
        10'b1000100101: data <= 14'h3fef; 
        10'b1000100110: data <= 14'h000d; 
        10'b1000100111: data <= 14'h0004; 
        10'b1000101000: data <= 14'h0011; 
        10'b1000101001: data <= 14'h0001; 
        10'b1000101010: data <= 14'h000b; 
        10'b1000101011: data <= 14'h3ff7; 
        10'b1000101100: data <= 14'h3fe8; 
        10'b1000101101: data <= 14'h3ff1; 
        10'b1000101110: data <= 14'h3ff4; 
        10'b1000101111: data <= 14'h0001; 
        10'b1000110000: data <= 14'h3ff4; 
        10'b1000110001: data <= 14'h3ffd; 
        10'b1000110010: data <= 14'h3ff5; 
        10'b1000110011: data <= 14'h3ff0; 
        10'b1000110100: data <= 14'h3fe0; 
        10'b1000110101: data <= 14'h3ffb; 
        10'b1000110110: data <= 14'h0005; 
        10'b1000110111: data <= 14'h002d; 
        10'b1000111000: data <= 14'h000d; 
        10'b1000111001: data <= 14'h3ffa; 
        10'b1000111010: data <= 14'h0000; 
        10'b1000111011: data <= 14'h3fda; 
        10'b1000111100: data <= 14'h0002; 
        10'b1000111101: data <= 14'h3fff; 
        10'b1000111110: data <= 14'h3fdc; 
        10'b1000111111: data <= 14'h3ff9; 
        10'b1001000000: data <= 14'h3fd6; 
        10'b1001000001: data <= 14'h3ff3; 
        10'b1001000010: data <= 14'h0007; 
        10'b1001000011: data <= 14'h0005; 
        10'b1001000100: data <= 14'h000d; 
        10'b1001000101: data <= 14'h0017; 
        10'b1001000110: data <= 14'h0017; 
        10'b1001000111: data <= 14'h3ffa; 
        10'b1001001000: data <= 14'h3ff1; 
        10'b1001001001: data <= 14'h3fec; 
        10'b1001001010: data <= 14'h3ffa; 
        10'b1001001011: data <= 14'h3ff5; 
        10'b1001001100: data <= 14'h0001; 
        10'b1001001101: data <= 14'h3ffa; 
        10'b1001001110: data <= 14'h0002; 
        10'b1001001111: data <= 14'h3fe7; 
        10'b1001010000: data <= 14'h3fdb; 
        10'b1001010001: data <= 14'h3ffc; 
        10'b1001010010: data <= 14'h0014; 
        10'b1001010011: data <= 14'h002a; 
        10'b1001010100: data <= 14'h0009; 
        10'b1001010101: data <= 14'h0012; 
        10'b1001010110: data <= 14'h3ffd; 
        10'b1001010111: data <= 14'h3fe4; 
        10'b1001011000: data <= 14'h3ff1; 
        10'b1001011001: data <= 14'h000a; 
        10'b1001011010: data <= 14'h3fff; 
        10'b1001011011: data <= 14'h3ffc; 
        10'b1001011100: data <= 14'h3fe0; 
        10'b1001011101: data <= 14'h3ff2; 
        10'b1001011110: data <= 14'h3ff7; 
        10'b1001011111: data <= 14'h3fff; 
        10'b1001100000: data <= 14'h3fff; 
        10'b1001100001: data <= 14'h0008; 
        10'b1001100010: data <= 14'h0007; 
        10'b1001100011: data <= 14'h3ff6; 
        10'b1001100100: data <= 14'h3ff4; 
        10'b1001100101: data <= 14'h3fff; 
        10'b1001100110: data <= 14'h3ffe; 
        10'b1001100111: data <= 14'h3ff8; 
        10'b1001101000: data <= 14'h3ffc; 
        10'b1001101001: data <= 14'h3ff2; 
        10'b1001101010: data <= 14'h3ff7; 
        10'b1001101011: data <= 14'h3ff0; 
        10'b1001101100: data <= 14'h3fe2; 
        10'b1001101101: data <= 14'h3fd4; 
        10'b1001101110: data <= 14'h0005; 
        10'b1001101111: data <= 14'h000c; 
        10'b1001110000: data <= 14'h3ffd; 
        10'b1001110001: data <= 14'h3ff2; 
        10'b1001110010: data <= 14'h0009; 
        10'b1001110011: data <= 14'h0003; 
        10'b1001110100: data <= 14'h0035; 
        10'b1001110101: data <= 14'h0037; 
        10'b1001110110: data <= 14'h0027; 
        10'b1001110111: data <= 14'h001f; 
        10'b1001111000: data <= 14'h3ffd; 
        10'b1001111001: data <= 14'h3ffd; 
        10'b1001111010: data <= 14'h000d; 
        10'b1001111011: data <= 14'h3ff0; 
        10'b1001111100: data <= 14'h3fee; 
        10'b1001111101: data <= 14'h0008; 
        10'b1001111110: data <= 14'h3ffd; 
        10'b1001111111: data <= 14'h3ff5; 
        10'b1010000000: data <= 14'h3ffd; 
        10'b1010000001: data <= 14'h3ffd; 
        10'b1010000010: data <= 14'h3ffd; 
        10'b1010000011: data <= 14'h3ff5; 
        10'b1010000100: data <= 14'h3ff5; 
        10'b1010000101: data <= 14'h3fff; 
        10'b1010000110: data <= 14'h3ffb; 
        10'b1010000111: data <= 14'h3ff2; 
        10'b1010001000: data <= 14'h3fe1; 
        10'b1010001001: data <= 14'h3fb6; 
        10'b1010001010: data <= 14'h3fc6; 
        10'b1010001011: data <= 14'h3fe3; 
        10'b1010001100: data <= 14'h000a; 
        10'b1010001101: data <= 14'h000a; 
        10'b1010001110: data <= 14'h0015; 
        10'b1010001111: data <= 14'h001c; 
        10'b1010010000: data <= 14'h003f; 
        10'b1010010001: data <= 14'h005a; 
        10'b1010010010: data <= 14'h004d; 
        10'b1010010011: data <= 14'h003d; 
        10'b1010010100: data <= 14'h0031; 
        10'b1010010101: data <= 14'h0023; 
        10'b1010010110: data <= 14'h001c; 
        10'b1010010111: data <= 14'h0024; 
        10'b1010011000: data <= 14'h001b; 
        10'b1010011001: data <= 14'h0006; 
        10'b1010011010: data <= 14'h3ffd; 
        10'b1010011011: data <= 14'h3ff8; 
        10'b1010011100: data <= 14'h3ff0; 
        10'b1010011101: data <= 14'h3ffe; 
        10'b1010011110: data <= 14'h3ff2; 
        10'b1010011111: data <= 14'h3ffd; 
        10'b1010100000: data <= 14'h3ffe; 
        10'b1010100001: data <= 14'h3ffd; 
        10'b1010100010: data <= 14'h0003; 
        10'b1010100011: data <= 14'h3ff3; 
        10'b1010100100: data <= 14'h3ff3; 
        10'b1010100101: data <= 14'h3fcf; 
        10'b1010100110: data <= 14'h3fbc; 
        10'b1010100111: data <= 14'h3fc7; 
        10'b1010101000: data <= 14'h3ffc; 
        10'b1010101001: data <= 14'h000d; 
        10'b1010101010: data <= 14'h3ffb; 
        10'b1010101011: data <= 14'h0018; 
        10'b1010101100: data <= 14'h0012; 
        10'b1010101101: data <= 14'h000c; 
        10'b1010101110: data <= 14'h001e; 
        10'b1010101111: data <= 14'h0040; 
        10'b1010110000: data <= 14'h0044; 
        10'b1010110001: data <= 14'h002e; 
        10'b1010110010: data <= 14'h0040; 
        10'b1010110011: data <= 14'h003c; 
        10'b1010110100: data <= 14'h0014; 
        10'b1010110101: data <= 14'h0001; 
        10'b1010110110: data <= 14'h3ff2; 
        10'b1010110111: data <= 14'h0001; 
        10'b1010111000: data <= 14'h3ffa; 
        10'b1010111001: data <= 14'h3ff7; 
        10'b1010111010: data <= 14'h0002; 
        10'b1010111011: data <= 14'h3ffc; 
        10'b1010111100: data <= 14'h0003; 
        10'b1010111101: data <= 14'h3ffe; 
        10'b1010111110: data <= 14'h0001; 
        10'b1010111111: data <= 14'h3ff3; 
        10'b1011000000: data <= 14'h3ff6; 
        10'b1011000001: data <= 14'h3fee; 
        10'b1011000010: data <= 14'h3fe6; 
        10'b1011000011: data <= 14'h3fe0; 
        10'b1011000100: data <= 14'h3fdc; 
        10'b1011000101: data <= 14'h3fdc; 
        10'b1011000110: data <= 14'h3ff3; 
        10'b1011000111: data <= 14'h3fe7; 
        10'b1011001000: data <= 14'h3ff1; 
        10'b1011001001: data <= 14'h3ff1; 
        10'b1011001010: data <= 14'h3ffe; 
        10'b1011001011: data <= 14'h0017; 
        10'b1011001100: data <= 14'h0010; 
        10'b1011001101: data <= 14'h0014; 
        10'b1011001110: data <= 14'h0017; 
        10'b1011001111: data <= 14'h0004; 
        10'b1011010000: data <= 14'h3ffb; 
        10'b1011010001: data <= 14'h3fff; 
        10'b1011010010: data <= 14'h3ff1; 
        10'b1011010011: data <= 14'h3ff1; 
        10'b1011010100: data <= 14'h3fff; 
        10'b1011010101: data <= 14'h3ffc; 
        10'b1011010110: data <= 14'h3ff6; 
        10'b1011010111: data <= 14'h3ffc; 
        10'b1011011000: data <= 14'h3ffe; 
        10'b1011011001: data <= 14'h0000; 
        10'b1011011010: data <= 14'h3ff9; 
        10'b1011011011: data <= 14'h3ff6; 
        10'b1011011100: data <= 14'h3ff1; 
        10'b1011011101: data <= 14'h3ff3; 
        10'b1011011110: data <= 14'h3fed; 
        10'b1011011111: data <= 14'h3ffb; 
        10'b1011100000: data <= 14'h3fee; 
        10'b1011100001: data <= 14'h3ff1; 
        10'b1011100010: data <= 14'h3fee; 
        10'b1011100011: data <= 14'h3ff6; 
        10'b1011100100: data <= 14'h3ff5; 
        10'b1011100101: data <= 14'h3ff6; 
        10'b1011100110: data <= 14'h3ff2; 
        10'b1011100111: data <= 14'h3ff6; 
        10'b1011101000: data <= 14'h3ff3; 
        10'b1011101001: data <= 14'h3fef; 
        10'b1011101010: data <= 14'h3fed; 
        10'b1011101011: data <= 14'h3ff4; 
        10'b1011101100: data <= 14'h3ff8; 
        10'b1011101101: data <= 14'h3ffd; 
        10'b1011101110: data <= 14'h3ff9; 
        10'b1011101111: data <= 14'h0003; 
        10'b1011110000: data <= 14'h0003; 
        10'b1011110001: data <= 14'h3ff2; 
        10'b1011110010: data <= 14'h3ffc; 
        10'b1011110011: data <= 14'h3ffa; 
        10'b1011110100: data <= 14'h3ffd; 
        10'b1011110101: data <= 14'h3ff5; 
        10'b1011110110: data <= 14'h3ff9; 
        10'b1011110111: data <= 14'h3ffc; 
        10'b1011111000: data <= 14'h3ffc; 
        10'b1011111001: data <= 14'h3ff2; 
        10'b1011111010: data <= 14'h3fff; 
        10'b1011111011: data <= 14'h3ff6; 
        10'b1011111100: data <= 14'h0002; 
        10'b1011111101: data <= 14'h3ff9; 
        10'b1011111110: data <= 14'h3ff4; 
        10'b1011111111: data <= 14'h3fff; 
        10'b1100000000: data <= 14'h3ff6; 
        10'b1100000001: data <= 14'h3ff4; 
        10'b1100000010: data <= 14'h3ff8; 
        10'b1100000011: data <= 14'h3ffd; 
        10'b1100000100: data <= 14'h3ffb; 
        10'b1100000101: data <= 14'h0000; 
        10'b1100000110: data <= 14'h0002; 
        10'b1100000111: data <= 14'h0003; 
        10'b1100001000: data <= 14'h3ffe; 
        10'b1100001001: data <= 14'h3ffc; 
        10'b1100001010: data <= 14'h3ffd; 
        10'b1100001011: data <= 14'h3ff5; 
        10'b1100001100: data <= 14'h3ffb; 
        10'b1100001101: data <= 14'h0002; 
        10'b1100001110: data <= 14'h3ff3; 
        10'b1100001111: data <= 14'h3ffb; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 9) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 15'h7ff2; 
        10'b0000000001: data <= 15'h7ff5; 
        10'b0000000010: data <= 15'h7ff2; 
        10'b0000000011: data <= 15'h7ff9; 
        10'b0000000100: data <= 15'h7ff8; 
        10'b0000000101: data <= 15'h0003; 
        10'b0000000110: data <= 15'h7fe3; 
        10'b0000000111: data <= 15'h7ffa; 
        10'b0000001000: data <= 15'h7fec; 
        10'b0000001001: data <= 15'h7fef; 
        10'b0000001010: data <= 15'h7fe8; 
        10'b0000001011: data <= 15'h0002; 
        10'b0000001100: data <= 15'h7ff7; 
        10'b0000001101: data <= 15'h7ffe; 
        10'b0000001110: data <= 15'h7fe8; 
        10'b0000001111: data <= 15'h7fff; 
        10'b0000010000: data <= 15'h7ff8; 
        10'b0000010001: data <= 15'h7fe6; 
        10'b0000010010: data <= 15'h0003; 
        10'b0000010011: data <= 15'h7ff4; 
        10'b0000010100: data <= 15'h7ff2; 
        10'b0000010101: data <= 15'h7ff1; 
        10'b0000010110: data <= 15'h7ff3; 
        10'b0000010111: data <= 15'h0005; 
        10'b0000011000: data <= 15'h0000; 
        10'b0000011001: data <= 15'h7fef; 
        10'b0000011010: data <= 15'h7feb; 
        10'b0000011011: data <= 15'h7ff3; 
        10'b0000011100: data <= 15'h7ff2; 
        10'b0000011101: data <= 15'h7fe3; 
        10'b0000011110: data <= 15'h0005; 
        10'b0000011111: data <= 15'h0000; 
        10'b0000100000: data <= 15'h7fe5; 
        10'b0000100001: data <= 15'h7fe6; 
        10'b0000100010: data <= 15'h7fe4; 
        10'b0000100011: data <= 15'h7fe6; 
        10'b0000100100: data <= 15'h0004; 
        10'b0000100101: data <= 15'h7ff5; 
        10'b0000100110: data <= 15'h7ff4; 
        10'b0000100111: data <= 15'h7fe3; 
        10'b0000101000: data <= 15'h0003; 
        10'b0000101001: data <= 15'h7ffb; 
        10'b0000101010: data <= 15'h7fec; 
        10'b0000101011: data <= 15'h7ff1; 
        10'b0000101100: data <= 15'h7ffc; 
        10'b0000101101: data <= 15'h7ff7; 
        10'b0000101110: data <= 15'h7fe9; 
        10'b0000101111: data <= 15'h7ff7; 
        10'b0000110000: data <= 15'h0003; 
        10'b0000110001: data <= 15'h7fe5; 
        10'b0000110010: data <= 15'h7ffb; 
        10'b0000110011: data <= 15'h7fea; 
        10'b0000110100: data <= 15'h7ffe; 
        10'b0000110101: data <= 15'h0006; 
        10'b0000110110: data <= 15'h7fec; 
        10'b0000110111: data <= 15'h7fea; 
        10'b0000111000: data <= 15'h7fe8; 
        10'b0000111001: data <= 15'h0000; 
        10'b0000111010: data <= 15'h7ff6; 
        10'b0000111011: data <= 15'h7ff4; 
        10'b0000111100: data <= 15'h7fe9; 
        10'b0000111101: data <= 15'h7fe3; 
        10'b0000111110: data <= 15'h7ff6; 
        10'b0000111111: data <= 15'h7fe3; 
        10'b0001000000: data <= 15'h0005; 
        10'b0001000001: data <= 15'h7fe2; 
        10'b0001000010: data <= 15'h7fe4; 
        10'b0001000011: data <= 15'h7ffa; 
        10'b0001000100: data <= 15'h7ff6; 
        10'b0001000101: data <= 15'h7fe2; 
        10'b0001000110: data <= 15'h7ffa; 
        10'b0001000111: data <= 15'h7ff8; 
        10'b0001001000: data <= 15'h7fe0; 
        10'b0001001001: data <= 15'h7fed; 
        10'b0001001010: data <= 15'h7fed; 
        10'b0001001011: data <= 15'h7ffc; 
        10'b0001001100: data <= 15'h7fff; 
        10'b0001001101: data <= 15'h7ffe; 
        10'b0001001110: data <= 15'h7ff9; 
        10'b0001001111: data <= 15'h7ff3; 
        10'b0001010000: data <= 15'h0003; 
        10'b0001010001: data <= 15'h7fec; 
        10'b0001010010: data <= 15'h7ffb; 
        10'b0001010011: data <= 15'h0004; 
        10'b0001010100: data <= 15'h7fea; 
        10'b0001010101: data <= 15'h7ff3; 
        10'b0001010110: data <= 15'h7ff4; 
        10'b0001010111: data <= 15'h7fe7; 
        10'b0001011000: data <= 15'h0005; 
        10'b0001011001: data <= 15'h7fe8; 
        10'b0001011010: data <= 15'h7fe4; 
        10'b0001011011: data <= 15'h7fef; 
        10'b0001011100: data <= 15'h7fe3; 
        10'b0001011101: data <= 15'h7ff6; 
        10'b0001011110: data <= 15'h7fea; 
        10'b0001011111: data <= 15'h7fd8; 
        10'b0001100000: data <= 15'h7fd3; 
        10'b0001100001: data <= 15'h7fca; 
        10'b0001100010: data <= 15'h7fd3; 
        10'b0001100011: data <= 15'h7fe5; 
        10'b0001100100: data <= 15'h7fd3; 
        10'b0001100101: data <= 15'h7fdd; 
        10'b0001100110: data <= 15'h7fe8; 
        10'b0001100111: data <= 15'h7ff1; 
        10'b0001101000: data <= 15'h7fde; 
        10'b0001101001: data <= 15'h0002; 
        10'b0001101010: data <= 15'h7fee; 
        10'b0001101011: data <= 15'h7ffe; 
        10'b0001101100: data <= 15'h7fed; 
        10'b0001101101: data <= 15'h7ffa; 
        10'b0001101110: data <= 15'h7ff7; 
        10'b0001101111: data <= 15'h7fe5; 
        10'b0001110000: data <= 15'h7ff4; 
        10'b0001110001: data <= 15'h7ffd; 
        10'b0001110010: data <= 15'h7fef; 
        10'b0001110011: data <= 15'h7fe5; 
        10'b0001110100: data <= 15'h7fff; 
        10'b0001110101: data <= 15'h7ffe; 
        10'b0001110110: data <= 15'h7ff4; 
        10'b0001110111: data <= 15'h7fe8; 
        10'b0001111000: data <= 15'h7fe8; 
        10'b0001111001: data <= 15'h7ff2; 
        10'b0001111010: data <= 15'h7ff3; 
        10'b0001111011: data <= 15'h7ff9; 
        10'b0001111100: data <= 15'h0027; 
        10'b0001111101: data <= 15'h0019; 
        10'b0001111110: data <= 15'h0055; 
        10'b0001111111: data <= 15'h0040; 
        10'b0010000000: data <= 15'h001d; 
        10'b0010000001: data <= 15'h0010; 
        10'b0010000010: data <= 15'h0018; 
        10'b0010000011: data <= 15'h7feb; 
        10'b0010000100: data <= 15'h7fe6; 
        10'b0010000101: data <= 15'h7ff2; 
        10'b0010000110: data <= 15'h7fd9; 
        10'b0010000111: data <= 15'h7fe4; 
        10'b0010001000: data <= 15'h7fff; 
        10'b0010001001: data <= 15'h0002; 
        10'b0010001010: data <= 15'h7ff1; 
        10'b0010001011: data <= 15'h7ff4; 
        10'b0010001100: data <= 15'h7ff5; 
        10'b0010001101: data <= 15'h7ffb; 
        10'b0010001110: data <= 15'h7ffd; 
        10'b0010001111: data <= 15'h7fff; 
        10'b0010010000: data <= 15'h7fe9; 
        10'b0010010001: data <= 15'h7ff2; 
        10'b0010010010: data <= 15'h7fec; 
        10'b0010010011: data <= 15'h7fca; 
        10'b0010010100: data <= 15'h7fea; 
        10'b0010010101: data <= 15'h0013; 
        10'b0010010110: data <= 15'h7fd4; 
        10'b0010010111: data <= 15'h003b; 
        10'b0010011000: data <= 15'h006f; 
        10'b0010011001: data <= 15'h005d; 
        10'b0010011010: data <= 15'h0060; 
        10'b0010011011: data <= 15'h002e; 
        10'b0010011100: data <= 15'h0026; 
        10'b0010011101: data <= 15'h0059; 
        10'b0010011110: data <= 15'h0004; 
        10'b0010011111: data <= 15'h7ffc; 
        10'b0010100000: data <= 15'h0020; 
        10'b0010100001: data <= 15'h0010; 
        10'b0010100010: data <= 15'h7fca; 
        10'b0010100011: data <= 15'h7fd3; 
        10'b0010100100: data <= 15'h7fe1; 
        10'b0010100101: data <= 15'h0018; 
        10'b0010100110: data <= 15'h7ff6; 
        10'b0010100111: data <= 15'h0004; 
        10'b0010101000: data <= 15'h7fea; 
        10'b0010101001: data <= 15'h7fe8; 
        10'b0010101010: data <= 15'h7fe3; 
        10'b0010101011: data <= 15'h7fe4; 
        10'b0010101100: data <= 15'h7fe0; 
        10'b0010101101: data <= 15'h7fe0; 
        10'b0010101110: data <= 15'h7fcd; 
        10'b0010101111: data <= 15'h7fcd; 
        10'b0010110000: data <= 15'h0004; 
        10'b0010110001: data <= 15'h000f; 
        10'b0010110010: data <= 15'h7ffc; 
        10'b0010110011: data <= 15'h001d; 
        10'b0010110100: data <= 15'h002d; 
        10'b0010110101: data <= 15'h0024; 
        10'b0010110110: data <= 15'h0033; 
        10'b0010110111: data <= 15'h0060; 
        10'b0010111000: data <= 15'h002e; 
        10'b0010111001: data <= 15'h0037; 
        10'b0010111010: data <= 15'h000c; 
        10'b0010111011: data <= 15'h003e; 
        10'b0010111100: data <= 15'h0018; 
        10'b0010111101: data <= 15'h001d; 
        10'b0010111110: data <= 15'h0024; 
        10'b0010111111: data <= 15'h0022; 
        10'b0011000000: data <= 15'h001d; 
        10'b0011000001: data <= 15'h000c; 
        10'b0011000010: data <= 15'h7ff4; 
        10'b0011000011: data <= 15'h7ffd; 
        10'b0011000100: data <= 15'h0004; 
        10'b0011000101: data <= 15'h7fea; 
        10'b0011000110: data <= 15'h7fe6; 
        10'b0011000111: data <= 15'h7fec; 
        10'b0011001000: data <= 15'h7fde; 
        10'b0011001001: data <= 15'h7ff4; 
        10'b0011001010: data <= 15'h7fdd; 
        10'b0011001011: data <= 15'h7ffe; 
        10'b0011001100: data <= 15'h0022; 
        10'b0011001101: data <= 15'h000e; 
        10'b0011001110: data <= 15'h0011; 
        10'b0011001111: data <= 15'h7ff5; 
        10'b0011010000: data <= 15'h7fd4; 
        10'b0011010001: data <= 15'h7fdf; 
        10'b0011010010: data <= 15'h7fd0; 
        10'b0011010011: data <= 15'h001d; 
        10'b0011010100: data <= 15'h0024; 
        10'b0011010101: data <= 15'h7ffe; 
        10'b0011010110: data <= 15'h0019; 
        10'b0011010111: data <= 15'h7fe5; 
        10'b0011011000: data <= 15'h0025; 
        10'b0011011001: data <= 15'h003a; 
        10'b0011011010: data <= 15'h000a; 
        10'b0011011011: data <= 15'h0078; 
        10'b0011011100: data <= 15'h004a; 
        10'b0011011101: data <= 15'h7ffd; 
        10'b0011011110: data <= 15'h0002; 
        10'b0011011111: data <= 15'h7ffb; 
        10'b0011100000: data <= 15'h7ffb; 
        10'b0011100001: data <= 15'h0002; 
        10'b0011100010: data <= 15'h7ffa; 
        10'b0011100011: data <= 15'h7fe8; 
        10'b0011100100: data <= 15'h7ffa; 
        10'b0011100101: data <= 15'h7ff5; 
        10'b0011100110: data <= 15'h0032; 
        10'b0011100111: data <= 15'h001f; 
        10'b0011101000: data <= 15'h000b; 
        10'b0011101001: data <= 15'h0056; 
        10'b0011101010: data <= 15'h0005; 
        10'b0011101011: data <= 15'h0003; 
        10'b0011101100: data <= 15'h003a; 
        10'b0011101101: data <= 15'h004b; 
        10'b0011101110: data <= 15'h7fc5; 
        10'b0011101111: data <= 15'h7fce; 
        10'b0011110000: data <= 15'h0029; 
        10'b0011110001: data <= 15'h7fe3; 
        10'b0011110010: data <= 15'h000e; 
        10'b0011110011: data <= 15'h0027; 
        10'b0011110100: data <= 15'h001a; 
        10'b0011110101: data <= 15'h0050; 
        10'b0011110110: data <= 15'h0035; 
        10'b0011110111: data <= 15'h005b; 
        10'b0011111000: data <= 15'h0053; 
        10'b0011111001: data <= 15'h7ff6; 
        10'b0011111010: data <= 15'h7ff9; 
        10'b0011111011: data <= 15'h0008; 
        10'b0011111100: data <= 15'h0000; 
        10'b0011111101: data <= 15'h0002; 
        10'b0011111110: data <= 15'h7ff3; 
        10'b0011111111: data <= 15'h7ff0; 
        10'b0100000000: data <= 15'h7ff7; 
        10'b0100000001: data <= 15'h0032; 
        10'b0100000010: data <= 15'h0025; 
        10'b0100000011: data <= 15'h004d; 
        10'b0100000100: data <= 15'h0067; 
        10'b0100000101: data <= 15'h0057; 
        10'b0100000110: data <= 15'h0037; 
        10'b0100000111: data <= 15'h0061; 
        10'b0100001000: data <= 15'h001a; 
        10'b0100001001: data <= 15'h001c; 
        10'b0100001010: data <= 15'h7f8f; 
        10'b0100001011: data <= 15'h7f62; 
        10'b0100001100: data <= 15'h7fc9; 
        10'b0100001101: data <= 15'h0008; 
        10'b0100001110: data <= 15'h0011; 
        10'b0100001111: data <= 15'h001f; 
        10'b0100010000: data <= 15'h0028; 
        10'b0100010001: data <= 15'h0023; 
        10'b0100010010: data <= 15'h0053; 
        10'b0100010011: data <= 15'h0056; 
        10'b0100010100: data <= 15'h7ff2; 
        10'b0100010101: data <= 15'h7ff4; 
        10'b0100010110: data <= 15'h0013; 
        10'b0100010111: data <= 15'h7fe6; 
        10'b0100011000: data <= 15'h7feb; 
        10'b0100011001: data <= 15'h0001; 
        10'b0100011010: data <= 15'h7fea; 
        10'b0100011011: data <= 15'h0002; 
        10'b0100011100: data <= 15'h0013; 
        10'b0100011101: data <= 15'h003e; 
        10'b0100011110: data <= 15'h003e; 
        10'b0100011111: data <= 15'h0071; 
        10'b0100100000: data <= 15'h0054; 
        10'b0100100001: data <= 15'h0062; 
        10'b0100100010: data <= 15'h008f; 
        10'b0100100011: data <= 15'h0045; 
        10'b0100100100: data <= 15'h0048; 
        10'b0100100101: data <= 15'h003a; 
        10'b0100100110: data <= 15'h7fed; 
        10'b0100100111: data <= 15'h7f6a; 
        10'b0100101000: data <= 15'h7f85; 
        10'b0100101001: data <= 15'h7fda; 
        10'b0100101010: data <= 15'h002b; 
        10'b0100101011: data <= 15'h002b; 
        10'b0100101100: data <= 15'h002c; 
        10'b0100101101: data <= 15'h0066; 
        10'b0100101110: data <= 15'h0070; 
        10'b0100101111: data <= 15'h005c; 
        10'b0100110000: data <= 15'h0001; 
        10'b0100110001: data <= 15'h7ff9; 
        10'b0100110010: data <= 15'h7ff4; 
        10'b0100110011: data <= 15'h7fec; 
        10'b0100110100: data <= 15'h7fea; 
        10'b0100110101: data <= 15'h0005; 
        10'b0100110110: data <= 15'h7ffe; 
        10'b0100110111: data <= 15'h7fdd; 
        10'b0100111000: data <= 15'h001e; 
        10'b0100111001: data <= 15'h0044; 
        10'b0100111010: data <= 15'h0082; 
        10'b0100111011: data <= 15'h00a9; 
        10'b0100111100: data <= 15'h0085; 
        10'b0100111101: data <= 15'h00a8; 
        10'b0100111110: data <= 15'h0073; 
        10'b0100111111: data <= 15'h0036; 
        10'b0101000000: data <= 15'h0046; 
        10'b0101000001: data <= 15'h00a7; 
        10'b0101000010: data <= 15'h00cb; 
        10'b0101000011: data <= 15'h7fe7; 
        10'b0101000100: data <= 15'h7f87; 
        10'b0101000101: data <= 15'h7fd6; 
        10'b0101000110: data <= 15'h7fd8; 
        10'b0101000111: data <= 15'h0011; 
        10'b0101001000: data <= 15'h005c; 
        10'b0101001001: data <= 15'h006e; 
        10'b0101001010: data <= 15'h0092; 
        10'b0101001011: data <= 15'h008a; 
        10'b0101001100: data <= 15'h0060; 
        10'b0101001101: data <= 15'h0010; 
        10'b0101001110: data <= 15'h0008; 
        10'b0101001111: data <= 15'h7ff8; 
        10'b0101010000: data <= 15'h7fed; 
        10'b0101010001: data <= 15'h7ffa; 
        10'b0101010010: data <= 15'h7ff0; 
        10'b0101010011: data <= 15'h7ff8; 
        10'b0101010100: data <= 15'h7ffa; 
        10'b0101010101: data <= 15'h0052; 
        10'b0101010110: data <= 15'h0044; 
        10'b0101010111: data <= 15'h0067; 
        10'b0101011000: data <= 15'h0062; 
        10'b0101011001: data <= 15'h007b; 
        10'b0101011010: data <= 15'h0015; 
        10'b0101011011: data <= 15'h001d; 
        10'b0101011100: data <= 15'h0010; 
        10'b0101011101: data <= 15'h00ca; 
        10'b0101011110: data <= 15'h00cb; 
        10'b0101011111: data <= 15'h002d; 
        10'b0101100000: data <= 15'h0008; 
        10'b0101100001: data <= 15'h7fee; 
        10'b0101100010: data <= 15'h7ff1; 
        10'b0101100011: data <= 15'h0033; 
        10'b0101100100: data <= 15'h0056; 
        10'b0101100101: data <= 15'h0094; 
        10'b0101100110: data <= 15'h00ad; 
        10'b0101100111: data <= 15'h0090; 
        10'b0101101000: data <= 15'h005a; 
        10'b0101101001: data <= 15'h0024; 
        10'b0101101010: data <= 15'h0012; 
        10'b0101101011: data <= 15'h7fe7; 
        10'b0101101100: data <= 15'h7fe4; 
        10'b0101101101: data <= 15'h7ff6; 
        10'b0101101110: data <= 15'h0006; 
        10'b0101101111: data <= 15'h7fe8; 
        10'b0101110000: data <= 15'h7fee; 
        10'b0101110001: data <= 15'h0000; 
        10'b0101110010: data <= 15'h7ff3; 
        10'b0101110011: data <= 15'h7ff4; 
        10'b0101110100: data <= 15'h000b; 
        10'b0101110101: data <= 15'h7ff1; 
        10'b0101110110: data <= 15'h7fd4; 
        10'b0101110111: data <= 15'h0011; 
        10'b0101111000: data <= 15'h004a; 
        10'b0101111001: data <= 15'h00bd; 
        10'b0101111010: data <= 15'h0039; 
        10'b0101111011: data <= 15'h008b; 
        10'b0101111100: data <= 15'h0037; 
        10'b0101111101: data <= 15'h7fdd; 
        10'b0101111110: data <= 15'h0003; 
        10'b0101111111: data <= 15'h0005; 
        10'b0110000000: data <= 15'h003e; 
        10'b0110000001: data <= 15'h0038; 
        10'b0110000010: data <= 15'h0020; 
        10'b0110000011: data <= 15'h002d; 
        10'b0110000100: data <= 15'h0018; 
        10'b0110000101: data <= 15'h0005; 
        10'b0110000110: data <= 15'h0005; 
        10'b0110000111: data <= 15'h7ffb; 
        10'b0110001000: data <= 15'h7fef; 
        10'b0110001001: data <= 15'h7fe3; 
        10'b0110001010: data <= 15'h7ffc; 
        10'b0110001011: data <= 15'h7ff4; 
        10'b0110001100: data <= 15'h7fe7; 
        10'b0110001101: data <= 15'h7fc9; 
        10'b0110001110: data <= 15'h7f9e; 
        10'b0110001111: data <= 15'h7f82; 
        10'b0110010000: data <= 15'h7f6c; 
        10'b0110010001: data <= 15'h7f89; 
        10'b0110010010: data <= 15'h7fef; 
        10'b0110010011: data <= 15'h004c; 
        10'b0110010100: data <= 15'h0049; 
        10'b0110010101: data <= 15'h009a; 
        10'b0110010110: data <= 15'h007b; 
        10'b0110010111: data <= 15'h0054; 
        10'b0110011000: data <= 15'h7ff6; 
        10'b0110011001: data <= 15'h000a; 
        10'b0110011010: data <= 15'h7fea; 
        10'b0110011011: data <= 15'h7fce; 
        10'b0110011100: data <= 15'h7fae; 
        10'b0110011101: data <= 15'h7fb7; 
        10'b0110011110: data <= 15'h7fc1; 
        10'b0110011111: data <= 15'h7fb5; 
        10'b0110100000: data <= 15'h7fde; 
        10'b0110100001: data <= 15'h7ffb; 
        10'b0110100010: data <= 15'h7fe2; 
        10'b0110100011: data <= 15'h0001; 
        10'b0110100100: data <= 15'h0002; 
        10'b0110100101: data <= 15'h7fee; 
        10'b0110100110: data <= 15'h7feb; 
        10'b0110100111: data <= 15'h7ff7; 
        10'b0110101000: data <= 15'h7fe4; 
        10'b0110101001: data <= 15'h7fc9; 
        10'b0110101010: data <= 15'h7f86; 
        10'b0110101011: data <= 15'h7f6a; 
        10'b0110101100: data <= 15'h7f78; 
        10'b0110101101: data <= 15'h7fdf; 
        10'b0110101110: data <= 15'h0005; 
        10'b0110101111: data <= 15'h0003; 
        10'b0110110000: data <= 15'h0069; 
        10'b0110110001: data <= 15'h007d; 
        10'b0110110010: data <= 15'h006d; 
        10'b0110110011: data <= 15'h003f; 
        10'b0110110100: data <= 15'h7fe0; 
        10'b0110110101: data <= 15'h7fe5; 
        10'b0110110110: data <= 15'h7fed; 
        10'b0110110111: data <= 15'h7f92; 
        10'b0110111000: data <= 15'h7f76; 
        10'b0110111001: data <= 15'h7f96; 
        10'b0110111010: data <= 15'h7fbd; 
        10'b0110111011: data <= 15'h7fc0; 
        10'b0110111100: data <= 15'h7fd0; 
        10'b0110111101: data <= 15'h7ff8; 
        10'b0110111110: data <= 15'h7fdf; 
        10'b0110111111: data <= 15'h0003; 
        10'b0111000000: data <= 15'h7ff1; 
        10'b0111000001: data <= 15'h7fe5; 
        10'b0111000010: data <= 15'h7fed; 
        10'b0111000011: data <= 15'h7ff6; 
        10'b0111000100: data <= 15'h7fd4; 
        10'b0111000101: data <= 15'h7fb1; 
        10'b0111000110: data <= 15'h7f81; 
        10'b0111000111: data <= 15'h7fb5; 
        10'b0111001000: data <= 15'h0032; 
        10'b0111001001: data <= 15'h0038; 
        10'b0111001010: data <= 15'h0017; 
        10'b0111001011: data <= 15'h0033; 
        10'b0111001100: data <= 15'h0066; 
        10'b0111001101: data <= 15'h0059; 
        10'b0111001110: data <= 15'h0020; 
        10'b0111001111: data <= 15'h0035; 
        10'b0111010000: data <= 15'h0012; 
        10'b0111010001: data <= 15'h7fd6; 
        10'b0111010010: data <= 15'h7fa7; 
        10'b0111010011: data <= 15'h7f81; 
        10'b0111010100: data <= 15'h7f81; 
        10'b0111010101: data <= 15'h7f7f; 
        10'b0111010110: data <= 15'h7f98; 
        10'b0111010111: data <= 15'h7fde; 
        10'b0111011000: data <= 15'h7fd3; 
        10'b0111011001: data <= 15'h7ff0; 
        10'b0111011010: data <= 15'h7ff0; 
        10'b0111011011: data <= 15'h7fe4; 
        10'b0111011100: data <= 15'h0006; 
        10'b0111011101: data <= 15'h0004; 
        10'b0111011110: data <= 15'h7fea; 
        10'b0111011111: data <= 15'h7fe5; 
        10'b0111100000: data <= 15'h7fe3; 
        10'b0111100001: data <= 15'h7fae; 
        10'b0111100010: data <= 15'h7f90; 
        10'b0111100011: data <= 15'h0014; 
        10'b0111100100: data <= 15'h0068; 
        10'b0111100101: data <= 15'h0081; 
        10'b0111100110: data <= 15'h0029; 
        10'b0111100111: data <= 15'h0062; 
        10'b0111101000: data <= 15'h009f; 
        10'b0111101001: data <= 15'h0060; 
        10'b0111101010: data <= 15'h0008; 
        10'b0111101011: data <= 15'h7fe6; 
        10'b0111101100: data <= 15'h000c; 
        10'b0111101101: data <= 15'h7fcf; 
        10'b0111101110: data <= 15'h7f7d; 
        10'b0111101111: data <= 15'h7fc2; 
        10'b0111110000: data <= 15'h7fc2; 
        10'b0111110001: data <= 15'h7fa9; 
        10'b0111110010: data <= 15'h7fc0; 
        10'b0111110011: data <= 15'h7fd7; 
        10'b0111110100: data <= 15'h7fe9; 
        10'b0111110101: data <= 15'h7fdf; 
        10'b0111110110: data <= 15'h7ffb; 
        10'b0111110111: data <= 15'h7fef; 
        10'b0111111000: data <= 15'h7fec; 
        10'b0111111001: data <= 15'h0001; 
        10'b0111111010: data <= 15'h7fe4; 
        10'b0111111011: data <= 15'h7fdc; 
        10'b0111111100: data <= 15'h7fce; 
        10'b0111111101: data <= 15'h7fcd; 
        10'b0111111110: data <= 15'h7fe0; 
        10'b0111111111: data <= 15'h001f; 
        10'b1000000000: data <= 15'h0056; 
        10'b1000000001: data <= 15'h009a; 
        10'b1000000010: data <= 15'h006c; 
        10'b1000000011: data <= 15'h0093; 
        10'b1000000100: data <= 15'h0060; 
        10'b1000000101: data <= 15'h0037; 
        10'b1000000110: data <= 15'h7fbd; 
        10'b1000000111: data <= 15'h7fef; 
        10'b1000001000: data <= 15'h7fda; 
        10'b1000001001: data <= 15'h7f9c; 
        10'b1000001010: data <= 15'h7fe8; 
        10'b1000001011: data <= 15'h7fed; 
        10'b1000001100: data <= 15'h0007; 
        10'b1000001101: data <= 15'h7fc9; 
        10'b1000001110: data <= 15'h7ff8; 
        10'b1000001111: data <= 15'h7fd1; 
        10'b1000010000: data <= 15'h7fc0; 
        10'b1000010001: data <= 15'h7fdf; 
        10'b1000010010: data <= 15'h7ffb; 
        10'b1000010011: data <= 15'h0004; 
        10'b1000010100: data <= 15'h7fed; 
        10'b1000010101: data <= 15'h7ff6; 
        10'b1000010110: data <= 15'h7ff9; 
        10'b1000010111: data <= 15'h7fd5; 
        10'b1000011000: data <= 15'h7fc9; 
        10'b1000011001: data <= 15'h7fea; 
        10'b1000011010: data <= 15'h000f; 
        10'b1000011011: data <= 15'h0029; 
        10'b1000011100: data <= 15'h002a; 
        10'b1000011101: data <= 15'h0069; 
        10'b1000011110: data <= 15'h0036; 
        10'b1000011111: data <= 15'h7ff9; 
        10'b1000100000: data <= 15'h001a; 
        10'b1000100001: data <= 15'h7fba; 
        10'b1000100010: data <= 15'h7fae; 
        10'b1000100011: data <= 15'h7fe1; 
        10'b1000100100: data <= 15'h7fe6; 
        10'b1000100101: data <= 15'h7fde; 
        10'b1000100110: data <= 15'h001a; 
        10'b1000100111: data <= 15'h0007; 
        10'b1000101000: data <= 15'h0021; 
        10'b1000101001: data <= 15'h0003; 
        10'b1000101010: data <= 15'h0016; 
        10'b1000101011: data <= 15'h7fee; 
        10'b1000101100: data <= 15'h7fcf; 
        10'b1000101101: data <= 15'h7fe3; 
        10'b1000101110: data <= 15'h7fe7; 
        10'b1000101111: data <= 15'h0003; 
        10'b1000110000: data <= 15'h7fe8; 
        10'b1000110001: data <= 15'h7ffb; 
        10'b1000110010: data <= 15'h7fea; 
        10'b1000110011: data <= 15'h7fe0; 
        10'b1000110100: data <= 15'h7fc0; 
        10'b1000110101: data <= 15'h7ff5; 
        10'b1000110110: data <= 15'h000a; 
        10'b1000110111: data <= 15'h005a; 
        10'b1000111000: data <= 15'h001b; 
        10'b1000111001: data <= 15'h7ff4; 
        10'b1000111010: data <= 15'h7fff; 
        10'b1000111011: data <= 15'h7fb3; 
        10'b1000111100: data <= 15'h0005; 
        10'b1000111101: data <= 15'h7ffe; 
        10'b1000111110: data <= 15'h7fb7; 
        10'b1000111111: data <= 15'h7ff3; 
        10'b1001000000: data <= 15'h7fab; 
        10'b1001000001: data <= 15'h7fe5; 
        10'b1001000010: data <= 15'h000f; 
        10'b1001000011: data <= 15'h0009; 
        10'b1001000100: data <= 15'h001b; 
        10'b1001000101: data <= 15'h002e; 
        10'b1001000110: data <= 15'h002d; 
        10'b1001000111: data <= 15'h7ff5; 
        10'b1001001000: data <= 15'h7fe2; 
        10'b1001001001: data <= 15'h7fd9; 
        10'b1001001010: data <= 15'h7ff4; 
        10'b1001001011: data <= 15'h7fe9; 
        10'b1001001100: data <= 15'h0002; 
        10'b1001001101: data <= 15'h7ff3; 
        10'b1001001110: data <= 15'h0004; 
        10'b1001001111: data <= 15'h7fce; 
        10'b1001010000: data <= 15'h7fb6; 
        10'b1001010001: data <= 15'h7ff9; 
        10'b1001010010: data <= 15'h0027; 
        10'b1001010011: data <= 15'h0054; 
        10'b1001010100: data <= 15'h0012; 
        10'b1001010101: data <= 15'h0024; 
        10'b1001010110: data <= 15'h7ff9; 
        10'b1001010111: data <= 15'h7fc9; 
        10'b1001011000: data <= 15'h7fe1; 
        10'b1001011001: data <= 15'h0013; 
        10'b1001011010: data <= 15'h7ffe; 
        10'b1001011011: data <= 15'h7ff7; 
        10'b1001011100: data <= 15'h7fbf; 
        10'b1001011101: data <= 15'h7fe5; 
        10'b1001011110: data <= 15'h7fee; 
        10'b1001011111: data <= 15'h7ffd; 
        10'b1001100000: data <= 15'h7ffe; 
        10'b1001100001: data <= 15'h0010; 
        10'b1001100010: data <= 15'h000d; 
        10'b1001100011: data <= 15'h7fec; 
        10'b1001100100: data <= 15'h7fe8; 
        10'b1001100101: data <= 15'h7fff; 
        10'b1001100110: data <= 15'h7ffb; 
        10'b1001100111: data <= 15'h7ff1; 
        10'b1001101000: data <= 15'h7ff8; 
        10'b1001101001: data <= 15'h7fe4; 
        10'b1001101010: data <= 15'h7fee; 
        10'b1001101011: data <= 15'h7fe0; 
        10'b1001101100: data <= 15'h7fc5; 
        10'b1001101101: data <= 15'h7fa7; 
        10'b1001101110: data <= 15'h000b; 
        10'b1001101111: data <= 15'h0018; 
        10'b1001110000: data <= 15'h7ffb; 
        10'b1001110001: data <= 15'h7fe4; 
        10'b1001110010: data <= 15'h0012; 
        10'b1001110011: data <= 15'h0006; 
        10'b1001110100: data <= 15'h006a; 
        10'b1001110101: data <= 15'h006f; 
        10'b1001110110: data <= 15'h004e; 
        10'b1001110111: data <= 15'h003d; 
        10'b1001111000: data <= 15'h7ffb; 
        10'b1001111001: data <= 15'h7ffa; 
        10'b1001111010: data <= 15'h001a; 
        10'b1001111011: data <= 15'h7fdf; 
        10'b1001111100: data <= 15'h7fdc; 
        10'b1001111101: data <= 15'h000f; 
        10'b1001111110: data <= 15'h7ffa; 
        10'b1001111111: data <= 15'h7fe9; 
        10'b1010000000: data <= 15'h7ffa; 
        10'b1010000001: data <= 15'h7ffa; 
        10'b1010000010: data <= 15'h7ff9; 
        10'b1010000011: data <= 15'h7fea; 
        10'b1010000100: data <= 15'h7fea; 
        10'b1010000101: data <= 15'h7ffd; 
        10'b1010000110: data <= 15'h7ff6; 
        10'b1010000111: data <= 15'h7fe4; 
        10'b1010001000: data <= 15'h7fc2; 
        10'b1010001001: data <= 15'h7f6c; 
        10'b1010001010: data <= 15'h7f8c; 
        10'b1010001011: data <= 15'h7fc6; 
        10'b1010001100: data <= 15'h0014; 
        10'b1010001101: data <= 15'h0014; 
        10'b1010001110: data <= 15'h002b; 
        10'b1010001111: data <= 15'h0038; 
        10'b1010010000: data <= 15'h007d; 
        10'b1010010001: data <= 15'h00b4; 
        10'b1010010010: data <= 15'h0099; 
        10'b1010010011: data <= 15'h007a; 
        10'b1010010100: data <= 15'h0063; 
        10'b1010010101: data <= 15'h0047; 
        10'b1010010110: data <= 15'h0038; 
        10'b1010010111: data <= 15'h0048; 
        10'b1010011000: data <= 15'h0035; 
        10'b1010011001: data <= 15'h000d; 
        10'b1010011010: data <= 15'h7ff9; 
        10'b1010011011: data <= 15'h7fef; 
        10'b1010011100: data <= 15'h7fdf; 
        10'b1010011101: data <= 15'h7ffd; 
        10'b1010011110: data <= 15'h7fe3; 
        10'b1010011111: data <= 15'h7ffa; 
        10'b1010100000: data <= 15'h7ffc; 
        10'b1010100001: data <= 15'h7ffa; 
        10'b1010100010: data <= 15'h0006; 
        10'b1010100011: data <= 15'h7fe7; 
        10'b1010100100: data <= 15'h7fe6; 
        10'b1010100101: data <= 15'h7f9e; 
        10'b1010100110: data <= 15'h7f78; 
        10'b1010100111: data <= 15'h7f8e; 
        10'b1010101000: data <= 15'h7ff9; 
        10'b1010101001: data <= 15'h001b; 
        10'b1010101010: data <= 15'h7ff6; 
        10'b1010101011: data <= 15'h0030; 
        10'b1010101100: data <= 15'h0024; 
        10'b1010101101: data <= 15'h0018; 
        10'b1010101110: data <= 15'h003b; 
        10'b1010101111: data <= 15'h0081; 
        10'b1010110000: data <= 15'h0089; 
        10'b1010110001: data <= 15'h005c; 
        10'b1010110010: data <= 15'h0081; 
        10'b1010110011: data <= 15'h0079; 
        10'b1010110100: data <= 15'h0028; 
        10'b1010110101: data <= 15'h0002; 
        10'b1010110110: data <= 15'h7fe5; 
        10'b1010110111: data <= 15'h0003; 
        10'b1010111000: data <= 15'h7ff5; 
        10'b1010111001: data <= 15'h7fed; 
        10'b1010111010: data <= 15'h0004; 
        10'b1010111011: data <= 15'h7ff9; 
        10'b1010111100: data <= 15'h0006; 
        10'b1010111101: data <= 15'h7ffc; 
        10'b1010111110: data <= 15'h0003; 
        10'b1010111111: data <= 15'h7fe6; 
        10'b1011000000: data <= 15'h7fed; 
        10'b1011000001: data <= 15'h7fdc; 
        10'b1011000010: data <= 15'h7fcd; 
        10'b1011000011: data <= 15'h7fc0; 
        10'b1011000100: data <= 15'h7fb9; 
        10'b1011000101: data <= 15'h7fb9; 
        10'b1011000110: data <= 15'h7fe5; 
        10'b1011000111: data <= 15'h7fce; 
        10'b1011001000: data <= 15'h7fe2; 
        10'b1011001001: data <= 15'h7fe2; 
        10'b1011001010: data <= 15'h7ffd; 
        10'b1011001011: data <= 15'h002d; 
        10'b1011001100: data <= 15'h0020; 
        10'b1011001101: data <= 15'h0029; 
        10'b1011001110: data <= 15'h002f; 
        10'b1011001111: data <= 15'h0007; 
        10'b1011010000: data <= 15'h7ff6; 
        10'b1011010001: data <= 15'h7fff; 
        10'b1011010010: data <= 15'h7fe1; 
        10'b1011010011: data <= 15'h7fe2; 
        10'b1011010100: data <= 15'h7ffd; 
        10'b1011010101: data <= 15'h7ff8; 
        10'b1011010110: data <= 15'h7fed; 
        10'b1011010111: data <= 15'h7ff7; 
        10'b1011011000: data <= 15'h7ffb; 
        10'b1011011001: data <= 15'h0001; 
        10'b1011011010: data <= 15'h7ff2; 
        10'b1011011011: data <= 15'h7feb; 
        10'b1011011100: data <= 15'h7fe2; 
        10'b1011011101: data <= 15'h7fe7; 
        10'b1011011110: data <= 15'h7fd9; 
        10'b1011011111: data <= 15'h7ff5; 
        10'b1011100000: data <= 15'h7fdd; 
        10'b1011100001: data <= 15'h7fe2; 
        10'b1011100010: data <= 15'h7fdc; 
        10'b1011100011: data <= 15'h7feb; 
        10'b1011100100: data <= 15'h7fe9; 
        10'b1011100101: data <= 15'h7fed; 
        10'b1011100110: data <= 15'h7fe3; 
        10'b1011100111: data <= 15'h7feb; 
        10'b1011101000: data <= 15'h7fe7; 
        10'b1011101001: data <= 15'h7fdf; 
        10'b1011101010: data <= 15'h7fdb; 
        10'b1011101011: data <= 15'h7fe9; 
        10'b1011101100: data <= 15'h7ff0; 
        10'b1011101101: data <= 15'h7ffb; 
        10'b1011101110: data <= 15'h7ff1; 
        10'b1011101111: data <= 15'h0007; 
        10'b1011110000: data <= 15'h0006; 
        10'b1011110001: data <= 15'h7fe4; 
        10'b1011110010: data <= 15'h7ff7; 
        10'b1011110011: data <= 15'h7ff4; 
        10'b1011110100: data <= 15'h7ffa; 
        10'b1011110101: data <= 15'h7fea; 
        10'b1011110110: data <= 15'h7ff3; 
        10'b1011110111: data <= 15'h7ff7; 
        10'b1011111000: data <= 15'h7ff9; 
        10'b1011111001: data <= 15'h7fe3; 
        10'b1011111010: data <= 15'h7fff; 
        10'b1011111011: data <= 15'h7fed; 
        10'b1011111100: data <= 15'h0005; 
        10'b1011111101: data <= 15'h7ff2; 
        10'b1011111110: data <= 15'h7fe7; 
        10'b1011111111: data <= 15'h7ffd; 
        10'b1100000000: data <= 15'h7fec; 
        10'b1100000001: data <= 15'h7fe8; 
        10'b1100000010: data <= 15'h7ff1; 
        10'b1100000011: data <= 15'h7ffa; 
        10'b1100000100: data <= 15'h7ff7; 
        10'b1100000101: data <= 15'h0001; 
        10'b1100000110: data <= 15'h0004; 
        10'b1100000111: data <= 15'h0006; 
        10'b1100001000: data <= 15'h7ffb; 
        10'b1100001001: data <= 15'h7ff8; 
        10'b1100001010: data <= 15'h7ffb; 
        10'b1100001011: data <= 15'h7fea; 
        10'b1100001100: data <= 15'h7ff6; 
        10'b1100001101: data <= 15'h0004; 
        10'b1100001110: data <= 15'h7fe5; 
        10'b1100001111: data <= 15'h7ff6; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 10) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 16'hffe3; 
        10'b0000000001: data <= 16'hffe9; 
        10'b0000000010: data <= 16'hffe4; 
        10'b0000000011: data <= 16'hfff3; 
        10'b0000000100: data <= 16'hffef; 
        10'b0000000101: data <= 16'h0006; 
        10'b0000000110: data <= 16'hffc5; 
        10'b0000000111: data <= 16'hfff3; 
        10'b0000001000: data <= 16'hffd9; 
        10'b0000001001: data <= 16'hffdf; 
        10'b0000001010: data <= 16'hffd1; 
        10'b0000001011: data <= 16'h0005; 
        10'b0000001100: data <= 16'hffed; 
        10'b0000001101: data <= 16'hfffd; 
        10'b0000001110: data <= 16'hffcf; 
        10'b0000001111: data <= 16'hfffd; 
        10'b0000010000: data <= 16'hfff1; 
        10'b0000010001: data <= 16'hffcb; 
        10'b0000010010: data <= 16'h0005; 
        10'b0000010011: data <= 16'hffe9; 
        10'b0000010100: data <= 16'hffe4; 
        10'b0000010101: data <= 16'hffe3; 
        10'b0000010110: data <= 16'hffe7; 
        10'b0000010111: data <= 16'h000b; 
        10'b0000011000: data <= 16'h0000; 
        10'b0000011001: data <= 16'hffde; 
        10'b0000011010: data <= 16'hffd6; 
        10'b0000011011: data <= 16'hffe6; 
        10'b0000011100: data <= 16'hffe4; 
        10'b0000011101: data <= 16'hffc6; 
        10'b0000011110: data <= 16'h000a; 
        10'b0000011111: data <= 16'h0000; 
        10'b0000100000: data <= 16'hffcb; 
        10'b0000100001: data <= 16'hffcc; 
        10'b0000100010: data <= 16'hffc7; 
        10'b0000100011: data <= 16'hffcc; 
        10'b0000100100: data <= 16'h0007; 
        10'b0000100101: data <= 16'hffea; 
        10'b0000100110: data <= 16'hffe8; 
        10'b0000100111: data <= 16'hffc6; 
        10'b0000101000: data <= 16'h0006; 
        10'b0000101001: data <= 16'hfff7; 
        10'b0000101010: data <= 16'hffd8; 
        10'b0000101011: data <= 16'hffe2; 
        10'b0000101100: data <= 16'hfff7; 
        10'b0000101101: data <= 16'hffed; 
        10'b0000101110: data <= 16'hffd3; 
        10'b0000101111: data <= 16'hffef; 
        10'b0000110000: data <= 16'h0006; 
        10'b0000110001: data <= 16'hffc9; 
        10'b0000110010: data <= 16'hfff6; 
        10'b0000110011: data <= 16'hffd3; 
        10'b0000110100: data <= 16'hfffc; 
        10'b0000110101: data <= 16'h000c; 
        10'b0000110110: data <= 16'hffd8; 
        10'b0000110111: data <= 16'hffd3; 
        10'b0000111000: data <= 16'hffcf; 
        10'b0000111001: data <= 16'hffff; 
        10'b0000111010: data <= 16'hffec; 
        10'b0000111011: data <= 16'hffe8; 
        10'b0000111100: data <= 16'hffd1; 
        10'b0000111101: data <= 16'hffc7; 
        10'b0000111110: data <= 16'hffed; 
        10'b0000111111: data <= 16'hffc5; 
        10'b0001000000: data <= 16'h000a; 
        10'b0001000001: data <= 16'hffc5; 
        10'b0001000010: data <= 16'hffc8; 
        10'b0001000011: data <= 16'hfff4; 
        10'b0001000100: data <= 16'hffec; 
        10'b0001000101: data <= 16'hffc3; 
        10'b0001000110: data <= 16'hfff4; 
        10'b0001000111: data <= 16'hfff0; 
        10'b0001001000: data <= 16'hffc0; 
        10'b0001001001: data <= 16'hffda; 
        10'b0001001010: data <= 16'hffda; 
        10'b0001001011: data <= 16'hfff8; 
        10'b0001001100: data <= 16'hfffe; 
        10'b0001001101: data <= 16'hfffd; 
        10'b0001001110: data <= 16'hfff2; 
        10'b0001001111: data <= 16'hffe6; 
        10'b0001010000: data <= 16'h0006; 
        10'b0001010001: data <= 16'hffd8; 
        10'b0001010010: data <= 16'hfff7; 
        10'b0001010011: data <= 16'h0008; 
        10'b0001010100: data <= 16'hffd4; 
        10'b0001010101: data <= 16'hffe7; 
        10'b0001010110: data <= 16'hffe7; 
        10'b0001010111: data <= 16'hffcd; 
        10'b0001011000: data <= 16'h000a; 
        10'b0001011001: data <= 16'hffd0; 
        10'b0001011010: data <= 16'hffc9; 
        10'b0001011011: data <= 16'hffdf; 
        10'b0001011100: data <= 16'hffc6; 
        10'b0001011101: data <= 16'hffec; 
        10'b0001011110: data <= 16'hffd5; 
        10'b0001011111: data <= 16'hffb0; 
        10'b0001100000: data <= 16'hffa7; 
        10'b0001100001: data <= 16'hff94; 
        10'b0001100010: data <= 16'hffa6; 
        10'b0001100011: data <= 16'hffcb; 
        10'b0001100100: data <= 16'hffa6; 
        10'b0001100101: data <= 16'hffba; 
        10'b0001100110: data <= 16'hffcf; 
        10'b0001100111: data <= 16'hffe2; 
        10'b0001101000: data <= 16'hffbc; 
        10'b0001101001: data <= 16'h0004; 
        10'b0001101010: data <= 16'hffdc; 
        10'b0001101011: data <= 16'hfffc; 
        10'b0001101100: data <= 16'hffd9; 
        10'b0001101101: data <= 16'hfff4; 
        10'b0001101110: data <= 16'hffee; 
        10'b0001101111: data <= 16'hffca; 
        10'b0001110000: data <= 16'hffe9; 
        10'b0001110001: data <= 16'hfff9; 
        10'b0001110010: data <= 16'hffde; 
        10'b0001110011: data <= 16'hffca; 
        10'b0001110100: data <= 16'hfffd; 
        10'b0001110101: data <= 16'hfffc; 
        10'b0001110110: data <= 16'hffe9; 
        10'b0001110111: data <= 16'hffcf; 
        10'b0001111000: data <= 16'hffcf; 
        10'b0001111001: data <= 16'hffe3; 
        10'b0001111010: data <= 16'hffe7; 
        10'b0001111011: data <= 16'hfff2; 
        10'b0001111100: data <= 16'h004e; 
        10'b0001111101: data <= 16'h0032; 
        10'b0001111110: data <= 16'h00aa; 
        10'b0001111111: data <= 16'h0081; 
        10'b0010000000: data <= 16'h003a; 
        10'b0010000001: data <= 16'h0020; 
        10'b0010000010: data <= 16'h0030; 
        10'b0010000011: data <= 16'hffd5; 
        10'b0010000100: data <= 16'hffcc; 
        10'b0010000101: data <= 16'hffe5; 
        10'b0010000110: data <= 16'hffb2; 
        10'b0010000111: data <= 16'hffc8; 
        10'b0010001000: data <= 16'hfffe; 
        10'b0010001001: data <= 16'h0004; 
        10'b0010001010: data <= 16'hffe2; 
        10'b0010001011: data <= 16'hffe9; 
        10'b0010001100: data <= 16'hffea; 
        10'b0010001101: data <= 16'hfff5; 
        10'b0010001110: data <= 16'hfff9; 
        10'b0010001111: data <= 16'hfffe; 
        10'b0010010000: data <= 16'hffd2; 
        10'b0010010001: data <= 16'hffe5; 
        10'b0010010010: data <= 16'hffd8; 
        10'b0010010011: data <= 16'hff94; 
        10'b0010010100: data <= 16'hffd5; 
        10'b0010010101: data <= 16'h0026; 
        10'b0010010110: data <= 16'hffa7; 
        10'b0010010111: data <= 16'h0076; 
        10'b0010011000: data <= 16'h00df; 
        10'b0010011001: data <= 16'h00b9; 
        10'b0010011010: data <= 16'h00c1; 
        10'b0010011011: data <= 16'h005c; 
        10'b0010011100: data <= 16'h004c; 
        10'b0010011101: data <= 16'h00b2; 
        10'b0010011110: data <= 16'h0009; 
        10'b0010011111: data <= 16'hfff8; 
        10'b0010100000: data <= 16'h0040; 
        10'b0010100001: data <= 16'h0021; 
        10'b0010100010: data <= 16'hff94; 
        10'b0010100011: data <= 16'hffa5; 
        10'b0010100100: data <= 16'hffc1; 
        10'b0010100101: data <= 16'h0030; 
        10'b0010100110: data <= 16'hffec; 
        10'b0010100111: data <= 16'h0008; 
        10'b0010101000: data <= 16'hffd4; 
        10'b0010101001: data <= 16'hffd0; 
        10'b0010101010: data <= 16'hffc6; 
        10'b0010101011: data <= 16'hffc8; 
        10'b0010101100: data <= 16'hffbf; 
        10'b0010101101: data <= 16'hffc1; 
        10'b0010101110: data <= 16'hff9a; 
        10'b0010101111: data <= 16'hff9a; 
        10'b0010110000: data <= 16'h0007; 
        10'b0010110001: data <= 16'h001e; 
        10'b0010110010: data <= 16'hfff8; 
        10'b0010110011: data <= 16'h0039; 
        10'b0010110100: data <= 16'h005b; 
        10'b0010110101: data <= 16'h0049; 
        10'b0010110110: data <= 16'h0066; 
        10'b0010110111: data <= 16'h00c0; 
        10'b0010111000: data <= 16'h005d; 
        10'b0010111001: data <= 16'h006d; 
        10'b0010111010: data <= 16'h0017; 
        10'b0010111011: data <= 16'h007d; 
        10'b0010111100: data <= 16'h0030; 
        10'b0010111101: data <= 16'h003a; 
        10'b0010111110: data <= 16'h0049; 
        10'b0010111111: data <= 16'h0044; 
        10'b0011000000: data <= 16'h0039; 
        10'b0011000001: data <= 16'h0018; 
        10'b0011000010: data <= 16'hffe9; 
        10'b0011000011: data <= 16'hfffa; 
        10'b0011000100: data <= 16'h0008; 
        10'b0011000101: data <= 16'hffd5; 
        10'b0011000110: data <= 16'hffcd; 
        10'b0011000111: data <= 16'hffd8; 
        10'b0011001000: data <= 16'hffbc; 
        10'b0011001001: data <= 16'hffe7; 
        10'b0011001010: data <= 16'hffbb; 
        10'b0011001011: data <= 16'hfffc; 
        10'b0011001100: data <= 16'h0045; 
        10'b0011001101: data <= 16'h001c; 
        10'b0011001110: data <= 16'h0022; 
        10'b0011001111: data <= 16'hffea; 
        10'b0011010000: data <= 16'hffa8; 
        10'b0011010001: data <= 16'hffbe; 
        10'b0011010010: data <= 16'hff9f; 
        10'b0011010011: data <= 16'h003a; 
        10'b0011010100: data <= 16'h0049; 
        10'b0011010101: data <= 16'hfffb; 
        10'b0011010110: data <= 16'h0032; 
        10'b0011010111: data <= 16'hffca; 
        10'b0011011000: data <= 16'h004a; 
        10'b0011011001: data <= 16'h0074; 
        10'b0011011010: data <= 16'h0015; 
        10'b0011011011: data <= 16'h00f0; 
        10'b0011011100: data <= 16'h0093; 
        10'b0011011101: data <= 16'hfffa; 
        10'b0011011110: data <= 16'h0004; 
        10'b0011011111: data <= 16'hfff6; 
        10'b0011100000: data <= 16'hfff6; 
        10'b0011100001: data <= 16'h0003; 
        10'b0011100010: data <= 16'hfff4; 
        10'b0011100011: data <= 16'hffd1; 
        10'b0011100100: data <= 16'hfff3; 
        10'b0011100101: data <= 16'hffea; 
        10'b0011100110: data <= 16'h0064; 
        10'b0011100111: data <= 16'h003d; 
        10'b0011101000: data <= 16'h0016; 
        10'b0011101001: data <= 16'h00ad; 
        10'b0011101010: data <= 16'h000a; 
        10'b0011101011: data <= 16'h0006; 
        10'b0011101100: data <= 16'h0073; 
        10'b0011101101: data <= 16'h0095; 
        10'b0011101110: data <= 16'hff8a; 
        10'b0011101111: data <= 16'hff9c; 
        10'b0011110000: data <= 16'h0052; 
        10'b0011110001: data <= 16'hffc6; 
        10'b0011110010: data <= 16'h001b; 
        10'b0011110011: data <= 16'h004e; 
        10'b0011110100: data <= 16'h0034; 
        10'b0011110101: data <= 16'h009f; 
        10'b0011110110: data <= 16'h006b; 
        10'b0011110111: data <= 16'h00b5; 
        10'b0011111000: data <= 16'h00a5; 
        10'b0011111001: data <= 16'hffec; 
        10'b0011111010: data <= 16'hfff2; 
        10'b0011111011: data <= 16'h0010; 
        10'b0011111100: data <= 16'h0001; 
        10'b0011111101: data <= 16'h0003; 
        10'b0011111110: data <= 16'hffe6; 
        10'b0011111111: data <= 16'hffe0; 
        10'b0100000000: data <= 16'hffef; 
        10'b0100000001: data <= 16'h0065; 
        10'b0100000010: data <= 16'h004b; 
        10'b0100000011: data <= 16'h009a; 
        10'b0100000100: data <= 16'h00cf; 
        10'b0100000101: data <= 16'h00ae; 
        10'b0100000110: data <= 16'h006e; 
        10'b0100000111: data <= 16'h00c2; 
        10'b0100001000: data <= 16'h0035; 
        10'b0100001001: data <= 16'h0038; 
        10'b0100001010: data <= 16'hff1d; 
        10'b0100001011: data <= 16'hfec4; 
        10'b0100001100: data <= 16'hff92; 
        10'b0100001101: data <= 16'h0011; 
        10'b0100001110: data <= 16'h0022; 
        10'b0100001111: data <= 16'h003d; 
        10'b0100010000: data <= 16'h0051; 
        10'b0100010001: data <= 16'h0046; 
        10'b0100010010: data <= 16'h00a7; 
        10'b0100010011: data <= 16'h00ab; 
        10'b0100010100: data <= 16'hffe4; 
        10'b0100010101: data <= 16'hffe8; 
        10'b0100010110: data <= 16'h0026; 
        10'b0100010111: data <= 16'hffcc; 
        10'b0100011000: data <= 16'hffd6; 
        10'b0100011001: data <= 16'h0002; 
        10'b0100011010: data <= 16'hffd4; 
        10'b0100011011: data <= 16'h0004; 
        10'b0100011100: data <= 16'h0027; 
        10'b0100011101: data <= 16'h007c; 
        10'b0100011110: data <= 16'h007b; 
        10'b0100011111: data <= 16'h00e2; 
        10'b0100100000: data <= 16'h00a7; 
        10'b0100100001: data <= 16'h00c4; 
        10'b0100100010: data <= 16'h011e; 
        10'b0100100011: data <= 16'h0089; 
        10'b0100100100: data <= 16'h008f; 
        10'b0100100101: data <= 16'h0075; 
        10'b0100100110: data <= 16'hffda; 
        10'b0100100111: data <= 16'hfed4; 
        10'b0100101000: data <= 16'hff0a; 
        10'b0100101001: data <= 16'hffb5; 
        10'b0100101010: data <= 16'h0056; 
        10'b0100101011: data <= 16'h0055; 
        10'b0100101100: data <= 16'h0057; 
        10'b0100101101: data <= 16'h00cb; 
        10'b0100101110: data <= 16'h00e1; 
        10'b0100101111: data <= 16'h00b8; 
        10'b0100110000: data <= 16'h0002; 
        10'b0100110001: data <= 16'hfff3; 
        10'b0100110010: data <= 16'hffe8; 
        10'b0100110011: data <= 16'hffd8; 
        10'b0100110100: data <= 16'hffd4; 
        10'b0100110101: data <= 16'h000a; 
        10'b0100110110: data <= 16'hfffc; 
        10'b0100110111: data <= 16'hffba; 
        10'b0100111000: data <= 16'h003b; 
        10'b0100111001: data <= 16'h0089; 
        10'b0100111010: data <= 16'h0104; 
        10'b0100111011: data <= 16'h0152; 
        10'b0100111100: data <= 16'h010a; 
        10'b0100111101: data <= 16'h014f; 
        10'b0100111110: data <= 16'h00e6; 
        10'b0100111111: data <= 16'h006d; 
        10'b0101000000: data <= 16'h008c; 
        10'b0101000001: data <= 16'h014e; 
        10'b0101000010: data <= 16'h0197; 
        10'b0101000011: data <= 16'hffce; 
        10'b0101000100: data <= 16'hff0e; 
        10'b0101000101: data <= 16'hffad; 
        10'b0101000110: data <= 16'hffb1; 
        10'b0101000111: data <= 16'h0021; 
        10'b0101001000: data <= 16'h00b8; 
        10'b0101001001: data <= 16'h00dc; 
        10'b0101001010: data <= 16'h0125; 
        10'b0101001011: data <= 16'h0114; 
        10'b0101001100: data <= 16'h00c0; 
        10'b0101001101: data <= 16'h001f; 
        10'b0101001110: data <= 16'h0011; 
        10'b0101001111: data <= 16'hfff0; 
        10'b0101010000: data <= 16'hffda; 
        10'b0101010001: data <= 16'hfff3; 
        10'b0101010010: data <= 16'hffe0; 
        10'b0101010011: data <= 16'hfff1; 
        10'b0101010100: data <= 16'hfff4; 
        10'b0101010101: data <= 16'h00a3; 
        10'b0101010110: data <= 16'h0087; 
        10'b0101010111: data <= 16'h00cf; 
        10'b0101011000: data <= 16'h00c3; 
        10'b0101011001: data <= 16'h00f5; 
        10'b0101011010: data <= 16'h002a; 
        10'b0101011011: data <= 16'h003b; 
        10'b0101011100: data <= 16'h0020; 
        10'b0101011101: data <= 16'h0193; 
        10'b0101011110: data <= 16'h0195; 
        10'b0101011111: data <= 16'h005b; 
        10'b0101100000: data <= 16'h000f; 
        10'b0101100001: data <= 16'hffdd; 
        10'b0101100010: data <= 16'hffe3; 
        10'b0101100011: data <= 16'h0066; 
        10'b0101100100: data <= 16'h00ac; 
        10'b0101100101: data <= 16'h0128; 
        10'b0101100110: data <= 16'h0159; 
        10'b0101100111: data <= 16'h0120; 
        10'b0101101000: data <= 16'h00b5; 
        10'b0101101001: data <= 16'h0048; 
        10'b0101101010: data <= 16'h0024; 
        10'b0101101011: data <= 16'hffcd; 
        10'b0101101100: data <= 16'hffc8; 
        10'b0101101101: data <= 16'hffec; 
        10'b0101101110: data <= 16'h000b; 
        10'b0101101111: data <= 16'hffd0; 
        10'b0101110000: data <= 16'hffdc; 
        10'b0101110001: data <= 16'hffff; 
        10'b0101110010: data <= 16'hffe6; 
        10'b0101110011: data <= 16'hffe7; 
        10'b0101110100: data <= 16'h0016; 
        10'b0101110101: data <= 16'hffe2; 
        10'b0101110110: data <= 16'hffa8; 
        10'b0101110111: data <= 16'h0022; 
        10'b0101111000: data <= 16'h0094; 
        10'b0101111001: data <= 16'h017a; 
        10'b0101111010: data <= 16'h0071; 
        10'b0101111011: data <= 16'h0116; 
        10'b0101111100: data <= 16'h006f; 
        10'b0101111101: data <= 16'hffba; 
        10'b0101111110: data <= 16'h0007; 
        10'b0101111111: data <= 16'h0009; 
        10'b0110000000: data <= 16'h007b; 
        10'b0110000001: data <= 16'h0070; 
        10'b0110000010: data <= 16'h003f; 
        10'b0110000011: data <= 16'h005a; 
        10'b0110000100: data <= 16'h0030; 
        10'b0110000101: data <= 16'h000b; 
        10'b0110000110: data <= 16'h000b; 
        10'b0110000111: data <= 16'hfff7; 
        10'b0110001000: data <= 16'hffde; 
        10'b0110001001: data <= 16'hffc7; 
        10'b0110001010: data <= 16'hfff8; 
        10'b0110001011: data <= 16'hffe8; 
        10'b0110001100: data <= 16'hffce; 
        10'b0110001101: data <= 16'hff92; 
        10'b0110001110: data <= 16'hff3c; 
        10'b0110001111: data <= 16'hff05; 
        10'b0110010000: data <= 16'hfed7; 
        10'b0110010001: data <= 16'hff12; 
        10'b0110010010: data <= 16'hffdf; 
        10'b0110010011: data <= 16'h0098; 
        10'b0110010100: data <= 16'h0092; 
        10'b0110010101: data <= 16'h0135; 
        10'b0110010110: data <= 16'h00f7; 
        10'b0110010111: data <= 16'h00a7; 
        10'b0110011000: data <= 16'hffec; 
        10'b0110011001: data <= 16'h0015; 
        10'b0110011010: data <= 16'hffd5; 
        10'b0110011011: data <= 16'hff9b; 
        10'b0110011100: data <= 16'hff5c; 
        10'b0110011101: data <= 16'hff6d; 
        10'b0110011110: data <= 16'hff82; 
        10'b0110011111: data <= 16'hff6b; 
        10'b0110100000: data <= 16'hffbc; 
        10'b0110100001: data <= 16'hfff6; 
        10'b0110100010: data <= 16'hffc4; 
        10'b0110100011: data <= 16'h0002; 
        10'b0110100100: data <= 16'h0005; 
        10'b0110100101: data <= 16'hffdb; 
        10'b0110100110: data <= 16'hffd6; 
        10'b0110100111: data <= 16'hffee; 
        10'b0110101000: data <= 16'hffc9; 
        10'b0110101001: data <= 16'hff93; 
        10'b0110101010: data <= 16'hff0c; 
        10'b0110101011: data <= 16'hfed5; 
        10'b0110101100: data <= 16'hfeef; 
        10'b0110101101: data <= 16'hffbd; 
        10'b0110101110: data <= 16'h000a; 
        10'b0110101111: data <= 16'h0007; 
        10'b0110110000: data <= 16'h00d3; 
        10'b0110110001: data <= 16'h00f9; 
        10'b0110110010: data <= 16'h00da; 
        10'b0110110011: data <= 16'h007e; 
        10'b0110110100: data <= 16'hffc1; 
        10'b0110110101: data <= 16'hffc9; 
        10'b0110110110: data <= 16'hffd9; 
        10'b0110110111: data <= 16'hff23; 
        10'b0110111000: data <= 16'hfeed; 
        10'b0110111001: data <= 16'hff2d; 
        10'b0110111010: data <= 16'hff7a; 
        10'b0110111011: data <= 16'hff81; 
        10'b0110111100: data <= 16'hffa0; 
        10'b0110111101: data <= 16'hffef; 
        10'b0110111110: data <= 16'hffbe; 
        10'b0110111111: data <= 16'h0005; 
        10'b0111000000: data <= 16'hffe2; 
        10'b0111000001: data <= 16'hffc9; 
        10'b0111000010: data <= 16'hffda; 
        10'b0111000011: data <= 16'hffec; 
        10'b0111000100: data <= 16'hffa8; 
        10'b0111000101: data <= 16'hff62; 
        10'b0111000110: data <= 16'hff02; 
        10'b0111000111: data <= 16'hff6a; 
        10'b0111001000: data <= 16'h0065; 
        10'b0111001001: data <= 16'h0070; 
        10'b0111001010: data <= 16'h002e; 
        10'b0111001011: data <= 16'h0066; 
        10'b0111001100: data <= 16'h00cc; 
        10'b0111001101: data <= 16'h00b3; 
        10'b0111001110: data <= 16'h0040; 
        10'b0111001111: data <= 16'h006b; 
        10'b0111010000: data <= 16'h0024; 
        10'b0111010001: data <= 16'hffac; 
        10'b0111010010: data <= 16'hff4e; 
        10'b0111010011: data <= 16'hff01; 
        10'b0111010100: data <= 16'hff01; 
        10'b0111010101: data <= 16'hfefd; 
        10'b0111010110: data <= 16'hff30; 
        10'b0111010111: data <= 16'hffbb; 
        10'b0111011000: data <= 16'hffa5; 
        10'b0111011001: data <= 16'hffe1; 
        10'b0111011010: data <= 16'hffe0; 
        10'b0111011011: data <= 16'hffc8; 
        10'b0111011100: data <= 16'h000c; 
        10'b0111011101: data <= 16'h0009; 
        10'b0111011110: data <= 16'hffd4; 
        10'b0111011111: data <= 16'hffcb; 
        10'b0111100000: data <= 16'hffc6; 
        10'b0111100001: data <= 16'hff5d; 
        10'b0111100010: data <= 16'hff20; 
        10'b0111100011: data <= 16'h0028; 
        10'b0111100100: data <= 16'h00d0; 
        10'b0111100101: data <= 16'h0102; 
        10'b0111100110: data <= 16'h0053; 
        10'b0111100111: data <= 16'h00c3; 
        10'b0111101000: data <= 16'h013e; 
        10'b0111101001: data <= 16'h00c1; 
        10'b0111101010: data <= 16'h0010; 
        10'b0111101011: data <= 16'hffcc; 
        10'b0111101100: data <= 16'h0017; 
        10'b0111101101: data <= 16'hff9d; 
        10'b0111101110: data <= 16'hfefa; 
        10'b0111101111: data <= 16'hff84; 
        10'b0111110000: data <= 16'hff85; 
        10'b0111110001: data <= 16'hff52; 
        10'b0111110010: data <= 16'hff7f; 
        10'b0111110011: data <= 16'hffaf; 
        10'b0111110100: data <= 16'hffd2; 
        10'b0111110101: data <= 16'hffbe; 
        10'b0111110110: data <= 16'hfff5; 
        10'b0111110111: data <= 16'hffde; 
        10'b0111111000: data <= 16'hffd8; 
        10'b0111111001: data <= 16'h0003; 
        10'b0111111010: data <= 16'hffc7; 
        10'b0111111011: data <= 16'hffb7; 
        10'b0111111100: data <= 16'hff9c; 
        10'b0111111101: data <= 16'hff9a; 
        10'b0111111110: data <= 16'hffc1; 
        10'b0111111111: data <= 16'h003e; 
        10'b1000000000: data <= 16'h00ab; 
        10'b1000000001: data <= 16'h0135; 
        10'b1000000010: data <= 16'h00d8; 
        10'b1000000011: data <= 16'h0126; 
        10'b1000000100: data <= 16'h00c0; 
        10'b1000000101: data <= 16'h006e; 
        10'b1000000110: data <= 16'hff7a; 
        10'b1000000111: data <= 16'hffdd; 
        10'b1000001000: data <= 16'hffb5; 
        10'b1000001001: data <= 16'hff37; 
        10'b1000001010: data <= 16'hffd0; 
        10'b1000001011: data <= 16'hffda; 
        10'b1000001100: data <= 16'h000f; 
        10'b1000001101: data <= 16'hff91; 
        10'b1000001110: data <= 16'hffef; 
        10'b1000001111: data <= 16'hffa2; 
        10'b1000010000: data <= 16'hff80; 
        10'b1000010001: data <= 16'hffbe; 
        10'b1000010010: data <= 16'hfff5; 
        10'b1000010011: data <= 16'h0008; 
        10'b1000010100: data <= 16'hffd9; 
        10'b1000010101: data <= 16'hffed; 
        10'b1000010110: data <= 16'hfff2; 
        10'b1000010111: data <= 16'hffa9; 
        10'b1000011000: data <= 16'hff92; 
        10'b1000011001: data <= 16'hffd4; 
        10'b1000011010: data <= 16'h001d; 
        10'b1000011011: data <= 16'h0052; 
        10'b1000011100: data <= 16'h0055; 
        10'b1000011101: data <= 16'h00d1; 
        10'b1000011110: data <= 16'h006b; 
        10'b1000011111: data <= 16'hfff1; 
        10'b1000100000: data <= 16'h0033; 
        10'b1000100001: data <= 16'hff74; 
        10'b1000100010: data <= 16'hff5c; 
        10'b1000100011: data <= 16'hffc1; 
        10'b1000100100: data <= 16'hffcd; 
        10'b1000100101: data <= 16'hffbd; 
        10'b1000100110: data <= 16'h0034; 
        10'b1000100111: data <= 16'h000f; 
        10'b1000101000: data <= 16'h0042; 
        10'b1000101001: data <= 16'h0006; 
        10'b1000101010: data <= 16'h002b; 
        10'b1000101011: data <= 16'hffdb; 
        10'b1000101100: data <= 16'hff9f; 
        10'b1000101101: data <= 16'hffc6; 
        10'b1000101110: data <= 16'hffce; 
        10'b1000101111: data <= 16'h0006; 
        10'b1000110000: data <= 16'hffd0; 
        10'b1000110001: data <= 16'hfff6; 
        10'b1000110010: data <= 16'hffd4; 
        10'b1000110011: data <= 16'hffc0; 
        10'b1000110100: data <= 16'hff80; 
        10'b1000110101: data <= 16'hffea; 
        10'b1000110110: data <= 16'h0014; 
        10'b1000110111: data <= 16'h00b5; 
        10'b1000111000: data <= 16'h0036; 
        10'b1000111001: data <= 16'hffe9; 
        10'b1000111010: data <= 16'hffff; 
        10'b1000111011: data <= 16'hff67; 
        10'b1000111100: data <= 16'h000a; 
        10'b1000111101: data <= 16'hfffc; 
        10'b1000111110: data <= 16'hff6f; 
        10'b1000111111: data <= 16'hffe6; 
        10'b1001000000: data <= 16'hff56; 
        10'b1001000001: data <= 16'hffca; 
        10'b1001000010: data <= 16'h001e; 
        10'b1001000011: data <= 16'h0013; 
        10'b1001000100: data <= 16'h0036; 
        10'b1001000101: data <= 16'h005b; 
        10'b1001000110: data <= 16'h005b; 
        10'b1001000111: data <= 16'hffea; 
        10'b1001001000: data <= 16'hffc4; 
        10'b1001001001: data <= 16'hffb1; 
        10'b1001001010: data <= 16'hffe9; 
        10'b1001001011: data <= 16'hffd2; 
        10'b1001001100: data <= 16'h0004; 
        10'b1001001101: data <= 16'hffe7; 
        10'b1001001110: data <= 16'h0009; 
        10'b1001001111: data <= 16'hff9c; 
        10'b1001010000: data <= 16'hff6b; 
        10'b1001010001: data <= 16'hfff1; 
        10'b1001010010: data <= 16'h004e; 
        10'b1001010011: data <= 16'h00a7; 
        10'b1001010100: data <= 16'h0023; 
        10'b1001010101: data <= 16'h0048; 
        10'b1001010110: data <= 16'hfff3; 
        10'b1001010111: data <= 16'hff91; 
        10'b1001011000: data <= 16'hffc2; 
        10'b1001011001: data <= 16'h0026; 
        10'b1001011010: data <= 16'hfffd; 
        10'b1001011011: data <= 16'hffef; 
        10'b1001011100: data <= 16'hff7e; 
        10'b1001011101: data <= 16'hffc9; 
        10'b1001011110: data <= 16'hffdc; 
        10'b1001011111: data <= 16'hfffb; 
        10'b1001100000: data <= 16'hfffd; 
        10'b1001100001: data <= 16'h001f; 
        10'b1001100010: data <= 16'h001b; 
        10'b1001100011: data <= 16'hffd9; 
        10'b1001100100: data <= 16'hffd1; 
        10'b1001100101: data <= 16'hfffd; 
        10'b1001100110: data <= 16'hfff6; 
        10'b1001100111: data <= 16'hffe2; 
        10'b1001101000: data <= 16'hfff1; 
        10'b1001101001: data <= 16'hffc7; 
        10'b1001101010: data <= 16'hffdc; 
        10'b1001101011: data <= 16'hffc0; 
        10'b1001101100: data <= 16'hff89; 
        10'b1001101101: data <= 16'hff4f; 
        10'b1001101110: data <= 16'h0015; 
        10'b1001101111: data <= 16'h0030; 
        10'b1001110000: data <= 16'hfff5; 
        10'b1001110001: data <= 16'hffc7; 
        10'b1001110010: data <= 16'h0024; 
        10'b1001110011: data <= 16'h000d; 
        10'b1001110100: data <= 16'h00d3; 
        10'b1001110101: data <= 16'h00de; 
        10'b1001110110: data <= 16'h009d; 
        10'b1001110111: data <= 16'h007b; 
        10'b1001111000: data <= 16'hfff5; 
        10'b1001111001: data <= 16'hfff4; 
        10'b1001111010: data <= 16'h0035; 
        10'b1001111011: data <= 16'hffbe; 
        10'b1001111100: data <= 16'hffb9; 
        10'b1001111101: data <= 16'h001e; 
        10'b1001111110: data <= 16'hfff3; 
        10'b1001111111: data <= 16'hffd3; 
        10'b1010000000: data <= 16'hfff5; 
        10'b1010000001: data <= 16'hfff4; 
        10'b1010000010: data <= 16'hfff3; 
        10'b1010000011: data <= 16'hffd4; 
        10'b1010000100: data <= 16'hffd4; 
        10'b1010000101: data <= 16'hfffa; 
        10'b1010000110: data <= 16'hffec; 
        10'b1010000111: data <= 16'hffc7; 
        10'b1010001000: data <= 16'hff84; 
        10'b1010001001: data <= 16'hfed8; 
        10'b1010001010: data <= 16'hff18; 
        10'b1010001011: data <= 16'hff8b; 
        10'b1010001100: data <= 16'h0028; 
        10'b1010001101: data <= 16'h0028; 
        10'b1010001110: data <= 16'h0056; 
        10'b1010001111: data <= 16'h0070; 
        10'b1010010000: data <= 16'h00fa; 
        10'b1010010001: data <= 16'h0168; 
        10'b1010010010: data <= 16'h0132; 
        10'b1010010011: data <= 16'h00f4; 
        10'b1010010100: data <= 16'h00c6; 
        10'b1010010101: data <= 16'h008e; 
        10'b1010010110: data <= 16'h0071; 
        10'b1010010111: data <= 16'h0090; 
        10'b1010011000: data <= 16'h006a; 
        10'b1010011001: data <= 16'h0019; 
        10'b1010011010: data <= 16'hfff3; 
        10'b1010011011: data <= 16'hffdf; 
        10'b1010011100: data <= 16'hffbf; 
        10'b1010011101: data <= 16'hfffa; 
        10'b1010011110: data <= 16'hffc6; 
        10'b1010011111: data <= 16'hfff4; 
        10'b1010100000: data <= 16'hfff9; 
        10'b1010100001: data <= 16'hfff5; 
        10'b1010100010: data <= 16'h000b; 
        10'b1010100011: data <= 16'hffcd; 
        10'b1010100100: data <= 16'hffcd; 
        10'b1010100101: data <= 16'hff3c; 
        10'b1010100110: data <= 16'hfef0; 
        10'b1010100111: data <= 16'hff1c; 
        10'b1010101000: data <= 16'hfff2; 
        10'b1010101001: data <= 16'h0035; 
        10'b1010101010: data <= 16'hffec; 
        10'b1010101011: data <= 16'h0061; 
        10'b1010101100: data <= 16'h0047; 
        10'b1010101101: data <= 16'h002f; 
        10'b1010101110: data <= 16'h0077; 
        10'b1010101111: data <= 16'h0102; 
        10'b1010110000: data <= 16'h0112; 
        10'b1010110001: data <= 16'h00b8; 
        10'b1010110010: data <= 16'h0102; 
        10'b1010110011: data <= 16'h00f2; 
        10'b1010110100: data <= 16'h0050; 
        10'b1010110101: data <= 16'h0005; 
        10'b1010110110: data <= 16'hffc9; 
        10'b1010110111: data <= 16'h0006; 
        10'b1010111000: data <= 16'hffea; 
        10'b1010111001: data <= 16'hffda; 
        10'b1010111010: data <= 16'h0009; 
        10'b1010111011: data <= 16'hfff1; 
        10'b1010111100: data <= 16'h000c; 
        10'b1010111101: data <= 16'hfff7; 
        10'b1010111110: data <= 16'h0006; 
        10'b1010111111: data <= 16'hffcd; 
        10'b1011000000: data <= 16'hffd9; 
        10'b1011000001: data <= 16'hffb7; 
        10'b1011000010: data <= 16'hff99; 
        10'b1011000011: data <= 16'hff80; 
        10'b1011000100: data <= 16'hff72; 
        10'b1011000101: data <= 16'hff71; 
        10'b1011000110: data <= 16'hffcb; 
        10'b1011000111: data <= 16'hff9b; 
        10'b1011001000: data <= 16'hffc4; 
        10'b1011001001: data <= 16'hffc3; 
        10'b1011001010: data <= 16'hfffa; 
        10'b1011001011: data <= 16'h005b; 
        10'b1011001100: data <= 16'h0041; 
        10'b1011001101: data <= 16'h0052; 
        10'b1011001110: data <= 16'h005d; 
        10'b1011001111: data <= 16'h000f; 
        10'b1011010000: data <= 16'hffec; 
        10'b1011010001: data <= 16'hfffd; 
        10'b1011010010: data <= 16'hffc2; 
        10'b1011010011: data <= 16'hffc5; 
        10'b1011010100: data <= 16'hfffb; 
        10'b1011010101: data <= 16'hfff0; 
        10'b1011010110: data <= 16'hffda; 
        10'b1011010111: data <= 16'hffee; 
        10'b1011011000: data <= 16'hfff6; 
        10'b1011011001: data <= 16'h0001; 
        10'b1011011010: data <= 16'hffe4; 
        10'b1011011011: data <= 16'hffd6; 
        10'b1011011100: data <= 16'hffc4; 
        10'b1011011101: data <= 16'hffcd; 
        10'b1011011110: data <= 16'hffb2; 
        10'b1011011111: data <= 16'hffea; 
        10'b1011100000: data <= 16'hffba; 
        10'b1011100001: data <= 16'hffc4; 
        10'b1011100010: data <= 16'hffb8; 
        10'b1011100011: data <= 16'hffd7; 
        10'b1011100100: data <= 16'hffd2; 
        10'b1011100101: data <= 16'hffd9; 
        10'b1011100110: data <= 16'hffc7; 
        10'b1011100111: data <= 16'hffd6; 
        10'b1011101000: data <= 16'hffce; 
        10'b1011101001: data <= 16'hffbd; 
        10'b1011101010: data <= 16'hffb6; 
        10'b1011101011: data <= 16'hffd1; 
        10'b1011101100: data <= 16'hffe0; 
        10'b1011101101: data <= 16'hfff6; 
        10'b1011101110: data <= 16'hffe3; 
        10'b1011101111: data <= 16'h000d; 
        10'b1011110000: data <= 16'h000c; 
        10'b1011110001: data <= 16'hffc8; 
        10'b1011110010: data <= 16'hffee; 
        10'b1011110011: data <= 16'hffe8; 
        10'b1011110100: data <= 16'hfff3; 
        10'b1011110101: data <= 16'hffd5; 
        10'b1011110110: data <= 16'hffe5; 
        10'b1011110111: data <= 16'hffef; 
        10'b1011111000: data <= 16'hfff1; 
        10'b1011111001: data <= 16'hffc7; 
        10'b1011111010: data <= 16'hfffe; 
        10'b1011111011: data <= 16'hffd9; 
        10'b1011111100: data <= 16'h0009; 
        10'b1011111101: data <= 16'hffe4; 
        10'b1011111110: data <= 16'hffce; 
        10'b1011111111: data <= 16'hfffb; 
        10'b1100000000: data <= 16'hffd8; 
        10'b1100000001: data <= 16'hffcf; 
        10'b1100000010: data <= 16'hffe2; 
        10'b1100000011: data <= 16'hfff3; 
        10'b1100000100: data <= 16'hffee; 
        10'b1100000101: data <= 16'h0001; 
        10'b1100000110: data <= 16'h0008; 
        10'b1100000111: data <= 16'h000b; 
        10'b1100001000: data <= 16'hfff6; 
        10'b1100001001: data <= 16'hfff0; 
        10'b1100001010: data <= 16'hfff6; 
        10'b1100001011: data <= 16'hffd4; 
        10'b1100001100: data <= 16'hffec; 
        10'b1100001101: data <= 16'h0008; 
        10'b1100001110: data <= 16'hffcb; 
        10'b1100001111: data <= 16'hffec; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 11) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 17'h1ffc7; 
        10'b0000000001: data <= 17'h1ffd2; 
        10'b0000000010: data <= 17'h1ffc8; 
        10'b0000000011: data <= 17'h1ffe6; 
        10'b0000000100: data <= 17'h1ffde; 
        10'b0000000101: data <= 17'h0000b; 
        10'b0000000110: data <= 17'h1ff8b; 
        10'b0000000111: data <= 17'h1ffe7; 
        10'b0000001000: data <= 17'h1ffb1; 
        10'b0000001001: data <= 17'h1ffbd; 
        10'b0000001010: data <= 17'h1ffa2; 
        10'b0000001011: data <= 17'h0000a; 
        10'b0000001100: data <= 17'h1ffdb; 
        10'b0000001101: data <= 17'h1fffa; 
        10'b0000001110: data <= 17'h1ff9e; 
        10'b0000001111: data <= 17'h1fffb; 
        10'b0000010000: data <= 17'h1ffe2; 
        10'b0000010001: data <= 17'h1ff97; 
        10'b0000010010: data <= 17'h0000b; 
        10'b0000010011: data <= 17'h1ffd2; 
        10'b0000010100: data <= 17'h1ffc9; 
        10'b0000010101: data <= 17'h1ffc5; 
        10'b0000010110: data <= 17'h1ffcd; 
        10'b0000010111: data <= 17'h00016; 
        10'b0000011000: data <= 17'h00001; 
        10'b0000011001: data <= 17'h1ffbd; 
        10'b0000011010: data <= 17'h1ffac; 
        10'b0000011011: data <= 17'h1ffcb; 
        10'b0000011100: data <= 17'h1ffc8; 
        10'b0000011101: data <= 17'h1ff8b; 
        10'b0000011110: data <= 17'h00014; 
        10'b0000011111: data <= 17'h00000; 
        10'b0000100000: data <= 17'h1ff95; 
        10'b0000100001: data <= 17'h1ff99; 
        10'b0000100010: data <= 17'h1ff8f; 
        10'b0000100011: data <= 17'h1ff99; 
        10'b0000100100: data <= 17'h0000f; 
        10'b0000100101: data <= 17'h1ffd5; 
        10'b0000100110: data <= 17'h1ffd0; 
        10'b0000100111: data <= 17'h1ff8c; 
        10'b0000101000: data <= 17'h0000d; 
        10'b0000101001: data <= 17'h1ffed; 
        10'b0000101010: data <= 17'h1ffb1; 
        10'b0000101011: data <= 17'h1ffc4; 
        10'b0000101100: data <= 17'h1ffee; 
        10'b0000101101: data <= 17'h1ffda; 
        10'b0000101110: data <= 17'h1ffa6; 
        10'b0000101111: data <= 17'h1ffde; 
        10'b0000110000: data <= 17'h0000b; 
        10'b0000110001: data <= 17'h1ff93; 
        10'b0000110010: data <= 17'h1ffec; 
        10'b0000110011: data <= 17'h1ffa7; 
        10'b0000110100: data <= 17'h1fff8; 
        10'b0000110101: data <= 17'h00018; 
        10'b0000110110: data <= 17'h1ffb1; 
        10'b0000110111: data <= 17'h1ffa6; 
        10'b0000111000: data <= 17'h1ff9e; 
        10'b0000111001: data <= 17'h1fffe; 
        10'b0000111010: data <= 17'h1ffd9; 
        10'b0000111011: data <= 17'h1ffcf; 
        10'b0000111100: data <= 17'h1ffa3; 
        10'b0000111101: data <= 17'h1ff8d; 
        10'b0000111110: data <= 17'h1ffd9; 
        10'b0000111111: data <= 17'h1ff8a; 
        10'b0001000000: data <= 17'h00015; 
        10'b0001000001: data <= 17'h1ff8a; 
        10'b0001000010: data <= 17'h1ff8f; 
        10'b0001000011: data <= 17'h1ffe9; 
        10'b0001000100: data <= 17'h1ffd8; 
        10'b0001000101: data <= 17'h1ff87; 
        10'b0001000110: data <= 17'h1ffe8; 
        10'b0001000111: data <= 17'h1ffdf; 
        10'b0001001000: data <= 17'h1ff80; 
        10'b0001001001: data <= 17'h1ffb4; 
        10'b0001001010: data <= 17'h1ffb5; 
        10'b0001001011: data <= 17'h1fff0; 
        10'b0001001100: data <= 17'h1fffc; 
        10'b0001001101: data <= 17'h1fffa; 
        10'b0001001110: data <= 17'h1ffe4; 
        10'b0001001111: data <= 17'h1ffcc; 
        10'b0001010000: data <= 17'h0000b; 
        10'b0001010001: data <= 17'h1ffb0; 
        10'b0001010010: data <= 17'h1ffee; 
        10'b0001010011: data <= 17'h0000f; 
        10'b0001010100: data <= 17'h1ffa8; 
        10'b0001010101: data <= 17'h1ffcd; 
        10'b0001010110: data <= 17'h1ffce; 
        10'b0001010111: data <= 17'h1ff9a; 
        10'b0001011000: data <= 17'h00014; 
        10'b0001011001: data <= 17'h1ffa0; 
        10'b0001011010: data <= 17'h1ff92; 
        10'b0001011011: data <= 17'h1ffbe; 
        10'b0001011100: data <= 17'h1ff8d; 
        10'b0001011101: data <= 17'h1ffd8; 
        10'b0001011110: data <= 17'h1ffa9; 
        10'b0001011111: data <= 17'h1ff5f; 
        10'b0001100000: data <= 17'h1ff4d; 
        10'b0001100001: data <= 17'h1ff27; 
        10'b0001100010: data <= 17'h1ff4c; 
        10'b0001100011: data <= 17'h1ff95; 
        10'b0001100100: data <= 17'h1ff4b; 
        10'b0001100101: data <= 17'h1ff74; 
        10'b0001100110: data <= 17'h1ff9e; 
        10'b0001100111: data <= 17'h1ffc4; 
        10'b0001101000: data <= 17'h1ff77; 
        10'b0001101001: data <= 17'h00008; 
        10'b0001101010: data <= 17'h1ffb8; 
        10'b0001101011: data <= 17'h1fff9; 
        10'b0001101100: data <= 17'h1ffb2; 
        10'b0001101101: data <= 17'h1ffe7; 
        10'b0001101110: data <= 17'h1ffdb; 
        10'b0001101111: data <= 17'h1ff95; 
        10'b0001110000: data <= 17'h1ffd1; 
        10'b0001110001: data <= 17'h1fff2; 
        10'b0001110010: data <= 17'h1ffbd; 
        10'b0001110011: data <= 17'h1ff95; 
        10'b0001110100: data <= 17'h1fffa; 
        10'b0001110101: data <= 17'h1fff8; 
        10'b0001110110: data <= 17'h1ffd1; 
        10'b0001110111: data <= 17'h1ff9f; 
        10'b0001111000: data <= 17'h1ff9f; 
        10'b0001111001: data <= 17'h1ffc7; 
        10'b0001111010: data <= 17'h1ffcd; 
        10'b0001111011: data <= 17'h1ffe4; 
        10'b0001111100: data <= 17'h0009c; 
        10'b0001111101: data <= 17'h00064; 
        10'b0001111110: data <= 17'h00153; 
        10'b0001111111: data <= 17'h00101; 
        10'b0010000000: data <= 17'h00075; 
        10'b0010000001: data <= 17'h00040; 
        10'b0010000010: data <= 17'h00060; 
        10'b0010000011: data <= 17'h1ffab; 
        10'b0010000100: data <= 17'h1ff98; 
        10'b0010000101: data <= 17'h1ffca; 
        10'b0010000110: data <= 17'h1ff63; 
        10'b0010000111: data <= 17'h1ff90; 
        10'b0010001000: data <= 17'h1fffc; 
        10'b0010001001: data <= 17'h00007; 
        10'b0010001010: data <= 17'h1ffc3; 
        10'b0010001011: data <= 17'h1ffd1; 
        10'b0010001100: data <= 17'h1ffd3; 
        10'b0010001101: data <= 17'h1ffeb; 
        10'b0010001110: data <= 17'h1fff3; 
        10'b0010001111: data <= 17'h1fffc; 
        10'b0010010000: data <= 17'h1ffa4; 
        10'b0010010001: data <= 17'h1ffc9; 
        10'b0010010010: data <= 17'h1ffb0; 
        10'b0010010011: data <= 17'h1ff29; 
        10'b0010010100: data <= 17'h1ffa9; 
        10'b0010010101: data <= 17'h0004d; 
        10'b0010010110: data <= 17'h1ff4e; 
        10'b0010010111: data <= 17'h000ed; 
        10'b0010011000: data <= 17'h001bd; 
        10'b0010011001: data <= 17'h00173; 
        10'b0010011010: data <= 17'h00182; 
        10'b0010011011: data <= 17'h000b8; 
        10'b0010011100: data <= 17'h00098; 
        10'b0010011101: data <= 17'h00165; 
        10'b0010011110: data <= 17'h00012; 
        10'b0010011111: data <= 17'h1fff0; 
        10'b0010100000: data <= 17'h0007f; 
        10'b0010100001: data <= 17'h00042; 
        10'b0010100010: data <= 17'h1ff28; 
        10'b0010100011: data <= 17'h1ff4a; 
        10'b0010100100: data <= 17'h1ff82; 
        10'b0010100101: data <= 17'h00060; 
        10'b0010100110: data <= 17'h1ffd9; 
        10'b0010100111: data <= 17'h00010; 
        10'b0010101000: data <= 17'h1ffa8; 
        10'b0010101001: data <= 17'h1ffa1; 
        10'b0010101010: data <= 17'h1ff8c; 
        10'b0010101011: data <= 17'h1ff8f; 
        10'b0010101100: data <= 17'h1ff7e; 
        10'b0010101101: data <= 17'h1ff81; 
        10'b0010101110: data <= 17'h1ff35; 
        10'b0010101111: data <= 17'h1ff34; 
        10'b0010110000: data <= 17'h0000e; 
        10'b0010110001: data <= 17'h0003c; 
        10'b0010110010: data <= 17'h1fff0; 
        10'b0010110011: data <= 17'h00073; 
        10'b0010110100: data <= 17'h000b5; 
        10'b0010110101: data <= 17'h00091; 
        10'b0010110110: data <= 17'h000cd; 
        10'b0010110111: data <= 17'h00180; 
        10'b0010111000: data <= 17'h000ba; 
        10'b0010111001: data <= 17'h000da; 
        10'b0010111010: data <= 17'h0002e; 
        10'b0010111011: data <= 17'h000f9; 
        10'b0010111100: data <= 17'h0005f; 
        10'b0010111101: data <= 17'h00075; 
        10'b0010111110: data <= 17'h00092; 
        10'b0010111111: data <= 17'h00088; 
        10'b0011000000: data <= 17'h00073; 
        10'b0011000001: data <= 17'h00030; 
        10'b0011000010: data <= 17'h1ffd1; 
        10'b0011000011: data <= 17'h1fff4; 
        10'b0011000100: data <= 17'h00011; 
        10'b0011000101: data <= 17'h1ffa9; 
        10'b0011000110: data <= 17'h1ff9a; 
        10'b0011000111: data <= 17'h1ffb0; 
        10'b0011001000: data <= 17'h1ff79; 
        10'b0011001001: data <= 17'h1ffcf; 
        10'b0011001010: data <= 17'h1ff75; 
        10'b0011001011: data <= 17'h1fff8; 
        10'b0011001100: data <= 17'h00089; 
        10'b0011001101: data <= 17'h00038; 
        10'b0011001110: data <= 17'h00045; 
        10'b0011001111: data <= 17'h1ffd5; 
        10'b0011010000: data <= 17'h1ff51; 
        10'b0011010001: data <= 17'h1ff7d; 
        10'b0011010010: data <= 17'h1ff3e; 
        10'b0011010011: data <= 17'h00074; 
        10'b0011010100: data <= 17'h00092; 
        10'b0011010101: data <= 17'h1fff7; 
        10'b0011010110: data <= 17'h00063; 
        10'b0011010111: data <= 17'h1ff94; 
        10'b0011011000: data <= 17'h00095; 
        10'b0011011001: data <= 17'h000e8; 
        10'b0011011010: data <= 17'h0002a; 
        10'b0011011011: data <= 17'h001e0; 
        10'b0011011100: data <= 17'h00126; 
        10'b0011011101: data <= 17'h1fff5; 
        10'b0011011110: data <= 17'h00007; 
        10'b0011011111: data <= 17'h1ffec; 
        10'b0011100000: data <= 17'h1ffec; 
        10'b0011100001: data <= 17'h00006; 
        10'b0011100010: data <= 17'h1ffe8; 
        10'b0011100011: data <= 17'h1ffa1; 
        10'b0011100100: data <= 17'h1ffe7; 
        10'b0011100101: data <= 17'h1ffd3; 
        10'b0011100110: data <= 17'h000c7; 
        10'b0011100111: data <= 17'h0007b; 
        10'b0011101000: data <= 17'h0002c; 
        10'b0011101001: data <= 17'h00159; 
        10'b0011101010: data <= 17'h00014; 
        10'b0011101011: data <= 17'h0000c; 
        10'b0011101100: data <= 17'h000e7; 
        10'b0011101101: data <= 17'h0012b; 
        10'b0011101110: data <= 17'h1ff14; 
        10'b0011101111: data <= 17'h1ff38; 
        10'b0011110000: data <= 17'h000a3; 
        10'b0011110001: data <= 17'h1ff8c; 
        10'b0011110010: data <= 17'h00036; 
        10'b0011110011: data <= 17'h0009c; 
        10'b0011110100: data <= 17'h00067; 
        10'b0011110101: data <= 17'h0013e; 
        10'b0011110110: data <= 17'h000d5; 
        10'b0011110111: data <= 17'h0016b; 
        10'b0011111000: data <= 17'h0014a; 
        10'b0011111001: data <= 17'h1ffd9; 
        10'b0011111010: data <= 17'h1ffe4; 
        10'b0011111011: data <= 17'h00021; 
        10'b0011111100: data <= 17'h00002; 
        10'b0011111101: data <= 17'h00007; 
        10'b0011111110: data <= 17'h1ffcc; 
        10'b0011111111: data <= 17'h1ffc0; 
        10'b0100000000: data <= 17'h1ffdd; 
        10'b0100000001: data <= 17'h000ca; 
        10'b0100000010: data <= 17'h00096; 
        10'b0100000011: data <= 17'h00134; 
        10'b0100000100: data <= 17'h0019d; 
        10'b0100000101: data <= 17'h0015c; 
        10'b0100000110: data <= 17'h000dd; 
        10'b0100000111: data <= 17'h00184; 
        10'b0100001000: data <= 17'h00069; 
        10'b0100001001: data <= 17'h00070; 
        10'b0100001010: data <= 17'h1fe3a; 
        10'b0100001011: data <= 17'h1fd89; 
        10'b0100001100: data <= 17'h1ff24; 
        10'b0100001101: data <= 17'h00022; 
        10'b0100001110: data <= 17'h00044; 
        10'b0100001111: data <= 17'h0007b; 
        10'b0100010000: data <= 17'h000a2; 
        10'b0100010001: data <= 17'h0008c; 
        10'b0100010010: data <= 17'h0014d; 
        10'b0100010011: data <= 17'h00156; 
        10'b0100010100: data <= 17'h1ffc8; 
        10'b0100010101: data <= 17'h1ffd1; 
        10'b0100010110: data <= 17'h0004c; 
        10'b0100010111: data <= 17'h1ff97; 
        10'b0100011000: data <= 17'h1ffad; 
        10'b0100011001: data <= 17'h00003; 
        10'b0100011010: data <= 17'h1ffa8; 
        10'b0100011011: data <= 17'h00009; 
        10'b0100011100: data <= 17'h0004e; 
        10'b0100011101: data <= 17'h000f8; 
        10'b0100011110: data <= 17'h000f6; 
        10'b0100011111: data <= 17'h001c3; 
        10'b0100100000: data <= 17'h0014f; 
        10'b0100100001: data <= 17'h00187; 
        10'b0100100010: data <= 17'h0023c; 
        10'b0100100011: data <= 17'h00112; 
        10'b0100100100: data <= 17'h0011e; 
        10'b0100100101: data <= 17'h000ea; 
        10'b0100100110: data <= 17'h1ffb4; 
        10'b0100100111: data <= 17'h1fda7; 
        10'b0100101000: data <= 17'h1fe14; 
        10'b0100101001: data <= 17'h1ff6a; 
        10'b0100101010: data <= 17'h000ab; 
        10'b0100101011: data <= 17'h000aa; 
        10'b0100101100: data <= 17'h000af; 
        10'b0100101101: data <= 17'h00197; 
        10'b0100101110: data <= 17'h001c2; 
        10'b0100101111: data <= 17'h0016f; 
        10'b0100110000: data <= 17'h00005; 
        10'b0100110001: data <= 17'h1ffe5; 
        10'b0100110010: data <= 17'h1ffd0; 
        10'b0100110011: data <= 17'h1ffb1; 
        10'b0100110100: data <= 17'h1ffa8; 
        10'b0100110101: data <= 17'h00014; 
        10'b0100110110: data <= 17'h1fff8; 
        10'b0100110111: data <= 17'h1ff75; 
        10'b0100111000: data <= 17'h00076; 
        10'b0100111001: data <= 17'h00111; 
        10'b0100111010: data <= 17'h00208; 
        10'b0100111011: data <= 17'h002a4; 
        10'b0100111100: data <= 17'h00213; 
        10'b0100111101: data <= 17'h0029f; 
        10'b0100111110: data <= 17'h001cb; 
        10'b0100111111: data <= 17'h000d9; 
        10'b0101000000: data <= 17'h00118; 
        10'b0101000001: data <= 17'h0029c; 
        10'b0101000010: data <= 17'h0032d; 
        10'b0101000011: data <= 17'h1ff9c; 
        10'b0101000100: data <= 17'h1fe1c; 
        10'b0101000101: data <= 17'h1ff59; 
        10'b0101000110: data <= 17'h1ff61; 
        10'b0101000111: data <= 17'h00043; 
        10'b0101001000: data <= 17'h00170; 
        10'b0101001001: data <= 17'h001b9; 
        10'b0101001010: data <= 17'h0024a; 
        10'b0101001011: data <= 17'h00229; 
        10'b0101001100: data <= 17'h00181; 
        10'b0101001101: data <= 17'h0003e; 
        10'b0101001110: data <= 17'h00022; 
        10'b0101001111: data <= 17'h1ffe0; 
        10'b0101010000: data <= 17'h1ffb3; 
        10'b0101010001: data <= 17'h1ffe6; 
        10'b0101010010: data <= 17'h1ffbf; 
        10'b0101010011: data <= 17'h1ffe2; 
        10'b0101010100: data <= 17'h1ffe7; 
        10'b0101010101: data <= 17'h00147; 
        10'b0101010110: data <= 17'h0010f; 
        10'b0101010111: data <= 17'h0019e; 
        10'b0101011000: data <= 17'h00187; 
        10'b0101011001: data <= 17'h001eb; 
        10'b0101011010: data <= 17'h00054; 
        10'b0101011011: data <= 17'h00075; 
        10'b0101011100: data <= 17'h00041; 
        10'b0101011101: data <= 17'h00327; 
        10'b0101011110: data <= 17'h0032b; 
        10'b0101011111: data <= 17'h000b6; 
        10'b0101100000: data <= 17'h0001f; 
        10'b0101100001: data <= 17'h1ffb9; 
        10'b0101100010: data <= 17'h1ffc6; 
        10'b0101100011: data <= 17'h000cb; 
        10'b0101100100: data <= 17'h00159; 
        10'b0101100101: data <= 17'h00251; 
        10'b0101100110: data <= 17'h002b2; 
        10'b0101100111: data <= 17'h00240; 
        10'b0101101000: data <= 17'h00169; 
        10'b0101101001: data <= 17'h00091; 
        10'b0101101010: data <= 17'h00048; 
        10'b0101101011: data <= 17'h1ff9a; 
        10'b0101101100: data <= 17'h1ff90; 
        10'b0101101101: data <= 17'h1ffd7; 
        10'b0101101110: data <= 17'h00017; 
        10'b0101101111: data <= 17'h1ffa0; 
        10'b0101110000: data <= 17'h1ffb7; 
        10'b0101110001: data <= 17'h1fffe; 
        10'b0101110010: data <= 17'h1ffcc; 
        10'b0101110011: data <= 17'h1ffcf; 
        10'b0101110100: data <= 17'h0002c; 
        10'b0101110101: data <= 17'h1ffc4; 
        10'b0101110110: data <= 17'h1ff4f; 
        10'b0101110111: data <= 17'h00043; 
        10'b0101111000: data <= 17'h00128; 
        10'b0101111001: data <= 17'h002f4; 
        10'b0101111010: data <= 17'h000e2; 
        10'b0101111011: data <= 17'h0022c; 
        10'b0101111100: data <= 17'h000dd; 
        10'b0101111101: data <= 17'h1ff73; 
        10'b0101111110: data <= 17'h0000d; 
        10'b0101111111: data <= 17'h00012; 
        10'b0110000000: data <= 17'h000f6; 
        10'b0110000001: data <= 17'h000df; 
        10'b0110000010: data <= 17'h0007f; 
        10'b0110000011: data <= 17'h000b4; 
        10'b0110000100: data <= 17'h00060; 
        10'b0110000101: data <= 17'h00015; 
        10'b0110000110: data <= 17'h00016; 
        10'b0110000111: data <= 17'h1ffed; 
        10'b0110001000: data <= 17'h1ffbc; 
        10'b0110001001: data <= 17'h1ff8e; 
        10'b0110001010: data <= 17'h1fff0; 
        10'b0110001011: data <= 17'h1ffd0; 
        10'b0110001100: data <= 17'h1ff9b; 
        10'b0110001101: data <= 17'h1ff24; 
        10'b0110001110: data <= 17'h1fe78; 
        10'b0110001111: data <= 17'h1fe0a; 
        10'b0110010000: data <= 17'h1fdaf; 
        10'b0110010001: data <= 17'h1fe25; 
        10'b0110010010: data <= 17'h1ffbe; 
        10'b0110010011: data <= 17'h00130; 
        10'b0110010100: data <= 17'h00124; 
        10'b0110010101: data <= 17'h0026a; 
        10'b0110010110: data <= 17'h001ee; 
        10'b0110010111: data <= 17'h0014e; 
        10'b0110011000: data <= 17'h1ffd7; 
        10'b0110011001: data <= 17'h0002a; 
        10'b0110011010: data <= 17'h1ffa9; 
        10'b0110011011: data <= 17'h1ff37; 
        10'b0110011100: data <= 17'h1feb8; 
        10'b0110011101: data <= 17'h1fedb; 
        10'b0110011110: data <= 17'h1ff04; 
        10'b0110011111: data <= 17'h1fed6; 
        10'b0110100000: data <= 17'h1ff79; 
        10'b0110100001: data <= 17'h1ffec; 
        10'b0110100010: data <= 17'h1ff87; 
        10'b0110100011: data <= 17'h00003; 
        10'b0110100100: data <= 17'h0000a; 
        10'b0110100101: data <= 17'h1ffb7; 
        10'b0110100110: data <= 17'h1ffac; 
        10'b0110100111: data <= 17'h1ffdd; 
        10'b0110101000: data <= 17'h1ff92; 
        10'b0110101001: data <= 17'h1ff26; 
        10'b0110101010: data <= 17'h1fe18; 
        10'b0110101011: data <= 17'h1fdaa; 
        10'b0110101100: data <= 17'h1fdde; 
        10'b0110101101: data <= 17'h1ff7b; 
        10'b0110101110: data <= 17'h00015; 
        10'b0110101111: data <= 17'h0000d; 
        10'b0110110000: data <= 17'h001a6; 
        10'b0110110001: data <= 17'h001f3; 
        10'b0110110010: data <= 17'h001b4; 
        10'b0110110011: data <= 17'h000fc; 
        10'b0110110100: data <= 17'h1ff82; 
        10'b0110110101: data <= 17'h1ff92; 
        10'b0110110110: data <= 17'h1ffb3; 
        10'b0110110111: data <= 17'h1fe46; 
        10'b0110111000: data <= 17'h1fdda; 
        10'b0110111001: data <= 17'h1fe5a; 
        10'b0110111010: data <= 17'h1fef4; 
        10'b0110111011: data <= 17'h1ff01; 
        10'b0110111100: data <= 17'h1ff40; 
        10'b0110111101: data <= 17'h1ffdf; 
        10'b0110111110: data <= 17'h1ff7b; 
        10'b0110111111: data <= 17'h0000b; 
        10'b0111000000: data <= 17'h1ffc5; 
        10'b0111000001: data <= 17'h1ff93; 
        10'b0111000010: data <= 17'h1ffb5; 
        10'b0111000011: data <= 17'h1ffd8; 
        10'b0111000100: data <= 17'h1ff50; 
        10'b0111000101: data <= 17'h1fec4; 
        10'b0111000110: data <= 17'h1fe05; 
        10'b0111000111: data <= 17'h1fed5; 
        10'b0111001000: data <= 17'h000c9; 
        10'b0111001001: data <= 17'h000df; 
        10'b0111001010: data <= 17'h0005b; 
        10'b0111001011: data <= 17'h000cd; 
        10'b0111001100: data <= 17'h00198; 
        10'b0111001101: data <= 17'h00165; 
        10'b0111001110: data <= 17'h00080; 
        10'b0111001111: data <= 17'h000d5; 
        10'b0111010000: data <= 17'h00048; 
        10'b0111010001: data <= 17'h1ff59; 
        10'b0111010010: data <= 17'h1fe9b; 
        10'b0111010011: data <= 17'h1fe02; 
        10'b0111010100: data <= 17'h1fe02; 
        10'b0111010101: data <= 17'h1fdfa; 
        10'b0111010110: data <= 17'h1fe61; 
        10'b0111010111: data <= 17'h1ff76; 
        10'b0111011000: data <= 17'h1ff4a; 
        10'b0111011001: data <= 17'h1ffc2; 
        10'b0111011010: data <= 17'h1ffc0; 
        10'b0111011011: data <= 17'h1ff90; 
        10'b0111011100: data <= 17'h00019; 
        10'b0111011101: data <= 17'h00011; 
        10'b0111011110: data <= 17'h1ffa9; 
        10'b0111011111: data <= 17'h1ff95; 
        10'b0111100000: data <= 17'h1ff8b; 
        10'b0111100001: data <= 17'h1feb9; 
        10'b0111100010: data <= 17'h1fe40; 
        10'b0111100011: data <= 17'h0004f; 
        10'b0111100100: data <= 17'h001a0; 
        10'b0111100101: data <= 17'h00204; 
        10'b0111100110: data <= 17'h000a5; 
        10'b0111100111: data <= 17'h00186; 
        10'b0111101000: data <= 17'h0027b; 
        10'b0111101001: data <= 17'h00181; 
        10'b0111101010: data <= 17'h00021; 
        10'b0111101011: data <= 17'h1ff99; 
        10'b0111101100: data <= 17'h0002e; 
        10'b0111101101: data <= 17'h1ff3a; 
        10'b0111101110: data <= 17'h1fdf4; 
        10'b0111101111: data <= 17'h1ff08; 
        10'b0111110000: data <= 17'h1ff0a; 
        10'b0111110001: data <= 17'h1fea4; 
        10'b0111110010: data <= 17'h1fefe; 
        10'b0111110011: data <= 17'h1ff5e; 
        10'b0111110100: data <= 17'h1ffa4; 
        10'b0111110101: data <= 17'h1ff7c; 
        10'b0111110110: data <= 17'h1ffea; 
        10'b0111110111: data <= 17'h1ffbc; 
        10'b0111111000: data <= 17'h1ffb1; 
        10'b0111111001: data <= 17'h00005; 
        10'b0111111010: data <= 17'h1ff8f; 
        10'b0111111011: data <= 17'h1ff6f; 
        10'b0111111100: data <= 17'h1ff39; 
        10'b0111111101: data <= 17'h1ff34; 
        10'b0111111110: data <= 17'h1ff82; 
        10'b0111111111: data <= 17'h0007b; 
        10'b1000000000: data <= 17'h00156; 
        10'b1000000001: data <= 17'h0026a; 
        10'b1000000010: data <= 17'h001b0; 
        10'b1000000011: data <= 17'h0024d; 
        10'b1000000100: data <= 17'h0017f; 
        10'b1000000101: data <= 17'h000dd; 
        10'b1000000110: data <= 17'h1fef4; 
        10'b1000000111: data <= 17'h1ffbb; 
        10'b1000001000: data <= 17'h1ff69; 
        10'b1000001001: data <= 17'h1fe6e; 
        10'b1000001010: data <= 17'h1ff9f; 
        10'b1000001011: data <= 17'h1ffb4; 
        10'b1000001100: data <= 17'h0001e; 
        10'b1000001101: data <= 17'h1ff23; 
        10'b1000001110: data <= 17'h1ffde; 
        10'b1000001111: data <= 17'h1ff44; 
        10'b1000010000: data <= 17'h1ff00; 
        10'b1000010001: data <= 17'h1ff7d; 
        10'b1000010010: data <= 17'h1ffeb; 
        10'b1000010011: data <= 17'h00010; 
        10'b1000010100: data <= 17'h1ffb2; 
        10'b1000010101: data <= 17'h1ffda; 
        10'b1000010110: data <= 17'h1ffe3; 
        10'b1000010111: data <= 17'h1ff53; 
        10'b1000011000: data <= 17'h1ff23; 
        10'b1000011001: data <= 17'h1ffa7; 
        10'b1000011010: data <= 17'h0003b; 
        10'b1000011011: data <= 17'h000a3; 
        10'b1000011100: data <= 17'h000aa; 
        10'b1000011101: data <= 17'h001a2; 
        10'b1000011110: data <= 17'h000d7; 
        10'b1000011111: data <= 17'h1ffe2; 
        10'b1000100000: data <= 17'h00066; 
        10'b1000100001: data <= 17'h1fee8; 
        10'b1000100010: data <= 17'h1feb8; 
        10'b1000100011: data <= 17'h1ff83; 
        10'b1000100100: data <= 17'h1ff99; 
        10'b1000100101: data <= 17'h1ff7a; 
        10'b1000100110: data <= 17'h00067; 
        10'b1000100111: data <= 17'h0001e; 
        10'b1000101000: data <= 17'h00085; 
        10'b1000101001: data <= 17'h0000b; 
        10'b1000101010: data <= 17'h00056; 
        10'b1000101011: data <= 17'h1ffb7; 
        10'b1000101100: data <= 17'h1ff3d; 
        10'b1000101101: data <= 17'h1ff8b; 
        10'b1000101110: data <= 17'h1ff9d; 
        10'b1000101111: data <= 17'h0000c; 
        10'b1000110000: data <= 17'h1ffa1; 
        10'b1000110001: data <= 17'h1ffeb; 
        10'b1000110010: data <= 17'h1ffa9; 
        10'b1000110011: data <= 17'h1ff81; 
        10'b1000110100: data <= 17'h1ff01; 
        10'b1000110101: data <= 17'h1ffd5; 
        10'b1000110110: data <= 17'h00029; 
        10'b1000110111: data <= 17'h0016a; 
        10'b1000111000: data <= 17'h0006c; 
        10'b1000111001: data <= 17'h1ffd1; 
        10'b1000111010: data <= 17'h1fffe; 
        10'b1000111011: data <= 17'h1fece; 
        10'b1000111100: data <= 17'h00013; 
        10'b1000111101: data <= 17'h1fff8; 
        10'b1000111110: data <= 17'h1fede; 
        10'b1000111111: data <= 17'h1ffcb; 
        10'b1001000000: data <= 17'h1fead; 
        10'b1001000001: data <= 17'h1ff95; 
        10'b1001000010: data <= 17'h0003c; 
        10'b1001000011: data <= 17'h00025; 
        10'b1001000100: data <= 17'h0006b; 
        10'b1001000101: data <= 17'h000b6; 
        10'b1001000110: data <= 17'h000b6; 
        10'b1001000111: data <= 17'h1ffd3; 
        10'b1001001000: data <= 17'h1ff88; 
        10'b1001001001: data <= 17'h1ff63; 
        10'b1001001010: data <= 17'h1ffd1; 
        10'b1001001011: data <= 17'h1ffa4; 
        10'b1001001100: data <= 17'h00008; 
        10'b1001001101: data <= 17'h1ffcd; 
        10'b1001001110: data <= 17'h00012; 
        10'b1001001111: data <= 17'h1ff38; 
        10'b1001010000: data <= 17'h1fed6; 
        10'b1001010001: data <= 17'h1ffe2; 
        10'b1001010010: data <= 17'h0009d; 
        10'b1001010011: data <= 17'h0014f; 
        10'b1001010100: data <= 17'h00046; 
        10'b1001010101: data <= 17'h0008f; 
        10'b1001010110: data <= 17'h1ffe6; 
        10'b1001010111: data <= 17'h1ff23; 
        10'b1001011000: data <= 17'h1ff84; 
        10'b1001011001: data <= 17'h0004c; 
        10'b1001011010: data <= 17'h1fff9; 
        10'b1001011011: data <= 17'h1ffdd; 
        10'b1001011100: data <= 17'h1fefc; 
        10'b1001011101: data <= 17'h1ff93; 
        10'b1001011110: data <= 17'h1ffb8; 
        10'b1001011111: data <= 17'h1fff6; 
        10'b1001100000: data <= 17'h1fffa; 
        10'b1001100001: data <= 17'h0003e; 
        10'b1001100010: data <= 17'h00036; 
        10'b1001100011: data <= 17'h1ffb2; 
        10'b1001100100: data <= 17'h1ffa2; 
        10'b1001100101: data <= 17'h1fffa; 
        10'b1001100110: data <= 17'h1ffec; 
        10'b1001100111: data <= 17'h1ffc4; 
        10'b1001101000: data <= 17'h1ffe2; 
        10'b1001101001: data <= 17'h1ff8e; 
        10'b1001101010: data <= 17'h1ffb7; 
        10'b1001101011: data <= 17'h1ff81; 
        10'b1001101100: data <= 17'h1ff13; 
        10'b1001101101: data <= 17'h1fe9e; 
        10'b1001101110: data <= 17'h0002a; 
        10'b1001101111: data <= 17'h0005f; 
        10'b1001110000: data <= 17'h1ffea; 
        10'b1001110001: data <= 17'h1ff8f; 
        10'b1001110010: data <= 17'h00048; 
        10'b1001110011: data <= 17'h0001a; 
        10'b1001110100: data <= 17'h001a7; 
        10'b1001110101: data <= 17'h001bc; 
        10'b1001110110: data <= 17'h00139; 
        10'b1001110111: data <= 17'h000f5; 
        10'b1001111000: data <= 17'h1ffeb; 
        10'b1001111001: data <= 17'h1ffe9; 
        10'b1001111010: data <= 17'h0006a; 
        10'b1001111011: data <= 17'h1ff7c; 
        10'b1001111100: data <= 17'h1ff72; 
        10'b1001111101: data <= 17'h0003d; 
        10'b1001111110: data <= 17'h1ffe7; 
        10'b1001111111: data <= 17'h1ffa5; 
        10'b1010000000: data <= 17'h1ffe9; 
        10'b1010000001: data <= 17'h1ffe9; 
        10'b1010000010: data <= 17'h1ffe6; 
        10'b1010000011: data <= 17'h1ffa8; 
        10'b1010000100: data <= 17'h1ffa7; 
        10'b1010000101: data <= 17'h1fff5; 
        10'b1010000110: data <= 17'h1ffd8; 
        10'b1010000111: data <= 17'h1ff8f; 
        10'b1010001000: data <= 17'h1ff08; 
        10'b1010001001: data <= 17'h1fdb0; 
        10'b1010001010: data <= 17'h1fe30; 
        10'b1010001011: data <= 17'h1ff16; 
        10'b1010001100: data <= 17'h00051; 
        10'b1010001101: data <= 17'h00050; 
        10'b1010001110: data <= 17'h000ac; 
        10'b1010001111: data <= 17'h000e0; 
        10'b1010010000: data <= 17'h001f5; 
        10'b1010010001: data <= 17'h002d0; 
        10'b1010010010: data <= 17'h00265; 
        10'b1010010011: data <= 17'h001e9; 
        10'b1010010100: data <= 17'h0018c; 
        10'b1010010101: data <= 17'h0011b; 
        10'b1010010110: data <= 17'h000e1; 
        10'b1010010111: data <= 17'h00120; 
        10'b1010011000: data <= 17'h000d4; 
        10'b1010011001: data <= 17'h00033; 
        10'b1010011010: data <= 17'h1ffe5; 
        10'b1010011011: data <= 17'h1ffbd; 
        10'b1010011100: data <= 17'h1ff7d; 
        10'b1010011101: data <= 17'h1fff4; 
        10'b1010011110: data <= 17'h1ff8c; 
        10'b1010011111: data <= 17'h1ffe9; 
        10'b1010100000: data <= 17'h1fff2; 
        10'b1010100001: data <= 17'h1ffe9; 
        10'b1010100010: data <= 17'h00016; 
        10'b1010100011: data <= 17'h1ff9a; 
        10'b1010100100: data <= 17'h1ff99; 
        10'b1010100101: data <= 17'h1fe78; 
        10'b1010100110: data <= 17'h1fde0; 
        10'b1010100111: data <= 17'h1fe37; 
        10'b1010101000: data <= 17'h1ffe4; 
        10'b1010101001: data <= 17'h0006b; 
        10'b1010101010: data <= 17'h1ffd8; 
        10'b1010101011: data <= 17'h000c2; 
        10'b1010101100: data <= 17'h0008f; 
        10'b1010101101: data <= 17'h0005e; 
        10'b1010101110: data <= 17'h000ed; 
        10'b1010101111: data <= 17'h00204; 
        10'b1010110000: data <= 17'h00224; 
        10'b1010110001: data <= 17'h00170; 
        10'b1010110010: data <= 17'h00203; 
        10'b1010110011: data <= 17'h001e4; 
        10'b1010110100: data <= 17'h0009f; 
        10'b1010110101: data <= 17'h00009; 
        10'b1010110110: data <= 17'h1ff93; 
        10'b1010110111: data <= 17'h0000b; 
        10'b1010111000: data <= 17'h1ffd3; 
        10'b1010111001: data <= 17'h1ffb5; 
        10'b1010111010: data <= 17'h00012; 
        10'b1010111011: data <= 17'h1ffe2; 
        10'b1010111100: data <= 17'h00018; 
        10'b1010111101: data <= 17'h1ffef; 
        10'b1010111110: data <= 17'h0000b; 
        10'b1010111111: data <= 17'h1ff99; 
        10'b1011000000: data <= 17'h1ffb2; 
        10'b1011000001: data <= 17'h1ff6e; 
        10'b1011000010: data <= 17'h1ff33; 
        10'b1011000011: data <= 17'h1ff01; 
        10'b1011000100: data <= 17'h1fee3; 
        10'b1011000101: data <= 17'h1fee3; 
        10'b1011000110: data <= 17'h1ff95; 
        10'b1011000111: data <= 17'h1ff36; 
        10'b1011001000: data <= 17'h1ff89; 
        10'b1011001001: data <= 17'h1ff87; 
        10'b1011001010: data <= 17'h1fff4; 
        10'b1011001011: data <= 17'h000b5; 
        10'b1011001100: data <= 17'h00081; 
        10'b1011001101: data <= 17'h000a4; 
        10'b1011001110: data <= 17'h000bb; 
        10'b1011001111: data <= 17'h0001e; 
        10'b1011010000: data <= 17'h1ffd8; 
        10'b1011010001: data <= 17'h1fffb; 
        10'b1011010010: data <= 17'h1ff84; 
        10'b1011010011: data <= 17'h1ff89; 
        10'b1011010100: data <= 17'h1fff6; 
        10'b1011010101: data <= 17'h1ffdf; 
        10'b1011010110: data <= 17'h1ffb3; 
        10'b1011010111: data <= 17'h1ffdc; 
        10'b1011011000: data <= 17'h1ffed; 
        10'b1011011001: data <= 17'h00003; 
        10'b1011011010: data <= 17'h1ffc7; 
        10'b1011011011: data <= 17'h1ffad; 
        10'b1011011100: data <= 17'h1ff87; 
        10'b1011011101: data <= 17'h1ff9a; 
        10'b1011011110: data <= 17'h1ff64; 
        10'b1011011111: data <= 17'h1ffd4; 
        10'b1011100000: data <= 17'h1ff73; 
        10'b1011100001: data <= 17'h1ff88; 
        10'b1011100010: data <= 17'h1ff6f; 
        10'b1011100011: data <= 17'h1ffad; 
        10'b1011100100: data <= 17'h1ffa5; 
        10'b1011100101: data <= 17'h1ffb2; 
        10'b1011100110: data <= 17'h1ff8d; 
        10'b1011100111: data <= 17'h1ffad; 
        10'b1011101000: data <= 17'h1ff9b; 
        10'b1011101001: data <= 17'h1ff7b; 
        10'b1011101010: data <= 17'h1ff6b; 
        10'b1011101011: data <= 17'h1ffa2; 
        10'b1011101100: data <= 17'h1ffbf; 
        10'b1011101101: data <= 17'h1ffec; 
        10'b1011101110: data <= 17'h1ffc5; 
        10'b1011101111: data <= 17'h0001a; 
        10'b1011110000: data <= 17'h00018; 
        10'b1011110001: data <= 17'h1ff90; 
        10'b1011110010: data <= 17'h1ffdd; 
        10'b1011110011: data <= 17'h1ffd1; 
        10'b1011110100: data <= 17'h1ffe7; 
        10'b1011110101: data <= 17'h1ffaa; 
        10'b1011110110: data <= 17'h1ffca; 
        10'b1011110111: data <= 17'h1ffde; 
        10'b1011111000: data <= 17'h1ffe3; 
        10'b1011111001: data <= 17'h1ff8d; 
        10'b1011111010: data <= 17'h1fffc; 
        10'b1011111011: data <= 17'h1ffb3; 
        10'b1011111100: data <= 17'h00013; 
        10'b1011111101: data <= 17'h1ffc7; 
        10'b1011111110: data <= 17'h1ff9d; 
        10'b1011111111: data <= 17'h1fff5; 
        10'b1100000000: data <= 17'h1ffaf; 
        10'b1100000001: data <= 17'h1ff9f; 
        10'b1100000010: data <= 17'h1ffc3; 
        10'b1100000011: data <= 17'h1ffe6; 
        10'b1100000100: data <= 17'h1ffdc; 
        10'b1100000101: data <= 17'h00002; 
        10'b1100000110: data <= 17'h00010; 
        10'b1100000111: data <= 17'h00017; 
        10'b1100001000: data <= 17'h1ffed; 
        10'b1100001001: data <= 17'h1ffdf; 
        10'b1100001010: data <= 17'h1ffeb; 
        10'b1100001011: data <= 17'h1ffa7; 
        10'b1100001100: data <= 17'h1ffd7; 
        10'b1100001101: data <= 17'h00011; 
        10'b1100001110: data <= 17'h1ff96; 
        10'b1100001111: data <= 17'h1ffd8; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 12) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 18'h3ff8d; 
        10'b0000000001: data <= 18'h3ffa4; 
        10'b0000000010: data <= 18'h3ff91; 
        10'b0000000011: data <= 18'h3ffcb; 
        10'b0000000100: data <= 18'h3ffbd; 
        10'b0000000101: data <= 18'h00017; 
        10'b0000000110: data <= 18'h3ff15; 
        10'b0000000111: data <= 18'h3ffce; 
        10'b0000001000: data <= 18'h3ff62; 
        10'b0000001001: data <= 18'h3ff7a; 
        10'b0000001010: data <= 18'h3ff43; 
        10'b0000001011: data <= 18'h00014; 
        10'b0000001100: data <= 18'h3ffb5; 
        10'b0000001101: data <= 18'h3fff3; 
        10'b0000001110: data <= 18'h3ff3c; 
        10'b0000001111: data <= 18'h3fff5; 
        10'b0000010000: data <= 18'h3ffc4; 
        10'b0000010001: data <= 18'h3ff2d; 
        10'b0000010010: data <= 18'h00015; 
        10'b0000010011: data <= 18'h3ffa3; 
        10'b0000010100: data <= 18'h3ff91; 
        10'b0000010101: data <= 18'h3ff8a; 
        10'b0000010110: data <= 18'h3ff9b; 
        10'b0000010111: data <= 18'h0002c; 
        10'b0000011000: data <= 18'h00001; 
        10'b0000011001: data <= 18'h3ff79; 
        10'b0000011010: data <= 18'h3ff58; 
        10'b0000011011: data <= 18'h3ff97; 
        10'b0000011100: data <= 18'h3ff91; 
        10'b0000011101: data <= 18'h3ff16; 
        10'b0000011110: data <= 18'h00027; 
        10'b0000011111: data <= 18'h00000; 
        10'b0000100000: data <= 18'h3ff2b; 
        10'b0000100001: data <= 18'h3ff31; 
        10'b0000100010: data <= 18'h3ff1e; 
        10'b0000100011: data <= 18'h3ff32; 
        10'b0000100100: data <= 18'h0001d; 
        10'b0000100101: data <= 18'h3ffaa; 
        10'b0000100110: data <= 18'h3ffa0; 
        10'b0000100111: data <= 18'h3ff18; 
        10'b0000101000: data <= 18'h0001a; 
        10'b0000101001: data <= 18'h3ffdb; 
        10'b0000101010: data <= 18'h3ff62; 
        10'b0000101011: data <= 18'h3ff88; 
        10'b0000101100: data <= 18'h3ffdc; 
        10'b0000101101: data <= 18'h3ffb5; 
        10'b0000101110: data <= 18'h3ff4c; 
        10'b0000101111: data <= 18'h3ffbb; 
        10'b0000110000: data <= 18'h00016; 
        10'b0000110001: data <= 18'h3ff26; 
        10'b0000110010: data <= 18'h3ffd9; 
        10'b0000110011: data <= 18'h3ff4e; 
        10'b0000110100: data <= 18'h3ffef; 
        10'b0000110101: data <= 18'h00030; 
        10'b0000110110: data <= 18'h3ff62; 
        10'b0000110111: data <= 18'h3ff4c; 
        10'b0000111000: data <= 18'h3ff3d; 
        10'b0000111001: data <= 18'h3fffc; 
        10'b0000111010: data <= 18'h3ffb2; 
        10'b0000111011: data <= 18'h3ff9f; 
        10'b0000111100: data <= 18'h3ff45; 
        10'b0000111101: data <= 18'h3ff1b; 
        10'b0000111110: data <= 18'h3ffb3; 
        10'b0000111111: data <= 18'h3ff14; 
        10'b0001000000: data <= 18'h0002a; 
        10'b0001000001: data <= 18'h3ff13; 
        10'b0001000010: data <= 18'h3ff1e; 
        10'b0001000011: data <= 18'h3ffd2; 
        10'b0001000100: data <= 18'h3ffb1; 
        10'b0001000101: data <= 18'h3ff0e; 
        10'b0001000110: data <= 18'h3ffcf; 
        10'b0001000111: data <= 18'h3ffbf; 
        10'b0001001000: data <= 18'h3feff; 
        10'b0001001001: data <= 18'h3ff69; 
        10'b0001001010: data <= 18'h3ff6a; 
        10'b0001001011: data <= 18'h3ffe0; 
        10'b0001001100: data <= 18'h3fff8; 
        10'b0001001101: data <= 18'h3fff4; 
        10'b0001001110: data <= 18'h3ffc7; 
        10'b0001001111: data <= 18'h3ff98; 
        10'b0001010000: data <= 18'h00016; 
        10'b0001010001: data <= 18'h3ff61; 
        10'b0001010010: data <= 18'h3ffdc; 
        10'b0001010011: data <= 18'h0001e; 
        10'b0001010100: data <= 18'h3ff51; 
        10'b0001010101: data <= 18'h3ff9b; 
        10'b0001010110: data <= 18'h3ff9d; 
        10'b0001010111: data <= 18'h3ff34; 
        10'b0001011000: data <= 18'h00029; 
        10'b0001011001: data <= 18'h3ff40; 
        10'b0001011010: data <= 18'h3ff24; 
        10'b0001011011: data <= 18'h3ff7b; 
        10'b0001011100: data <= 18'h3ff19; 
        10'b0001011101: data <= 18'h3ffb0; 
        10'b0001011110: data <= 18'h3ff53; 
        10'b0001011111: data <= 18'h3febe; 
        10'b0001100000: data <= 18'h3fe9a; 
        10'b0001100001: data <= 18'h3fe4e; 
        10'b0001100010: data <= 18'h3fe98; 
        10'b0001100011: data <= 18'h3ff2b; 
        10'b0001100100: data <= 18'h3fe97; 
        10'b0001100101: data <= 18'h3fee7; 
        10'b0001100110: data <= 18'h3ff3d; 
        10'b0001100111: data <= 18'h3ff88; 
        10'b0001101000: data <= 18'h3feef; 
        10'b0001101001: data <= 18'h00011; 
        10'b0001101010: data <= 18'h3ff71; 
        10'b0001101011: data <= 18'h3fff2; 
        10'b0001101100: data <= 18'h3ff64; 
        10'b0001101101: data <= 18'h3ffce; 
        10'b0001101110: data <= 18'h3ffb7; 
        10'b0001101111: data <= 18'h3ff29; 
        10'b0001110000: data <= 18'h3ffa2; 
        10'b0001110001: data <= 18'h3ffe5; 
        10'b0001110010: data <= 18'h3ff79; 
        10'b0001110011: data <= 18'h3ff2a; 
        10'b0001110100: data <= 18'h3fff4; 
        10'b0001110101: data <= 18'h3fff0; 
        10'b0001110110: data <= 18'h3ffa3; 
        10'b0001110111: data <= 18'h3ff3e; 
        10'b0001111000: data <= 18'h3ff3d; 
        10'b0001111001: data <= 18'h3ff8d; 
        10'b0001111010: data <= 18'h3ff9b; 
        10'b0001111011: data <= 18'h3ffc8; 
        10'b0001111100: data <= 18'h00137; 
        10'b0001111101: data <= 18'h000c9; 
        10'b0001111110: data <= 18'h002a6; 
        10'b0001111111: data <= 18'h00203; 
        10'b0010000000: data <= 18'h000ea; 
        10'b0010000001: data <= 18'h00080; 
        10'b0010000010: data <= 18'h000c0; 
        10'b0010000011: data <= 18'h3ff55; 
        10'b0010000100: data <= 18'h3ff30; 
        10'b0010000101: data <= 18'h3ff94; 
        10'b0010000110: data <= 18'h3fec6; 
        10'b0010000111: data <= 18'h3ff1f; 
        10'b0010001000: data <= 18'h3fff9; 
        10'b0010001001: data <= 18'h0000f; 
        10'b0010001010: data <= 18'h3ff87; 
        10'b0010001011: data <= 18'h3ffa3; 
        10'b0010001100: data <= 18'h3ffa7; 
        10'b0010001101: data <= 18'h3ffd6; 
        10'b0010001110: data <= 18'h3ffe5; 
        10'b0010001111: data <= 18'h3fff8; 
        10'b0010010000: data <= 18'h3ff47; 
        10'b0010010001: data <= 18'h3ff93; 
        10'b0010010010: data <= 18'h3ff61; 
        10'b0010010011: data <= 18'h3fe51; 
        10'b0010010100: data <= 18'h3ff53; 
        10'b0010010101: data <= 18'h0009a; 
        10'b0010010110: data <= 18'h3fe9c; 
        10'b0010010111: data <= 18'h001da; 
        10'b0010011000: data <= 18'h0037b; 
        10'b0010011001: data <= 18'h002e5; 
        10'b0010011010: data <= 18'h00303; 
        10'b0010011011: data <= 18'h00170; 
        10'b0010011100: data <= 18'h00130; 
        10'b0010011101: data <= 18'h002ca; 
        10'b0010011110: data <= 18'h00024; 
        10'b0010011111: data <= 18'h3ffdf; 
        10'b0010100000: data <= 18'h000ff; 
        10'b0010100001: data <= 18'h00084; 
        10'b0010100010: data <= 18'h3fe50; 
        10'b0010100011: data <= 18'h3fe95; 
        10'b0010100100: data <= 18'h3ff05; 
        10'b0010100101: data <= 18'h000bf; 
        10'b0010100110: data <= 18'h3ffb2; 
        10'b0010100111: data <= 18'h00021; 
        10'b0010101000: data <= 18'h3ff50; 
        10'b0010101001: data <= 18'h3ff42; 
        10'b0010101010: data <= 18'h3ff19; 
        10'b0010101011: data <= 18'h3ff1e; 
        10'b0010101100: data <= 18'h3fefd; 
        10'b0010101101: data <= 18'h3ff03; 
        10'b0010101110: data <= 18'h3fe69; 
        10'b0010101111: data <= 18'h3fe68; 
        10'b0010110000: data <= 18'h0001c; 
        10'b0010110001: data <= 18'h00078; 
        10'b0010110010: data <= 18'h3ffe0; 
        10'b0010110011: data <= 18'h000e5; 
        10'b0010110100: data <= 18'h0016b; 
        10'b0010110101: data <= 18'h00123; 
        10'b0010110110: data <= 18'h0019a; 
        10'b0010110111: data <= 18'h002ff; 
        10'b0010111000: data <= 18'h00173; 
        10'b0010111001: data <= 18'h001b5; 
        10'b0010111010: data <= 18'h0005c; 
        10'b0010111011: data <= 18'h001f2; 
        10'b0010111100: data <= 18'h000be; 
        10'b0010111101: data <= 18'h000ea; 
        10'b0010111110: data <= 18'h00123; 
        10'b0010111111: data <= 18'h00110; 
        10'b0011000000: data <= 18'h000e5; 
        10'b0011000001: data <= 18'h00060; 
        10'b0011000010: data <= 18'h3ffa2; 
        10'b0011000011: data <= 18'h3ffe9; 
        10'b0011000100: data <= 18'h00022; 
        10'b0011000101: data <= 18'h3ff52; 
        10'b0011000110: data <= 18'h3ff34; 
        10'b0011000111: data <= 18'h3ff61; 
        10'b0011001000: data <= 18'h3fef2; 
        10'b0011001001: data <= 18'h3ff9e; 
        10'b0011001010: data <= 18'h3feea; 
        10'b0011001011: data <= 18'h3fff0; 
        10'b0011001100: data <= 18'h00112; 
        10'b0011001101: data <= 18'h00070; 
        10'b0011001110: data <= 18'h0008a; 
        10'b0011001111: data <= 18'h3ffaa; 
        10'b0011010000: data <= 18'h3fea1; 
        10'b0011010001: data <= 18'h3fef9; 
        10'b0011010010: data <= 18'h3fe7d; 
        10'b0011010011: data <= 18'h000e8; 
        10'b0011010100: data <= 18'h00123; 
        10'b0011010101: data <= 18'h3ffee; 
        10'b0011010110: data <= 18'h000c7; 
        10'b0011010111: data <= 18'h3ff27; 
        10'b0011011000: data <= 18'h00129; 
        10'b0011011001: data <= 18'h001cf; 
        10'b0011011010: data <= 18'h00053; 
        10'b0011011011: data <= 18'h003c1; 
        10'b0011011100: data <= 18'h0024c; 
        10'b0011011101: data <= 18'h3ffea; 
        10'b0011011110: data <= 18'h0000e; 
        10'b0011011111: data <= 18'h3ffd8; 
        10'b0011100000: data <= 18'h3ffd7; 
        10'b0011100001: data <= 18'h0000d; 
        10'b0011100010: data <= 18'h3ffd1; 
        10'b0011100011: data <= 18'h3ff42; 
        10'b0011100100: data <= 18'h3ffce; 
        10'b0011100101: data <= 18'h3ffa7; 
        10'b0011100110: data <= 18'h0018e; 
        10'b0011100111: data <= 18'h000f6; 
        10'b0011101000: data <= 18'h00059; 
        10'b0011101001: data <= 18'h002b2; 
        10'b0011101010: data <= 18'h00027; 
        10'b0011101011: data <= 18'h00017; 
        10'b0011101100: data <= 18'h001cd; 
        10'b0011101101: data <= 18'h00255; 
        10'b0011101110: data <= 18'h3fe28; 
        10'b0011101111: data <= 18'h3fe6f; 
        10'b0011110000: data <= 18'h00147; 
        10'b0011110001: data <= 18'h3ff19; 
        10'b0011110010: data <= 18'h0006d; 
        10'b0011110011: data <= 18'h00139; 
        10'b0011110100: data <= 18'h000ce; 
        10'b0011110101: data <= 18'h0027d; 
        10'b0011110110: data <= 18'h001ab; 
        10'b0011110111: data <= 18'h002d6; 
        10'b0011111000: data <= 18'h00294; 
        10'b0011111001: data <= 18'h3ffb1; 
        10'b0011111010: data <= 18'h3ffc8; 
        10'b0011111011: data <= 18'h00041; 
        10'b0011111100: data <= 18'h00004; 
        10'b0011111101: data <= 18'h0000d; 
        10'b0011111110: data <= 18'h3ff99; 
        10'b0011111111: data <= 18'h3ff80; 
        10'b0100000000: data <= 18'h3ffba; 
        10'b0100000001: data <= 18'h00193; 
        10'b0100000010: data <= 18'h0012b; 
        10'b0100000011: data <= 18'h00268; 
        10'b0100000100: data <= 18'h0033b; 
        10'b0100000101: data <= 18'h002b9; 
        10'b0100000110: data <= 18'h001ba; 
        10'b0100000111: data <= 18'h00308; 
        10'b0100001000: data <= 18'h000d2; 
        10'b0100001001: data <= 18'h000e1; 
        10'b0100001010: data <= 18'h3fc74; 
        10'b0100001011: data <= 18'h3fb11; 
        10'b0100001100: data <= 18'h3fe48; 
        10'b0100001101: data <= 18'h00043; 
        10'b0100001110: data <= 18'h00089; 
        10'b0100001111: data <= 18'h000f5; 
        10'b0100010000: data <= 18'h00144; 
        10'b0100010001: data <= 18'h00117; 
        10'b0100010010: data <= 18'h0029b; 
        10'b0100010011: data <= 18'h002ad; 
        10'b0100010100: data <= 18'h3ff91; 
        10'b0100010101: data <= 18'h3ffa2; 
        10'b0100010110: data <= 18'h00098; 
        10'b0100010111: data <= 18'h3ff2f; 
        10'b0100011000: data <= 18'h3ff5a; 
        10'b0100011001: data <= 18'h00007; 
        10'b0100011010: data <= 18'h3ff4f; 
        10'b0100011011: data <= 18'h00012; 
        10'b0100011100: data <= 18'h0009b; 
        10'b0100011101: data <= 18'h001ef; 
        10'b0100011110: data <= 18'h001ec; 
        10'b0100011111: data <= 18'h00386; 
        10'b0100100000: data <= 18'h0029e; 
        10'b0100100001: data <= 18'h0030f; 
        10'b0100100010: data <= 18'h00477; 
        10'b0100100011: data <= 18'h00224; 
        10'b0100100100: data <= 18'h0023d; 
        10'b0100100101: data <= 18'h001d3; 
        10'b0100100110: data <= 18'h3ff68; 
        10'b0100100111: data <= 18'h3fb4e; 
        10'b0100101000: data <= 18'h3fc27; 
        10'b0100101001: data <= 18'h3fed4; 
        10'b0100101010: data <= 18'h00157; 
        10'b0100101011: data <= 18'h00155; 
        10'b0100101100: data <= 18'h0015e; 
        10'b0100101101: data <= 18'h0032d; 
        10'b0100101110: data <= 18'h00384; 
        10'b0100101111: data <= 18'h002de; 
        10'b0100110000: data <= 18'h00009; 
        10'b0100110001: data <= 18'h3ffca; 
        10'b0100110010: data <= 18'h3ffa1; 
        10'b0100110011: data <= 18'h3ff62; 
        10'b0100110100: data <= 18'h3ff4f; 
        10'b0100110101: data <= 18'h00028; 
        10'b0100110110: data <= 18'h3fff0; 
        10'b0100110111: data <= 18'h3fee9; 
        10'b0100111000: data <= 18'h000ec; 
        10'b0100111001: data <= 18'h00223; 
        10'b0100111010: data <= 18'h00411; 
        10'b0100111011: data <= 18'h00547; 
        10'b0100111100: data <= 18'h00426; 
        10'b0100111101: data <= 18'h0053e; 
        10'b0100111110: data <= 18'h00397; 
        10'b0100111111: data <= 18'h001b2; 
        10'b0101000000: data <= 18'h00230; 
        10'b0101000001: data <= 18'h00538; 
        10'b0101000010: data <= 18'h0065b; 
        10'b0101000011: data <= 18'h3ff38; 
        10'b0101000100: data <= 18'h3fc38; 
        10'b0101000101: data <= 18'h3feb3; 
        10'b0101000110: data <= 18'h3fec3; 
        10'b0101000111: data <= 18'h00085; 
        10'b0101001000: data <= 18'h002e0; 
        10'b0101001001: data <= 18'h00372; 
        10'b0101001010: data <= 18'h00493; 
        10'b0101001011: data <= 18'h00451; 
        10'b0101001100: data <= 18'h00301; 
        10'b0101001101: data <= 18'h0007d; 
        10'b0101001110: data <= 18'h00044; 
        10'b0101001111: data <= 18'h3ffc1; 
        10'b0101010000: data <= 18'h3ff66; 
        10'b0101010001: data <= 18'h3ffcc; 
        10'b0101010010: data <= 18'h3ff7e; 
        10'b0101010011: data <= 18'h3ffc4; 
        10'b0101010100: data <= 18'h3ffce; 
        10'b0101010101: data <= 18'h0028e; 
        10'b0101010110: data <= 18'h0021e; 
        10'b0101010111: data <= 18'h0033c; 
        10'b0101011000: data <= 18'h0030d; 
        10'b0101011001: data <= 18'h003d5; 
        10'b0101011010: data <= 18'h000a7; 
        10'b0101011011: data <= 18'h000ea; 
        10'b0101011100: data <= 18'h00082; 
        10'b0101011101: data <= 18'h0064d; 
        10'b0101011110: data <= 18'h00655; 
        10'b0101011111: data <= 18'h0016b; 
        10'b0101100000: data <= 18'h0003e; 
        10'b0101100001: data <= 18'h3ff72; 
        10'b0101100010: data <= 18'h3ff8b; 
        10'b0101100011: data <= 18'h00196; 
        10'b0101100100: data <= 18'h002b2; 
        10'b0101100101: data <= 18'h004a2; 
        10'b0101100110: data <= 18'h00565; 
        10'b0101100111: data <= 18'h00480; 
        10'b0101101000: data <= 18'h002d3; 
        10'b0101101001: data <= 18'h00121; 
        10'b0101101010: data <= 18'h0008f; 
        10'b0101101011: data <= 18'h3ff34; 
        10'b0101101100: data <= 18'h3ff1f; 
        10'b0101101101: data <= 18'h3ffaf; 
        10'b0101101110: data <= 18'h0002e; 
        10'b0101101111: data <= 18'h3ff3f; 
        10'b0101110000: data <= 18'h3ff6e; 
        10'b0101110001: data <= 18'h3fffd; 
        10'b0101110010: data <= 18'h3ff97; 
        10'b0101110011: data <= 18'h3ff9d; 
        10'b0101110100: data <= 18'h00059; 
        10'b0101110101: data <= 18'h3ff89; 
        10'b0101110110: data <= 18'h3fe9e; 
        10'b0101110111: data <= 18'h00087; 
        10'b0101111000: data <= 18'h00251; 
        10'b0101111001: data <= 18'h005e7; 
        10'b0101111010: data <= 18'h001c4; 
        10'b0101111011: data <= 18'h00458; 
        10'b0101111100: data <= 18'h001ba; 
        10'b0101111101: data <= 18'h3fee7; 
        10'b0101111110: data <= 18'h0001a; 
        10'b0101111111: data <= 18'h00025; 
        10'b0110000000: data <= 18'h001ec; 
        10'b0110000001: data <= 18'h001bf; 
        10'b0110000010: data <= 18'h000fd; 
        10'b0110000011: data <= 18'h00168; 
        10'b0110000100: data <= 18'h000c0; 
        10'b0110000101: data <= 18'h0002b; 
        10'b0110000110: data <= 18'h0002c; 
        10'b0110000111: data <= 18'h3ffdb; 
        10'b0110001000: data <= 18'h3ff77; 
        10'b0110001001: data <= 18'h3ff1c; 
        10'b0110001010: data <= 18'h3ffe1; 
        10'b0110001011: data <= 18'h3ffa1; 
        10'b0110001100: data <= 18'h3ff36; 
        10'b0110001101: data <= 18'h3fe49; 
        10'b0110001110: data <= 18'h3fcf0; 
        10'b0110001111: data <= 18'h3fc13; 
        10'b0110010000: data <= 18'h3fb5e; 
        10'b0110010001: data <= 18'h3fc4a; 
        10'b0110010010: data <= 18'h3ff7b; 
        10'b0110010011: data <= 18'h00260; 
        10'b0110010100: data <= 18'h00249; 
        10'b0110010101: data <= 18'h004d3; 
        10'b0110010110: data <= 18'h003dc; 
        10'b0110010111: data <= 18'h0029c; 
        10'b0110011000: data <= 18'h3ffaf; 
        10'b0110011001: data <= 18'h00053; 
        10'b0110011010: data <= 18'h3ff52; 
        10'b0110011011: data <= 18'h3fe6d; 
        10'b0110011100: data <= 18'h3fd70; 
        10'b0110011101: data <= 18'h3fdb5; 
        10'b0110011110: data <= 18'h3fe07; 
        10'b0110011111: data <= 18'h3fdac; 
        10'b0110100000: data <= 18'h3fef2; 
        10'b0110100001: data <= 18'h3ffd9; 
        10'b0110100010: data <= 18'h3ff0f; 
        10'b0110100011: data <= 18'h00007; 
        10'b0110100100: data <= 18'h00013; 
        10'b0110100101: data <= 18'h3ff6e; 
        10'b0110100110: data <= 18'h3ff58; 
        10'b0110100111: data <= 18'h3ffba; 
        10'b0110101000: data <= 18'h3ff23; 
        10'b0110101001: data <= 18'h3fe4c; 
        10'b0110101010: data <= 18'h3fc2f; 
        10'b0110101011: data <= 18'h3fb53; 
        10'b0110101100: data <= 18'h3fbbd; 
        10'b0110101101: data <= 18'h3fef6; 
        10'b0110101110: data <= 18'h00029; 
        10'b0110101111: data <= 18'h0001b; 
        10'b0110110000: data <= 18'h0034c; 
        10'b0110110001: data <= 18'h003e6; 
        10'b0110110010: data <= 18'h00369; 
        10'b0110110011: data <= 18'h001f7; 
        10'b0110110100: data <= 18'h3ff04; 
        10'b0110110101: data <= 18'h3ff24; 
        10'b0110110110: data <= 18'h3ff66; 
        10'b0110110111: data <= 18'h3fc8c; 
        10'b0110111000: data <= 18'h3fbb3; 
        10'b0110111001: data <= 18'h3fcb4; 
        10'b0110111010: data <= 18'h3fde9; 
        10'b0110111011: data <= 18'h3fe02; 
        10'b0110111100: data <= 18'h3fe7f; 
        10'b0110111101: data <= 18'h3ffbd; 
        10'b0110111110: data <= 18'h3fef6; 
        10'b0110111111: data <= 18'h00016; 
        10'b0111000000: data <= 18'h3ff8a; 
        10'b0111000001: data <= 18'h3ff26; 
        10'b0111000010: data <= 18'h3ff69; 
        10'b0111000011: data <= 18'h3ffb1; 
        10'b0111000100: data <= 18'h3fe9f; 
        10'b0111000101: data <= 18'h3fd89; 
        10'b0111000110: data <= 18'h3fc0a; 
        10'b0111000111: data <= 18'h3fda9; 
        10'b0111001000: data <= 18'h00192; 
        10'b0111001001: data <= 18'h001bf; 
        10'b0111001010: data <= 18'h000b7; 
        10'b0111001011: data <= 18'h0019a; 
        10'b0111001100: data <= 18'h00330; 
        10'b0111001101: data <= 18'h002cb; 
        10'b0111001110: data <= 18'h00100; 
        10'b0111001111: data <= 18'h001ab; 
        10'b0111010000: data <= 18'h00091; 
        10'b0111010001: data <= 18'h3feb2; 
        10'b0111010010: data <= 18'h3fd37; 
        10'b0111010011: data <= 18'h3fc05; 
        10'b0111010100: data <= 18'h3fc05; 
        10'b0111010101: data <= 18'h3fbf4; 
        10'b0111010110: data <= 18'h3fcc1; 
        10'b0111010111: data <= 18'h3feec; 
        10'b0111011000: data <= 18'h3fe95; 
        10'b0111011001: data <= 18'h3ff84; 
        10'b0111011010: data <= 18'h3ff7f; 
        10'b0111011011: data <= 18'h3ff20; 
        10'b0111011100: data <= 18'h00032; 
        10'b0111011101: data <= 18'h00023; 
        10'b0111011110: data <= 18'h3ff51; 
        10'b0111011111: data <= 18'h3ff2a; 
        10'b0111100000: data <= 18'h3ff16; 
        10'b0111100001: data <= 18'h3fd73; 
        10'b0111100010: data <= 18'h3fc80; 
        10'b0111100011: data <= 18'h0009e; 
        10'b0111100100: data <= 18'h00341; 
        10'b0111100101: data <= 18'h00408; 
        10'b0111100110: data <= 18'h0014a; 
        10'b0111100111: data <= 18'h0030d; 
        10'b0111101000: data <= 18'h004f6; 
        10'b0111101001: data <= 18'h00303; 
        10'b0111101010: data <= 18'h00041; 
        10'b0111101011: data <= 18'h3ff32; 
        10'b0111101100: data <= 18'h0005c; 
        10'b0111101101: data <= 18'h3fe74; 
        10'b0111101110: data <= 18'h3fbe9; 
        10'b0111101111: data <= 18'h3fe10; 
        10'b0111110000: data <= 18'h3fe14; 
        10'b0111110001: data <= 18'h3fd48; 
        10'b0111110010: data <= 18'h3fdfd; 
        10'b0111110011: data <= 18'h3febb; 
        10'b0111110100: data <= 18'h3ff47; 
        10'b0111110101: data <= 18'h3fef8; 
        10'b0111110110: data <= 18'h3ffd4; 
        10'b0111110111: data <= 18'h3ff77; 
        10'b0111111000: data <= 18'h3ff61; 
        10'b0111111001: data <= 18'h0000a; 
        10'b0111111010: data <= 18'h3ff1d; 
        10'b0111111011: data <= 18'h3fede; 
        10'b0111111100: data <= 18'h3fe72; 
        10'b0111111101: data <= 18'h3fe68; 
        10'b0111111110: data <= 18'h3ff04; 
        10'b0111111111: data <= 18'h000f6; 
        10'b1000000000: data <= 18'h002ad; 
        10'b1000000001: data <= 18'h004d3; 
        10'b1000000010: data <= 18'h0035f; 
        10'b1000000011: data <= 18'h0049a; 
        10'b1000000100: data <= 18'h002ff; 
        10'b1000000101: data <= 18'h001ba; 
        10'b1000000110: data <= 18'h3fde9; 
        10'b1000000111: data <= 18'h3ff76; 
        10'b1000001000: data <= 18'h3fed2; 
        10'b1000001001: data <= 18'h3fcdc; 
        10'b1000001010: data <= 18'h3ff3e; 
        10'b1000001011: data <= 18'h3ff69; 
        10'b1000001100: data <= 18'h0003b; 
        10'b1000001101: data <= 18'h3fe45; 
        10'b1000001110: data <= 18'h3ffbd; 
        10'b1000001111: data <= 18'h3fe88; 
        10'b1000010000: data <= 18'h3fe01; 
        10'b1000010001: data <= 18'h3fef9; 
        10'b1000010010: data <= 18'h3ffd6; 
        10'b1000010011: data <= 18'h00020; 
        10'b1000010100: data <= 18'h3ff65; 
        10'b1000010101: data <= 18'h3ffb3; 
        10'b1000010110: data <= 18'h3ffc6; 
        10'b1000010111: data <= 18'h3fea6; 
        10'b1000011000: data <= 18'h3fe46; 
        10'b1000011001: data <= 18'h3ff4e; 
        10'b1000011010: data <= 18'h00076; 
        10'b1000011011: data <= 18'h00146; 
        10'b1000011100: data <= 18'h00154; 
        10'b1000011101: data <= 18'h00345; 
        10'b1000011110: data <= 18'h001ae; 
        10'b1000011111: data <= 18'h3ffc5; 
        10'b1000100000: data <= 18'h000cc; 
        10'b1000100001: data <= 18'h3fdd0; 
        10'b1000100010: data <= 18'h3fd70; 
        10'b1000100011: data <= 18'h3ff05; 
        10'b1000100100: data <= 18'h3ff32; 
        10'b1000100101: data <= 18'h3fef3; 
        10'b1000100110: data <= 18'h000ce; 
        10'b1000100111: data <= 18'h0003b; 
        10'b1000101000: data <= 18'h00109; 
        10'b1000101001: data <= 18'h00016; 
        10'b1000101010: data <= 18'h000ac; 
        10'b1000101011: data <= 18'h3ff6d; 
        10'b1000101100: data <= 18'h3fe7a; 
        10'b1000101101: data <= 18'h3ff17; 
        10'b1000101110: data <= 18'h3ff3a; 
        10'b1000101111: data <= 18'h00018; 
        10'b1000110000: data <= 18'h3ff42; 
        10'b1000110001: data <= 18'h3ffd7; 
        10'b1000110010: data <= 18'h3ff52; 
        10'b1000110011: data <= 18'h3ff02; 
        10'b1000110100: data <= 18'h3fe02; 
        10'b1000110101: data <= 18'h3ffaa; 
        10'b1000110110: data <= 18'h00051; 
        10'b1000110111: data <= 18'h002d4; 
        10'b1000111000: data <= 18'h000d8; 
        10'b1000111001: data <= 18'h3ffa3; 
        10'b1000111010: data <= 18'h3fffc; 
        10'b1000111011: data <= 18'h3fd9c; 
        10'b1000111100: data <= 18'h00027; 
        10'b1000111101: data <= 18'h3fff0; 
        10'b1000111110: data <= 18'h3fdbb; 
        10'b1000111111: data <= 18'h3ff96; 
        10'b1001000000: data <= 18'h3fd59; 
        10'b1001000001: data <= 18'h3ff29; 
        10'b1001000010: data <= 18'h00078; 
        10'b1001000011: data <= 18'h0004a; 
        10'b1001000100: data <= 18'h000d7; 
        10'b1001000101: data <= 18'h0016d; 
        10'b1001000110: data <= 18'h0016c; 
        10'b1001000111: data <= 18'h3ffa6; 
        10'b1001001000: data <= 18'h3ff11; 
        10'b1001001001: data <= 18'h3fec6; 
        10'b1001001010: data <= 18'h3ffa3; 
        10'b1001001011: data <= 18'h3ff48; 
        10'b1001001100: data <= 18'h00011; 
        10'b1001001101: data <= 18'h3ff9a; 
        10'b1001001110: data <= 18'h00024; 
        10'b1001001111: data <= 18'h3fe6f; 
        10'b1001010000: data <= 18'h3fdad; 
        10'b1001010001: data <= 18'h3ffc5; 
        10'b1001010010: data <= 18'h0013a; 
        10'b1001010011: data <= 18'h0029e; 
        10'b1001010100: data <= 18'h0008c; 
        10'b1001010101: data <= 18'h0011f; 
        10'b1001010110: data <= 18'h3ffcb; 
        10'b1001010111: data <= 18'h3fe46; 
        10'b1001011000: data <= 18'h3ff08; 
        10'b1001011001: data <= 18'h00099; 
        10'b1001011010: data <= 18'h3fff2; 
        10'b1001011011: data <= 18'h3ffba; 
        10'b1001011100: data <= 18'h3fdf8; 
        10'b1001011101: data <= 18'h3ff26; 
        10'b1001011110: data <= 18'h3ff6f; 
        10'b1001011111: data <= 18'h3ffeb; 
        10'b1001100000: data <= 18'h3fff4; 
        10'b1001100001: data <= 18'h0007d; 
        10'b1001100010: data <= 18'h0006c; 
        10'b1001100011: data <= 18'h3ff64; 
        10'b1001100100: data <= 18'h3ff44; 
        10'b1001100101: data <= 18'h3fff4; 
        10'b1001100110: data <= 18'h3ffd9; 
        10'b1001100111: data <= 18'h3ff87; 
        10'b1001101000: data <= 18'h3ffc3; 
        10'b1001101001: data <= 18'h3ff1c; 
        10'b1001101010: data <= 18'h3ff6f; 
        10'b1001101011: data <= 18'h3ff01; 
        10'b1001101100: data <= 18'h3fe25; 
        10'b1001101101: data <= 18'h3fd3c; 
        10'b1001101110: data <= 18'h00054; 
        10'b1001101111: data <= 18'h000bf; 
        10'b1001110000: data <= 18'h3ffd4; 
        10'b1001110001: data <= 18'h3ff1e; 
        10'b1001110010: data <= 18'h0008f; 
        10'b1001110011: data <= 18'h00033; 
        10'b1001110100: data <= 18'h0034e; 
        10'b1001110101: data <= 18'h00377; 
        10'b1001110110: data <= 18'h00273; 
        10'b1001110111: data <= 18'h001ea; 
        10'b1001111000: data <= 18'h3ffd6; 
        10'b1001111001: data <= 18'h3ffd2; 
        10'b1001111010: data <= 18'h000d4; 
        10'b1001111011: data <= 18'h3fef8; 
        10'b1001111100: data <= 18'h3fee3; 
        10'b1001111101: data <= 18'h00079; 
        10'b1001111110: data <= 18'h3ffcd; 
        10'b1001111111: data <= 18'h3ff4a; 
        10'b1010000000: data <= 18'h3ffd3; 
        10'b1010000001: data <= 18'h3ffd1; 
        10'b1010000010: data <= 18'h3ffcb; 
        10'b1010000011: data <= 18'h3ff50; 
        10'b1010000100: data <= 18'h3ff4e; 
        10'b1010000101: data <= 18'h3ffea; 
        10'b1010000110: data <= 18'h3ffb0; 
        10'b1010000111: data <= 18'h3ff1d; 
        10'b1010001000: data <= 18'h3fe0f; 
        10'b1010001001: data <= 18'h3fb5f; 
        10'b1010001010: data <= 18'h3fc5f; 
        10'b1010001011: data <= 18'h3fe2c; 
        10'b1010001100: data <= 18'h000a2; 
        10'b1010001101: data <= 18'h000a0; 
        10'b1010001110: data <= 18'h00158; 
        10'b1010001111: data <= 18'h001c1; 
        10'b1010010000: data <= 18'h003ea; 
        10'b1010010001: data <= 18'h005a0; 
        10'b1010010010: data <= 18'h004ca; 
        10'b1010010011: data <= 18'h003d1; 
        10'b1010010100: data <= 18'h00317; 
        10'b1010010101: data <= 18'h00237; 
        10'b1010010110: data <= 18'h001c2; 
        10'b1010010111: data <= 18'h0023f; 
        10'b1010011000: data <= 18'h001a8; 
        10'b1010011001: data <= 18'h00066; 
        10'b1010011010: data <= 18'h3ffca; 
        10'b1010011011: data <= 18'h3ff7a; 
        10'b1010011100: data <= 18'h3fefa; 
        10'b1010011101: data <= 18'h3ffe7; 
        10'b1010011110: data <= 18'h3ff18; 
        10'b1010011111: data <= 18'h3ffd2; 
        10'b1010100000: data <= 18'h3ffe4; 
        10'b1010100001: data <= 18'h3ffd2; 
        10'b1010100010: data <= 18'h0002c; 
        10'b1010100011: data <= 18'h3ff34; 
        10'b1010100100: data <= 18'h3ff32; 
        10'b1010100101: data <= 18'h3fcf0; 
        10'b1010100110: data <= 18'h3fbc0; 
        10'b1010100111: data <= 18'h3fc6f; 
        10'b1010101000: data <= 18'h3ffc8; 
        10'b1010101001: data <= 18'h000d5; 
        10'b1010101010: data <= 18'h3ffaf; 
        10'b1010101011: data <= 18'h00184; 
        10'b1010101100: data <= 18'h0011e; 
        10'b1010101101: data <= 18'h000bd; 
        10'b1010101110: data <= 18'h001db; 
        10'b1010101111: data <= 18'h00408; 
        10'b1010110000: data <= 18'h00448; 
        10'b1010110001: data <= 18'h002e0; 
        10'b1010110010: data <= 18'h00406; 
        10'b1010110011: data <= 18'h003c7; 
        10'b1010110100: data <= 18'h0013f; 
        10'b1010110101: data <= 18'h00012; 
        10'b1010110110: data <= 18'h3ff25; 
        10'b1010110111: data <= 18'h00016; 
        10'b1010111000: data <= 18'h3ffa6; 
        10'b1010111001: data <= 18'h3ff6a; 
        10'b1010111010: data <= 18'h00023; 
        10'b1010111011: data <= 18'h3ffc4; 
        10'b1010111100: data <= 18'h00030; 
        10'b1010111101: data <= 18'h3ffdd; 
        10'b1010111110: data <= 18'h00017; 
        10'b1010111111: data <= 18'h3ff32; 
        10'b1011000000: data <= 18'h3ff65; 
        10'b1011000001: data <= 18'h3fedd; 
        10'b1011000010: data <= 18'h3fe66; 
        10'b1011000011: data <= 18'h3fe02; 
        10'b1011000100: data <= 18'h3fdc7; 
        10'b1011000101: data <= 18'h3fdc5; 
        10'b1011000110: data <= 18'h3ff2b; 
        10'b1011000111: data <= 18'h3fe6c; 
        10'b1011001000: data <= 18'h3ff11; 
        10'b1011001001: data <= 18'h3ff0d; 
        10'b1011001010: data <= 18'h3ffe8; 
        10'b1011001011: data <= 18'h0016a; 
        10'b1011001100: data <= 18'h00102; 
        10'b1011001101: data <= 18'h00148; 
        10'b1011001110: data <= 18'h00176; 
        10'b1011001111: data <= 18'h0003b; 
        10'b1011010000: data <= 18'h3ffb0; 
        10'b1011010001: data <= 18'h3fff6; 
        10'b1011010010: data <= 18'h3ff09; 
        10'b1011010011: data <= 18'h3ff12; 
        10'b1011010100: data <= 18'h3ffec; 
        10'b1011010101: data <= 18'h3ffbe; 
        10'b1011010110: data <= 18'h3ff67; 
        10'b1011010111: data <= 18'h3ffb9; 
        10'b1011011000: data <= 18'h3ffda; 
        10'b1011011001: data <= 18'h00005; 
        10'b1011011010: data <= 18'h3ff8e; 
        10'b1011011011: data <= 18'h3ff5a; 
        10'b1011011100: data <= 18'h3ff0e; 
        10'b1011011101: data <= 18'h3ff35; 
        10'b1011011110: data <= 18'h3fec9; 
        10'b1011011111: data <= 18'h3ffa8; 
        10'b1011100000: data <= 18'h3fee6; 
        10'b1011100001: data <= 18'h3ff10; 
        10'b1011100010: data <= 18'h3fede; 
        10'b1011100011: data <= 18'h3ff5a; 
        10'b1011100100: data <= 18'h3ff49; 
        10'b1011100101: data <= 18'h3ff65; 
        10'b1011100110: data <= 18'h3ff1a; 
        10'b1011100111: data <= 18'h3ff59; 
        10'b1011101000: data <= 18'h3ff37; 
        10'b1011101001: data <= 18'h3fef5; 
        10'b1011101010: data <= 18'h3fed6; 
        10'b1011101011: data <= 18'h3ff45; 
        10'b1011101100: data <= 18'h3ff7e; 
        10'b1011101101: data <= 18'h3ffd8; 
        10'b1011101110: data <= 18'h3ff8b; 
        10'b1011101111: data <= 18'h00035; 
        10'b1011110000: data <= 18'h00030; 
        10'b1011110001: data <= 18'h3ff20; 
        10'b1011110010: data <= 18'h3ffb9; 
        10'b1011110011: data <= 18'h3ffa2; 
        10'b1011110100: data <= 18'h3ffcd; 
        10'b1011110101: data <= 18'h3ff54; 
        10'b1011110110: data <= 18'h3ff94; 
        10'b1011110111: data <= 18'h3ffbc; 
        10'b1011111000: data <= 18'h3ffc5; 
        10'b1011111001: data <= 18'h3ff1a; 
        10'b1011111010: data <= 18'h3fff8; 
        10'b1011111011: data <= 18'h3ff65; 
        10'b1011111100: data <= 18'h00026; 
        10'b1011111101: data <= 18'h3ff8e; 
        10'b1011111110: data <= 18'h3ff3a; 
        10'b1011111111: data <= 18'h3ffeb; 
        10'b1100000000: data <= 18'h3ff5f; 
        10'b1100000001: data <= 18'h3ff3d; 
        10'b1100000010: data <= 18'h3ff87; 
        10'b1100000011: data <= 18'h3ffcc; 
        10'b1100000100: data <= 18'h3ffb8; 
        10'b1100000101: data <= 18'h00004; 
        10'b1100000110: data <= 18'h00020; 
        10'b1100000111: data <= 18'h0002d; 
        10'b1100001000: data <= 18'h3ffda; 
        10'b1100001001: data <= 18'h3ffbf; 
        10'b1100001010: data <= 18'h3ffd7; 
        10'b1100001011: data <= 18'h3ff4f; 
        10'b1100001100: data <= 18'h3ffae; 
        10'b1100001101: data <= 18'h00021; 
        10'b1100001110: data <= 18'h3ff2c; 
        10'b1100001111: data <= 18'h3ffb0; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 13) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 19'h7ff1a; 
        10'b0000000001: data <= 19'h7ff49; 
        10'b0000000010: data <= 19'h7ff21; 
        10'b0000000011: data <= 19'h7ff96; 
        10'b0000000100: data <= 19'h7ff7a; 
        10'b0000000101: data <= 19'h0002e; 
        10'b0000000110: data <= 19'h7fe2a; 
        10'b0000000111: data <= 19'h7ff9b; 
        10'b0000001000: data <= 19'h7fec4; 
        10'b0000001001: data <= 19'h7fef4; 
        10'b0000001010: data <= 19'h7fe87; 
        10'b0000001011: data <= 19'h00027; 
        10'b0000001100: data <= 19'h7ff6a; 
        10'b0000001101: data <= 19'h7ffe7; 
        10'b0000001110: data <= 19'h7fe79; 
        10'b0000001111: data <= 19'h7ffeb; 
        10'b0000010000: data <= 19'h7ff87; 
        10'b0000010001: data <= 19'h7fe5b; 
        10'b0000010010: data <= 19'h0002a; 
        10'b0000010011: data <= 19'h7ff47; 
        10'b0000010100: data <= 19'h7ff22; 
        10'b0000010101: data <= 19'h7ff15; 
        10'b0000010110: data <= 19'h7ff36; 
        10'b0000010111: data <= 19'h00057; 
        10'b0000011000: data <= 19'h00002; 
        10'b0000011001: data <= 19'h7fef2; 
        10'b0000011010: data <= 19'h7feb0; 
        10'b0000011011: data <= 19'h7ff2d; 
        10'b0000011100: data <= 19'h7ff22; 
        10'b0000011101: data <= 19'h7fe2c; 
        10'b0000011110: data <= 19'h0004f; 
        10'b0000011111: data <= 19'h00001; 
        10'b0000100000: data <= 19'h7fe55; 
        10'b0000100001: data <= 19'h7fe62; 
        10'b0000100010: data <= 19'h7fe3c; 
        10'b0000100011: data <= 19'h7fe63; 
        10'b0000100100: data <= 19'h0003a; 
        10'b0000100101: data <= 19'h7ff53; 
        10'b0000100110: data <= 19'h7ff41; 
        10'b0000100111: data <= 19'h7fe2f; 
        10'b0000101000: data <= 19'h00033; 
        10'b0000101001: data <= 19'h7ffb6; 
        10'b0000101010: data <= 19'h7fec3; 
        10'b0000101011: data <= 19'h7ff10; 
        10'b0000101100: data <= 19'h7ffb8; 
        10'b0000101101: data <= 19'h7ff69; 
        10'b0000101110: data <= 19'h7fe98; 
        10'b0000101111: data <= 19'h7ff77; 
        10'b0000110000: data <= 19'h0002d; 
        10'b0000110001: data <= 19'h7fe4b; 
        10'b0000110010: data <= 19'h7ffb2; 
        10'b0000110011: data <= 19'h7fe9c; 
        10'b0000110100: data <= 19'h7ffde; 
        10'b0000110101: data <= 19'h00061; 
        10'b0000110110: data <= 19'h7fec3; 
        10'b0000110111: data <= 19'h7fe99; 
        10'b0000111000: data <= 19'h7fe79; 
        10'b0000111001: data <= 19'h7fff9; 
        10'b0000111010: data <= 19'h7ff64; 
        10'b0000111011: data <= 19'h7ff3e; 
        10'b0000111100: data <= 19'h7fe8b; 
        10'b0000111101: data <= 19'h7fe35; 
        10'b0000111110: data <= 19'h7ff66; 
        10'b0000111111: data <= 19'h7fe28; 
        10'b0001000000: data <= 19'h00054; 
        10'b0001000001: data <= 19'h7fe26; 
        10'b0001000010: data <= 19'h7fe3d; 
        10'b0001000011: data <= 19'h7ffa3; 
        10'b0001000100: data <= 19'h7ff62; 
        10'b0001000101: data <= 19'h7fe1b; 
        10'b0001000110: data <= 19'h7ff9e; 
        10'b0001000111: data <= 19'h7ff7e; 
        10'b0001001000: data <= 19'h7fdfe; 
        10'b0001001001: data <= 19'h7fed2; 
        10'b0001001010: data <= 19'h7fed3; 
        10'b0001001011: data <= 19'h7ffc0; 
        10'b0001001100: data <= 19'h7fff1; 
        10'b0001001101: data <= 19'h7ffe8; 
        10'b0001001110: data <= 19'h7ff8f; 
        10'b0001001111: data <= 19'h7ff30; 
        10'b0001010000: data <= 19'h0002d; 
        10'b0001010001: data <= 19'h7fec2; 
        10'b0001010010: data <= 19'h7ffb8; 
        10'b0001010011: data <= 19'h0003c; 
        10'b0001010100: data <= 19'h7fea1; 
        10'b0001010101: data <= 19'h7ff35; 
        10'b0001010110: data <= 19'h7ff3a; 
        10'b0001010111: data <= 19'h7fe69; 
        10'b0001011000: data <= 19'h00052; 
        10'b0001011001: data <= 19'h7fe7f; 
        10'b0001011010: data <= 19'h7fe47; 
        10'b0001011011: data <= 19'h7fef7; 
        10'b0001011100: data <= 19'h7fe32; 
        10'b0001011101: data <= 19'h7ff5f; 
        10'b0001011110: data <= 19'h7fea5; 
        10'b0001011111: data <= 19'h7fd7c; 
        10'b0001100000: data <= 19'h7fd34; 
        10'b0001100001: data <= 19'h7fc9c; 
        10'b0001100010: data <= 19'h7fd30; 
        10'b0001100011: data <= 19'h7fe55; 
        10'b0001100100: data <= 19'h7fd2d; 
        10'b0001100101: data <= 19'h7fdcf; 
        10'b0001100110: data <= 19'h7fe79; 
        10'b0001100111: data <= 19'h7ff10; 
        10'b0001101000: data <= 19'h7fddd; 
        10'b0001101001: data <= 19'h00022; 
        10'b0001101010: data <= 19'h7fee2; 
        10'b0001101011: data <= 19'h7ffe3; 
        10'b0001101100: data <= 19'h7fec8; 
        10'b0001101101: data <= 19'h7ff9c; 
        10'b0001101110: data <= 19'h7ff6e; 
        10'b0001101111: data <= 19'h7fe53; 
        10'b0001110000: data <= 19'h7ff45; 
        10'b0001110001: data <= 19'h7ffca; 
        10'b0001110010: data <= 19'h7fef3; 
        10'b0001110011: data <= 19'h7fe54; 
        10'b0001110100: data <= 19'h7ffe9; 
        10'b0001110101: data <= 19'h7ffdf; 
        10'b0001110110: data <= 19'h7ff46; 
        10'b0001110111: data <= 19'h7fe7c; 
        10'b0001111000: data <= 19'h7fe7a; 
        10'b0001111001: data <= 19'h7ff1b; 
        10'b0001111010: data <= 19'h7ff35; 
        10'b0001111011: data <= 19'h7ff90; 
        10'b0001111100: data <= 19'h0026f; 
        10'b0001111101: data <= 19'h00192; 
        10'b0001111110: data <= 19'h0054c; 
        10'b0001111111: data <= 19'h00405; 
        10'b0010000000: data <= 19'h001d4; 
        10'b0010000001: data <= 19'h00100; 
        10'b0010000010: data <= 19'h00180; 
        10'b0010000011: data <= 19'h7feaa; 
        10'b0010000100: data <= 19'h7fe60; 
        10'b0010000101: data <= 19'h7ff28; 
        10'b0010000110: data <= 19'h7fd8c; 
        10'b0010000111: data <= 19'h7fe3e; 
        10'b0010001000: data <= 19'h7fff2; 
        10'b0010001001: data <= 19'h0001e; 
        10'b0010001010: data <= 19'h7ff0d; 
        10'b0010001011: data <= 19'h7ff45; 
        10'b0010001100: data <= 19'h7ff4e; 
        10'b0010001101: data <= 19'h7ffac; 
        10'b0010001110: data <= 19'h7ffcb; 
        10'b0010001111: data <= 19'h7fff0; 
        10'b0010010000: data <= 19'h7fe8e; 
        10'b0010010001: data <= 19'h7ff26; 
        10'b0010010010: data <= 19'h7fec1; 
        10'b0010010011: data <= 19'h7fca3; 
        10'b0010010100: data <= 19'h7fea6; 
        10'b0010010101: data <= 19'h00133; 
        10'b0010010110: data <= 19'h7fd38; 
        10'b0010010111: data <= 19'h003b4; 
        10'b0010011000: data <= 19'h006f6; 
        10'b0010011001: data <= 19'h005ca; 
        10'b0010011010: data <= 19'h00606; 
        10'b0010011011: data <= 19'h002e0; 
        10'b0010011100: data <= 19'h0025f; 
        10'b0010011101: data <= 19'h00593; 
        10'b0010011110: data <= 19'h00047; 
        10'b0010011111: data <= 19'h7ffbf; 
        10'b0010100000: data <= 19'h001fd; 
        10'b0010100001: data <= 19'h00108; 
        10'b0010100010: data <= 19'h7fc9f; 
        10'b0010100011: data <= 19'h7fd2a; 
        10'b0010100100: data <= 19'h7fe0a; 
        10'b0010100101: data <= 19'h0017f; 
        10'b0010100110: data <= 19'h7ff64; 
        10'b0010100111: data <= 19'h00042; 
        10'b0010101000: data <= 19'h7fea1; 
        10'b0010101001: data <= 19'h7fe84; 
        10'b0010101010: data <= 19'h7fe32; 
        10'b0010101011: data <= 19'h7fe3c; 
        10'b0010101100: data <= 19'h7fdfa; 
        10'b0010101101: data <= 19'h7fe05; 
        10'b0010101110: data <= 19'h7fcd2; 
        10'b0010101111: data <= 19'h7fccf; 
        10'b0010110000: data <= 19'h00039; 
        10'b0010110001: data <= 19'h000f0; 
        10'b0010110010: data <= 19'h7ffc1; 
        10'b0010110011: data <= 19'h001cb; 
        10'b0010110100: data <= 19'h002d6; 
        10'b0010110101: data <= 19'h00246; 
        10'b0010110110: data <= 19'h00334; 
        10'b0010110111: data <= 19'h005ff; 
        10'b0010111000: data <= 19'h002e7; 
        10'b0010111001: data <= 19'h00369; 
        10'b0010111010: data <= 19'h000b8; 
        10'b0010111011: data <= 19'h003e5; 
        10'b0010111100: data <= 19'h0017c; 
        10'b0010111101: data <= 19'h001d4; 
        10'b0010111110: data <= 19'h00246; 
        10'b0010111111: data <= 19'h0021f; 
        10'b0011000000: data <= 19'h001ca; 
        10'b0011000001: data <= 19'h000c1; 
        10'b0011000010: data <= 19'h7ff45; 
        10'b0011000011: data <= 19'h7ffd1; 
        10'b0011000100: data <= 19'h00044; 
        10'b0011000101: data <= 19'h7fea4; 
        10'b0011000110: data <= 19'h7fe68; 
        10'b0011000111: data <= 19'h7fec2; 
        10'b0011001000: data <= 19'h7fde4; 
        10'b0011001001: data <= 19'h7ff3b; 
        10'b0011001010: data <= 19'h7fdd5; 
        10'b0011001011: data <= 19'h7ffdf; 
        10'b0011001100: data <= 19'h00225; 
        10'b0011001101: data <= 19'h000e0; 
        10'b0011001110: data <= 19'h00114; 
        10'b0011001111: data <= 19'h7ff53; 
        10'b0011010000: data <= 19'h7fd42; 
        10'b0011010001: data <= 19'h7fdf2; 
        10'b0011010010: data <= 19'h7fcfa; 
        10'b0011010011: data <= 19'h001d1; 
        10'b0011010100: data <= 19'h00247; 
        10'b0011010101: data <= 19'h7ffdc; 
        10'b0011010110: data <= 19'h0018d; 
        10'b0011010111: data <= 19'h7fe4e; 
        10'b0011011000: data <= 19'h00253; 
        10'b0011011001: data <= 19'h0039f; 
        10'b0011011010: data <= 19'h000a7; 
        10'b0011011011: data <= 19'h00781; 
        10'b0011011100: data <= 19'h00499; 
        10'b0011011101: data <= 19'h7ffd3; 
        10'b0011011110: data <= 19'h0001c; 
        10'b0011011111: data <= 19'h7ffaf; 
        10'b0011100000: data <= 19'h7ffae; 
        10'b0011100001: data <= 19'h0001a; 
        10'b0011100010: data <= 19'h7ffa1; 
        10'b0011100011: data <= 19'h7fe85; 
        10'b0011100100: data <= 19'h7ff9b; 
        10'b0011100101: data <= 19'h7ff4e; 
        10'b0011100110: data <= 19'h0031c; 
        10'b0011100111: data <= 19'h001ec; 
        10'b0011101000: data <= 19'h000b1; 
        10'b0011101001: data <= 19'h00565; 
        10'b0011101010: data <= 19'h0004f; 
        10'b0011101011: data <= 19'h0002e; 
        10'b0011101100: data <= 19'h0039a; 
        10'b0011101101: data <= 19'h004ab; 
        10'b0011101110: data <= 19'h7fc51; 
        10'b0011101111: data <= 19'h7fcdf; 
        10'b0011110000: data <= 19'h0028d; 
        10'b0011110001: data <= 19'h7fe31; 
        10'b0011110010: data <= 19'h000d9; 
        10'b0011110011: data <= 19'h00271; 
        10'b0011110100: data <= 19'h0019d; 
        10'b0011110101: data <= 19'h004f9; 
        10'b0011110110: data <= 19'h00356; 
        10'b0011110111: data <= 19'h005ab; 
        10'b0011111000: data <= 19'h00528; 
        10'b0011111001: data <= 19'h7ff63; 
        10'b0011111010: data <= 19'h7ff90; 
        10'b0011111011: data <= 19'h00082; 
        10'b0011111100: data <= 19'h00008; 
        10'b0011111101: data <= 19'h0001a; 
        10'b0011111110: data <= 19'h7ff31; 
        10'b0011111111: data <= 19'h7ff01; 
        10'b0100000000: data <= 19'h7ff75; 
        10'b0100000001: data <= 19'h00326; 
        10'b0100000010: data <= 19'h00256; 
        10'b0100000011: data <= 19'h004d0; 
        10'b0100000100: data <= 19'h00675; 
        10'b0100000101: data <= 19'h00572; 
        10'b0100000110: data <= 19'h00373; 
        10'b0100000111: data <= 19'h00610; 
        10'b0100001000: data <= 19'h001a5; 
        10'b0100001001: data <= 19'h001c1; 
        10'b0100001010: data <= 19'h7f8e8; 
        10'b0100001011: data <= 19'h7f623; 
        10'b0100001100: data <= 19'h7fc90; 
        10'b0100001101: data <= 19'h00087; 
        10'b0100001110: data <= 19'h00112; 
        10'b0100001111: data <= 19'h001ea; 
        10'b0100010000: data <= 19'h00287; 
        10'b0100010001: data <= 19'h0022e; 
        10'b0100010010: data <= 19'h00536; 
        10'b0100010011: data <= 19'h0055a; 
        10'b0100010100: data <= 19'h7ff21; 
        10'b0100010101: data <= 19'h7ff44; 
        10'b0100010110: data <= 19'h00131; 
        10'b0100010111: data <= 19'h7fe5e; 
        10'b0100011000: data <= 19'h7feb4; 
        10'b0100011001: data <= 19'h0000d; 
        10'b0100011010: data <= 19'h7fe9f; 
        10'b0100011011: data <= 19'h00023; 
        10'b0100011100: data <= 19'h00137; 
        10'b0100011101: data <= 19'h003df; 
        10'b0100011110: data <= 19'h003d8; 
        10'b0100011111: data <= 19'h0070c; 
        10'b0100100000: data <= 19'h0053b; 
        10'b0100100001: data <= 19'h0061d; 
        10'b0100100010: data <= 19'h008ef; 
        10'b0100100011: data <= 19'h00448; 
        10'b0100100100: data <= 19'h0047a; 
        10'b0100100101: data <= 19'h003a6; 
        10'b0100100110: data <= 19'h7fed1; 
        10'b0100100111: data <= 19'h7f69c; 
        10'b0100101000: data <= 19'h7f84e; 
        10'b0100101001: data <= 19'h7fda8; 
        10'b0100101010: data <= 19'h002ad; 
        10'b0100101011: data <= 19'h002aa; 
        10'b0100101100: data <= 19'h002bb; 
        10'b0100101101: data <= 19'h0065b; 
        10'b0100101110: data <= 19'h00708; 
        10'b0100101111: data <= 19'h005bc; 
        10'b0100110000: data <= 19'h00013; 
        10'b0100110001: data <= 19'h7ff95; 
        10'b0100110010: data <= 19'h7ff41; 
        10'b0100110011: data <= 19'h7fec3; 
        10'b0100110100: data <= 19'h7fe9f; 
        10'b0100110101: data <= 19'h00050; 
        10'b0100110110: data <= 19'h7ffe0; 
        10'b0100110111: data <= 19'h7fdd3; 
        10'b0100111000: data <= 19'h001d8; 
        10'b0100111001: data <= 19'h00445; 
        10'b0100111010: data <= 19'h00822; 
        10'b0100111011: data <= 19'h00a8e; 
        10'b0100111100: data <= 19'h0084c; 
        10'b0100111101: data <= 19'h00a7c; 
        10'b0100111110: data <= 19'h0072e; 
        10'b0100111111: data <= 19'h00365; 
        10'b0101000000: data <= 19'h0045f; 
        10'b0101000001: data <= 19'h00a70; 
        10'b0101000010: data <= 19'h00cb6; 
        10'b0101000011: data <= 19'h7fe70; 
        10'b0101000100: data <= 19'h7f86f; 
        10'b0101000101: data <= 19'h7fd66; 
        10'b0101000110: data <= 19'h7fd86; 
        10'b0101000111: data <= 19'h0010b; 
        10'b0101001000: data <= 19'h005c0; 
        10'b0101001001: data <= 19'h006e3; 
        10'b0101001010: data <= 19'h00926; 
        10'b0101001011: data <= 19'h008a3; 
        10'b0101001100: data <= 19'h00602; 
        10'b0101001101: data <= 19'h000fa; 
        10'b0101001110: data <= 19'h00087; 
        10'b0101001111: data <= 19'h7ff82; 
        10'b0101010000: data <= 19'h7fecd; 
        10'b0101010001: data <= 19'h7ff98; 
        10'b0101010010: data <= 19'h7fefc; 
        10'b0101010011: data <= 19'h7ff87; 
        10'b0101010100: data <= 19'h7ff9d; 
        10'b0101010101: data <= 19'h0051b; 
        10'b0101010110: data <= 19'h0043c; 
        10'b0101010111: data <= 19'h00677; 
        10'b0101011000: data <= 19'h0061a; 
        10'b0101011001: data <= 19'h007ab; 
        10'b0101011010: data <= 19'h0014e; 
        10'b0101011011: data <= 19'h001d4; 
        10'b0101011100: data <= 19'h00104; 
        10'b0101011101: data <= 19'h00c9b; 
        10'b0101011110: data <= 19'h00cab; 
        10'b0101011111: data <= 19'h002d7; 
        10'b0101100000: data <= 19'h0007b; 
        10'b0101100001: data <= 19'h7fee4; 
        10'b0101100010: data <= 19'h7ff17; 
        10'b0101100011: data <= 19'h0032c; 
        10'b0101100100: data <= 19'h00564; 
        10'b0101100101: data <= 19'h00943; 
        10'b0101100110: data <= 19'h00ac9; 
        10'b0101100111: data <= 19'h00900; 
        10'b0101101000: data <= 19'h005a6; 
        10'b0101101001: data <= 19'h00243; 
        10'b0101101010: data <= 19'h0011f; 
        10'b0101101011: data <= 19'h7fe69; 
        10'b0101101100: data <= 19'h7fe3f; 
        10'b0101101101: data <= 19'h7ff5e; 
        10'b0101101110: data <= 19'h0005b; 
        10'b0101101111: data <= 19'h7fe7f; 
        10'b0101110000: data <= 19'h7fedc; 
        10'b0101110001: data <= 19'h7fff9; 
        10'b0101110010: data <= 19'h7ff2e; 
        10'b0101110011: data <= 19'h7ff3b; 
        10'b0101110100: data <= 19'h000b2; 
        10'b0101110101: data <= 19'h7ff12; 
        10'b0101110110: data <= 19'h7fd3d; 
        10'b0101110111: data <= 19'h0010d; 
        10'b0101111000: data <= 19'h004a1; 
        10'b0101111001: data <= 19'h00bcf; 
        10'b0101111010: data <= 19'h00388; 
        10'b0101111011: data <= 19'h008af; 
        10'b0101111100: data <= 19'h00375; 
        10'b0101111101: data <= 19'h7fdce; 
        10'b0101111110: data <= 19'h00035; 
        10'b0101111111: data <= 19'h0004a; 
        10'b0110000000: data <= 19'h003d8; 
        10'b0110000001: data <= 19'h0037d; 
        10'b0110000010: data <= 19'h001fb; 
        10'b0110000011: data <= 19'h002d0; 
        10'b0110000100: data <= 19'h0017f; 
        10'b0110000101: data <= 19'h00055; 
        10'b0110000110: data <= 19'h00057; 
        10'b0110000111: data <= 19'h7ffb6; 
        10'b0110001000: data <= 19'h7feee; 
        10'b0110001001: data <= 19'h7fe37; 
        10'b0110001010: data <= 19'h7ffc2; 
        10'b0110001011: data <= 19'h7ff42; 
        10'b0110001100: data <= 19'h7fe6d; 
        10'b0110001101: data <= 19'h7fc92; 
        10'b0110001110: data <= 19'h7f9e0; 
        10'b0110001111: data <= 19'h7f826; 
        10'b0110010000: data <= 19'h7f6bb; 
        10'b0110010001: data <= 19'h7f893; 
        10'b0110010010: data <= 19'h7fef6; 
        10'b0110010011: data <= 19'h004bf; 
        10'b0110010100: data <= 19'h00491; 
        10'b0110010101: data <= 19'h009a7; 
        10'b0110010110: data <= 19'h007b8; 
        10'b0110010111: data <= 19'h00538; 
        10'b0110011000: data <= 19'h7ff5d; 
        10'b0110011001: data <= 19'h000a6; 
        10'b0110011010: data <= 19'h7fea5; 
        10'b0110011011: data <= 19'h7fcda; 
        10'b0110011100: data <= 19'h7fae0; 
        10'b0110011101: data <= 19'h7fb6a; 
        10'b0110011110: data <= 19'h7fc0f; 
        10'b0110011111: data <= 19'h7fb57; 
        10'b0110100000: data <= 19'h7fde3; 
        10'b0110100001: data <= 19'h7ffb1; 
        10'b0110100010: data <= 19'h7fe1d; 
        10'b0110100011: data <= 19'h0000e; 
        10'b0110100100: data <= 19'h00026; 
        10'b0110100101: data <= 19'h7fedb; 
        10'b0110100110: data <= 19'h7feaf; 
        10'b0110100111: data <= 19'h7ff73; 
        10'b0110101000: data <= 19'h7fe47; 
        10'b0110101001: data <= 19'h7fc98; 
        10'b0110101010: data <= 19'h7f85f; 
        10'b0110101011: data <= 19'h7f6a6; 
        10'b0110101100: data <= 19'h7f77a; 
        10'b0110101101: data <= 19'h7fdec; 
        10'b0110101110: data <= 19'h00052; 
        10'b0110101111: data <= 19'h00035; 
        10'b0110110000: data <= 19'h00698; 
        10'b0110110001: data <= 19'h007cb; 
        10'b0110110010: data <= 19'h006d2; 
        10'b0110110011: data <= 19'h003ef; 
        10'b0110110100: data <= 19'h7fe07; 
        10'b0110110101: data <= 19'h7fe48; 
        10'b0110110110: data <= 19'h7fecc; 
        10'b0110110111: data <= 19'h7f918; 
        10'b0110111000: data <= 19'h7f767; 
        10'b0110111001: data <= 19'h7f968; 
        10'b0110111010: data <= 19'h7fbd1; 
        10'b0110111011: data <= 19'h7fc05; 
        10'b0110111100: data <= 19'h7fcff; 
        10'b0110111101: data <= 19'h7ff7b; 
        10'b0110111110: data <= 19'h7fdec; 
        10'b0110111111: data <= 19'h0002b; 
        10'b0111000000: data <= 19'h7ff14; 
        10'b0111000001: data <= 19'h7fe4c; 
        10'b0111000010: data <= 19'h7fed3; 
        10'b0111000011: data <= 19'h7ff61; 
        10'b0111000100: data <= 19'h7fd3e; 
        10'b0111000101: data <= 19'h7fb12; 
        10'b0111000110: data <= 19'h7f813; 
        10'b0111000111: data <= 19'h7fb52; 
        10'b0111001000: data <= 19'h00324; 
        10'b0111001001: data <= 19'h0037e; 
        10'b0111001010: data <= 19'h0016e; 
        10'b0111001011: data <= 19'h00333; 
        10'b0111001100: data <= 19'h00660; 
        10'b0111001101: data <= 19'h00596; 
        10'b0111001110: data <= 19'h00201; 
        10'b0111001111: data <= 19'h00355; 
        10'b0111010000: data <= 19'h00121; 
        10'b0111010001: data <= 19'h7fd64; 
        10'b0111010010: data <= 19'h7fa6e; 
        10'b0111010011: data <= 19'h7f80a; 
        10'b0111010100: data <= 19'h7f80a; 
        10'b0111010101: data <= 19'h7f7e9; 
        10'b0111010110: data <= 19'h7f983; 
        10'b0111010111: data <= 19'h7fdd9; 
        10'b0111011000: data <= 19'h7fd2a; 
        10'b0111011001: data <= 19'h7ff08; 
        10'b0111011010: data <= 19'h7fefe; 
        10'b0111011011: data <= 19'h7fe40; 
        10'b0111011100: data <= 19'h00064; 
        10'b0111011101: data <= 19'h00045; 
        10'b0111011110: data <= 19'h7fea2; 
        10'b0111011111: data <= 19'h7fe54; 
        10'b0111100000: data <= 19'h7fe2d; 
        10'b0111100001: data <= 19'h7fae5; 
        10'b0111100010: data <= 19'h7f901; 
        10'b0111100011: data <= 19'h0013d; 
        10'b0111100100: data <= 19'h00681; 
        10'b0111100101: data <= 19'h0080f; 
        10'b0111100110: data <= 19'h00294; 
        10'b0111100111: data <= 19'h00619; 
        10'b0111101000: data <= 19'h009ed; 
        10'b0111101001: data <= 19'h00605; 
        10'b0111101010: data <= 19'h00082; 
        10'b0111101011: data <= 19'h7fe63; 
        10'b0111101100: data <= 19'h000b9; 
        10'b0111101101: data <= 19'h7fce9; 
        10'b0111101110: data <= 19'h7f7d1; 
        10'b0111101111: data <= 19'h7fc20; 
        10'b0111110000: data <= 19'h7fc27; 
        10'b0111110001: data <= 19'h7fa90; 
        10'b0111110010: data <= 19'h7fbf9; 
        10'b0111110011: data <= 19'h7fd77; 
        10'b0111110100: data <= 19'h7fe8e; 
        10'b0111110101: data <= 19'h7fdf0; 
        10'b0111110110: data <= 19'h7ffa9; 
        10'b0111110111: data <= 19'h7feee; 
        10'b0111111000: data <= 19'h7fec3; 
        10'b0111111001: data <= 19'h00014; 
        10'b0111111010: data <= 19'h7fe3b; 
        10'b0111111011: data <= 19'h7fdbb; 
        10'b0111111100: data <= 19'h7fce3; 
        10'b0111111101: data <= 19'h7fcd0; 
        10'b0111111110: data <= 19'h7fe07; 
        10'b0111111111: data <= 19'h001ec; 
        10'b1000000000: data <= 19'h00559; 
        10'b1000000001: data <= 19'h009a7; 
        10'b1000000010: data <= 19'h006bf; 
        10'b1000000011: data <= 19'h00934; 
        10'b1000000100: data <= 19'h005fe; 
        10'b1000000101: data <= 19'h00374; 
        10'b1000000110: data <= 19'h7fbd1; 
        10'b1000000111: data <= 19'h7feeb; 
        10'b1000001000: data <= 19'h7fda5; 
        10'b1000001001: data <= 19'h7f9b8; 
        10'b1000001010: data <= 19'h7fe7d; 
        10'b1000001011: data <= 19'h7fed1; 
        10'b1000001100: data <= 19'h00077; 
        10'b1000001101: data <= 19'h7fc8b; 
        10'b1000001110: data <= 19'h7ff7a; 
        10'b1000001111: data <= 19'h7fd10; 
        10'b1000010000: data <= 19'h7fc02; 
        10'b1000010001: data <= 19'h7fdf3; 
        10'b1000010010: data <= 19'h7ffac; 
        10'b1000010011: data <= 19'h00041; 
        10'b1000010100: data <= 19'h7feca; 
        10'b1000010101: data <= 19'h7ff66; 
        10'b1000010110: data <= 19'h7ff8d; 
        10'b1000010111: data <= 19'h7fd4c; 
        10'b1000011000: data <= 19'h7fc8d; 
        10'b1000011001: data <= 19'h7fe9c; 
        10'b1000011010: data <= 19'h000ec; 
        10'b1000011011: data <= 19'h0028d; 
        10'b1000011100: data <= 19'h002a8; 
        10'b1000011101: data <= 19'h00689; 
        10'b1000011110: data <= 19'h0035b; 
        10'b1000011111: data <= 19'h7ff89; 
        10'b1000100000: data <= 19'h00199; 
        10'b1000100001: data <= 19'h7fba0; 
        10'b1000100010: data <= 19'h7fae0; 
        10'b1000100011: data <= 19'h7fe0a; 
        10'b1000100100: data <= 19'h7fe64; 
        10'b1000100101: data <= 19'h7fde6; 
        10'b1000100110: data <= 19'h0019d; 
        10'b1000100111: data <= 19'h00077; 
        10'b1000101000: data <= 19'h00213; 
        10'b1000101001: data <= 19'h0002d; 
        10'b1000101010: data <= 19'h00158; 
        10'b1000101011: data <= 19'h7feda; 
        10'b1000101100: data <= 19'h7fcf4; 
        10'b1000101101: data <= 19'h7fe2e; 
        10'b1000101110: data <= 19'h7fe73; 
        10'b1000101111: data <= 19'h0002f; 
        10'b1000110000: data <= 19'h7fe83; 
        10'b1000110001: data <= 19'h7ffad; 
        10'b1000110010: data <= 19'h7fea3; 
        10'b1000110011: data <= 19'h7fe04; 
        10'b1000110100: data <= 19'h7fc04; 
        10'b1000110101: data <= 19'h7ff54; 
        10'b1000110110: data <= 19'h000a3; 
        10'b1000110111: data <= 19'h005a8; 
        10'b1000111000: data <= 19'h001b0; 
        10'b1000111001: data <= 19'h7ff45; 
        10'b1000111010: data <= 19'h7fff8; 
        10'b1000111011: data <= 19'h7fb38; 
        10'b1000111100: data <= 19'h0004d; 
        10'b1000111101: data <= 19'h7ffe0; 
        10'b1000111110: data <= 19'h7fb76; 
        10'b1000111111: data <= 19'h7ff2d; 
        10'b1001000000: data <= 19'h7fab3; 
        10'b1001000001: data <= 19'h7fe52; 
        10'b1001000010: data <= 19'h000f0; 
        10'b1001000011: data <= 19'h00095; 
        10'b1001000100: data <= 19'h001ae; 
        10'b1001000101: data <= 19'h002d9; 
        10'b1001000110: data <= 19'h002d7; 
        10'b1001000111: data <= 19'h7ff4c; 
        10'b1001001000: data <= 19'h7fe21; 
        10'b1001001001: data <= 19'h7fd8b; 
        10'b1001001010: data <= 19'h7ff46; 
        10'b1001001011: data <= 19'h7fe91; 
        10'b1001001100: data <= 19'h00021; 
        10'b1001001101: data <= 19'h7ff35; 
        10'b1001001110: data <= 19'h00048; 
        10'b1001001111: data <= 19'h7fcdf; 
        10'b1001010000: data <= 19'h7fb5a; 
        10'b1001010001: data <= 19'h7ff89; 
        10'b1001010010: data <= 19'h00273; 
        10'b1001010011: data <= 19'h0053c; 
        10'b1001010100: data <= 19'h00118; 
        10'b1001010101: data <= 19'h0023e; 
        10'b1001010110: data <= 19'h7ff96; 
        10'b1001010111: data <= 19'h7fc8c; 
        10'b1001011000: data <= 19'h7fe11; 
        10'b1001011001: data <= 19'h00131; 
        10'b1001011010: data <= 19'h7ffe5; 
        10'b1001011011: data <= 19'h7ff74; 
        10'b1001011100: data <= 19'h7fbf1; 
        10'b1001011101: data <= 19'h7fe4c; 
        10'b1001011110: data <= 19'h7fede; 
        10'b1001011111: data <= 19'h7ffd6; 
        10'b1001100000: data <= 19'h7ffe8; 
        10'b1001100001: data <= 19'h000f9; 
        10'b1001100010: data <= 19'h000d7; 
        10'b1001100011: data <= 19'h7fec8; 
        10'b1001100100: data <= 19'h7fe87; 
        10'b1001100101: data <= 19'h7ffe9; 
        10'b1001100110: data <= 19'h7ffb2; 
        10'b1001100111: data <= 19'h7ff0f; 
        10'b1001101000: data <= 19'h7ff87; 
        10'b1001101001: data <= 19'h7fe39; 
        10'b1001101010: data <= 19'h7fedd; 
        10'b1001101011: data <= 19'h7fe02; 
        10'b1001101100: data <= 19'h7fc4a; 
        10'b1001101101: data <= 19'h7fa77; 
        10'b1001101110: data <= 19'h000a8; 
        10'b1001101111: data <= 19'h0017d; 
        10'b1001110000: data <= 19'h7ffa9; 
        10'b1001110001: data <= 19'h7fe3b; 
        10'b1001110010: data <= 19'h0011f; 
        10'b1001110011: data <= 19'h00066; 
        10'b1001110100: data <= 19'h0069c; 
        10'b1001110101: data <= 19'h006ee; 
        10'b1001110110: data <= 19'h004e6; 
        10'b1001110111: data <= 19'h003d4; 
        10'b1001111000: data <= 19'h7ffac; 
        10'b1001111001: data <= 19'h7ffa3; 
        10'b1001111010: data <= 19'h001a8; 
        10'b1001111011: data <= 19'h7fdf1; 
        10'b1001111100: data <= 19'h7fdc6; 
        10'b1001111101: data <= 19'h000f3; 
        10'b1001111110: data <= 19'h7ff9a; 
        10'b1001111111: data <= 19'h7fe95; 
        10'b1010000000: data <= 19'h7ffa5; 
        10'b1010000001: data <= 19'h7ffa3; 
        10'b1010000010: data <= 19'h7ff97; 
        10'b1010000011: data <= 19'h7fea1; 
        10'b1010000100: data <= 19'h7fe9c; 
        10'b1010000101: data <= 19'h7ffd3; 
        10'b1010000110: data <= 19'h7ff5f; 
        10'b1010000111: data <= 19'h7fe3b; 
        10'b1010001000: data <= 19'h7fc1e; 
        10'b1010001001: data <= 19'h7f6bf; 
        10'b1010001010: data <= 19'h7f8be; 
        10'b1010001011: data <= 19'h7fc58; 
        10'b1010001100: data <= 19'h00143; 
        10'b1010001101: data <= 19'h0013f; 
        10'b1010001110: data <= 19'h002af; 
        10'b1010001111: data <= 19'h00381; 
        10'b1010010000: data <= 19'h007d3; 
        10'b1010010001: data <= 19'h00b40; 
        10'b1010010010: data <= 19'h00993; 
        10'b1010010011: data <= 19'h007a2; 
        10'b1010010100: data <= 19'h0062e; 
        10'b1010010101: data <= 19'h0046e; 
        10'b1010010110: data <= 19'h00384; 
        10'b1010010111: data <= 19'h0047f; 
        10'b1010011000: data <= 19'h00351; 
        10'b1010011001: data <= 19'h000cc; 
        10'b1010011010: data <= 19'h7ff95; 
        10'b1010011011: data <= 19'h7fef4; 
        10'b1010011100: data <= 19'h7fdf4; 
        10'b1010011101: data <= 19'h7ffcf; 
        10'b1010011110: data <= 19'h7fe30; 
        10'b1010011111: data <= 19'h7ffa4; 
        10'b1010100000: data <= 19'h7ffc7; 
        10'b1010100001: data <= 19'h7ffa4; 
        10'b1010100010: data <= 19'h00058; 
        10'b1010100011: data <= 19'h7fe69; 
        10'b1010100100: data <= 19'h7fe64; 
        10'b1010100101: data <= 19'h7f9e0; 
        10'b1010100110: data <= 19'h7f781; 
        10'b1010100111: data <= 19'h7f8dd; 
        10'b1010101000: data <= 19'h7ff90; 
        10'b1010101001: data <= 19'h001ab; 
        10'b1010101010: data <= 19'h7ff5e; 
        10'b1010101011: data <= 19'h00308; 
        10'b1010101100: data <= 19'h0023c; 
        10'b1010101101: data <= 19'h00179; 
        10'b1010101110: data <= 19'h003b6; 
        10'b1010101111: data <= 19'h00810; 
        10'b1010110000: data <= 19'h0088f; 
        10'b1010110001: data <= 19'h005bf; 
        10'b1010110010: data <= 19'h0080d; 
        10'b1010110011: data <= 19'h0078e; 
        10'b1010110100: data <= 19'h0027d; 
        10'b1010110101: data <= 19'h00025; 
        10'b1010110110: data <= 19'h7fe4a; 
        10'b1010110111: data <= 19'h0002c; 
        10'b1010111000: data <= 19'h7ff4c; 
        10'b1010111001: data <= 19'h7fed3; 
        10'b1010111010: data <= 19'h00047; 
        10'b1010111011: data <= 19'h7ff88; 
        10'b1010111100: data <= 19'h0005f; 
        10'b1010111101: data <= 19'h7ffbb; 
        10'b1010111110: data <= 19'h0002e; 
        10'b1010111111: data <= 19'h7fe65; 
        10'b1011000000: data <= 19'h7fec9; 
        10'b1011000001: data <= 19'h7fdba; 
        10'b1011000010: data <= 19'h7fccb; 
        10'b1011000011: data <= 19'h7fc03; 
        10'b1011000100: data <= 19'h7fb8e; 
        10'b1011000101: data <= 19'h7fb8a; 
        10'b1011000110: data <= 19'h7fe55; 
        10'b1011000111: data <= 19'h7fcd9; 
        10'b1011001000: data <= 19'h7fe22; 
        10'b1011001001: data <= 19'h7fe1b; 
        10'b1011001010: data <= 19'h7ffd0; 
        10'b1011001011: data <= 19'h002d5; 
        10'b1011001100: data <= 19'h00204; 
        10'b1011001101: data <= 19'h00290; 
        10'b1011001110: data <= 19'h002eb; 
        10'b1011001111: data <= 19'h00076; 
        10'b1011010000: data <= 19'h7ff61; 
        10'b1011010001: data <= 19'h7ffec; 
        10'b1011010010: data <= 19'h7fe11; 
        10'b1011010011: data <= 19'h7fe24; 
        10'b1011010100: data <= 19'h7ffd7; 
        10'b1011010101: data <= 19'h7ff7c; 
        10'b1011010110: data <= 19'h7fece; 
        10'b1011010111: data <= 19'h7ff72; 
        10'b1011011000: data <= 19'h7ffb4; 
        10'b1011011001: data <= 19'h0000b; 
        10'b1011011010: data <= 19'h7ff1c; 
        10'b1011011011: data <= 19'h7feb4; 
        10'b1011011100: data <= 19'h7fe1c; 
        10'b1011011101: data <= 19'h7fe6a; 
        10'b1011011110: data <= 19'h7fd92; 
        10'b1011011111: data <= 19'h7ff51; 
        10'b1011100000: data <= 19'h7fdcd; 
        10'b1011100001: data <= 19'h7fe20; 
        10'b1011100010: data <= 19'h7fdbc; 
        10'b1011100011: data <= 19'h7feb5; 
        10'b1011100100: data <= 19'h7fe93; 
        10'b1011100101: data <= 19'h7fec9; 
        10'b1011100110: data <= 19'h7fe34; 
        10'b1011100111: data <= 19'h7feb3; 
        10'b1011101000: data <= 19'h7fe6e; 
        10'b1011101001: data <= 19'h7fdea; 
        10'b1011101010: data <= 19'h7fdac; 
        10'b1011101011: data <= 19'h7fe8a; 
        10'b1011101100: data <= 19'h7fefd; 
        10'b1011101101: data <= 19'h7ffaf; 
        10'b1011101110: data <= 19'h7ff16; 
        10'b1011101111: data <= 19'h0006a; 
        10'b1011110000: data <= 19'h00060; 
        10'b1011110001: data <= 19'h7fe41; 
        10'b1011110010: data <= 19'h7ff72; 
        10'b1011110011: data <= 19'h7ff43; 
        10'b1011110100: data <= 19'h7ff9b; 
        10'b1011110101: data <= 19'h7fea8; 
        10'b1011110110: data <= 19'h7ff29; 
        10'b1011110111: data <= 19'h7ff78; 
        10'b1011111000: data <= 19'h7ff8a; 
        10'b1011111001: data <= 19'h7fe34; 
        10'b1011111010: data <= 19'h7ffef; 
        10'b1011111011: data <= 19'h7fecb; 
        10'b1011111100: data <= 19'h0004c; 
        10'b1011111101: data <= 19'h7ff1d; 
        10'b1011111110: data <= 19'h7fe73; 
        10'b1011111111: data <= 19'h7ffd6; 
        10'b1100000000: data <= 19'h7febd; 
        10'b1100000001: data <= 19'h7fe7a; 
        10'b1100000010: data <= 19'h7ff0e; 
        10'b1100000011: data <= 19'h7ff98; 
        10'b1100000100: data <= 19'h7ff6f; 
        10'b1100000101: data <= 19'h00008; 
        10'b1100000110: data <= 19'h0003f; 
        10'b1100000111: data <= 19'h0005a; 
        10'b1100001000: data <= 19'h7ffb3; 
        10'b1100001001: data <= 19'h7ff7e; 
        10'b1100001010: data <= 19'h7ffae; 
        10'b1100001011: data <= 19'h7fe9e; 
        10'b1100001100: data <= 19'h7ff5c; 
        10'b1100001101: data <= 19'h00042; 
        10'b1100001110: data <= 19'h7fe57; 
        10'b1100001111: data <= 19'h7ff60; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 14) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 20'hffe34; 
        10'b0000000001: data <= 20'hffe91; 
        10'b0000000010: data <= 20'hffe43; 
        10'b0000000011: data <= 20'hfff2c; 
        10'b0000000100: data <= 20'hffef4; 
        10'b0000000101: data <= 20'h0005c; 
        10'b0000000110: data <= 20'hffc55; 
        10'b0000000111: data <= 20'hfff36; 
        10'b0000001000: data <= 20'hffd88; 
        10'b0000001001: data <= 20'hffde8; 
        10'b0000001010: data <= 20'hffd0d; 
        10'b0000001011: data <= 20'h0004e; 
        10'b0000001100: data <= 20'hffed4; 
        10'b0000001101: data <= 20'hfffcd; 
        10'b0000001110: data <= 20'hffcf1; 
        10'b0000001111: data <= 20'hfffd6; 
        10'b0000010000: data <= 20'hfff0e; 
        10'b0000010001: data <= 20'hffcb5; 
        10'b0000010010: data <= 20'h00054; 
        10'b0000010011: data <= 20'hffe8e; 
        10'b0000010100: data <= 20'hffe45; 
        10'b0000010101: data <= 20'hffe29; 
        10'b0000010110: data <= 20'hffe6c; 
        10'b0000010111: data <= 20'h000ae; 
        10'b0000011000: data <= 20'h00004; 
        10'b0000011001: data <= 20'hffde5; 
        10'b0000011010: data <= 20'hffd60; 
        10'b0000011011: data <= 20'hffe5a; 
        10'b0000011100: data <= 20'hffe44; 
        10'b0000011101: data <= 20'hffc59; 
        10'b0000011110: data <= 20'h0009e; 
        10'b0000011111: data <= 20'h00001; 
        10'b0000100000: data <= 20'hffcab; 
        10'b0000100001: data <= 20'hffcc4; 
        10'b0000100010: data <= 20'hffc77; 
        10'b0000100011: data <= 20'hffcc6; 
        10'b0000100100: data <= 20'h00074; 
        10'b0000100101: data <= 20'hffea6; 
        10'b0000100110: data <= 20'hffe81; 
        10'b0000100111: data <= 20'hffc5e; 
        10'b0000101000: data <= 20'h00066; 
        10'b0000101001: data <= 20'hfff6c; 
        10'b0000101010: data <= 20'hffd86; 
        10'b0000101011: data <= 20'hffe1f; 
        10'b0000101100: data <= 20'hfff70; 
        10'b0000101101: data <= 20'hffed3; 
        10'b0000101110: data <= 20'hffd2f; 
        10'b0000101111: data <= 20'hffeed; 
        10'b0000110000: data <= 20'h00059; 
        10'b0000110001: data <= 20'hffc97; 
        10'b0000110010: data <= 20'hfff63; 
        10'b0000110011: data <= 20'hffd37; 
        10'b0000110100: data <= 20'hfffbd; 
        10'b0000110101: data <= 20'h000c1; 
        10'b0000110110: data <= 20'hffd86; 
        10'b0000110111: data <= 20'hffd32; 
        10'b0000111000: data <= 20'hffcf2; 
        10'b0000111001: data <= 20'hffff1; 
        10'b0000111010: data <= 20'hffec7; 
        10'b0000111011: data <= 20'hffe7b; 
        10'b0000111100: data <= 20'hffd16; 
        10'b0000111101: data <= 20'hffc6a; 
        10'b0000111110: data <= 20'hffecc; 
        10'b0000111111: data <= 20'hffc50; 
        10'b0001000000: data <= 20'h000a8; 
        10'b0001000001: data <= 20'hffc4d; 
        10'b0001000010: data <= 20'hffc79; 
        10'b0001000011: data <= 20'hfff47; 
        10'b0001000100: data <= 20'hffec3; 
        10'b0001000101: data <= 20'hffc37; 
        10'b0001000110: data <= 20'hfff3d; 
        10'b0001000111: data <= 20'hffefc; 
        10'b0001001000: data <= 20'hffbfc; 
        10'b0001001001: data <= 20'hffda3; 
        10'b0001001010: data <= 20'hffda7; 
        10'b0001001011: data <= 20'hfff7f; 
        10'b0001001100: data <= 20'hfffe1; 
        10'b0001001101: data <= 20'hfffd0; 
        10'b0001001110: data <= 20'hfff1d; 
        10'b0001001111: data <= 20'hffe60; 
        10'b0001010000: data <= 20'h00059; 
        10'b0001010001: data <= 20'hffd84; 
        10'b0001010010: data <= 20'hfff70; 
        10'b0001010011: data <= 20'h00078; 
        10'b0001010100: data <= 20'hffd42; 
        10'b0001010101: data <= 20'hffe6b; 
        10'b0001010110: data <= 20'hffe73; 
        10'b0001010111: data <= 20'hffcd1; 
        10'b0001011000: data <= 20'h000a4; 
        10'b0001011001: data <= 20'hffcfe; 
        10'b0001011010: data <= 20'hffc8e; 
        10'b0001011011: data <= 20'hffded; 
        10'b0001011100: data <= 20'hffc65; 
        10'b0001011101: data <= 20'hffebe; 
        10'b0001011110: data <= 20'hffd4b; 
        10'b0001011111: data <= 20'hffaf9; 
        10'b0001100000: data <= 20'hffa69; 
        10'b0001100001: data <= 20'hff939; 
        10'b0001100010: data <= 20'hffa60; 
        10'b0001100011: data <= 20'hffcaa; 
        10'b0001100100: data <= 20'hffa5b; 
        10'b0001100101: data <= 20'hffb9e; 
        10'b0001100110: data <= 20'hffcf2; 
        10'b0001100111: data <= 20'hffe21; 
        10'b0001101000: data <= 20'hffbbb; 
        10'b0001101001: data <= 20'h00044; 
        10'b0001101010: data <= 20'hffdc4; 
        10'b0001101011: data <= 20'hfffc7; 
        10'b0001101100: data <= 20'hffd91; 
        10'b0001101101: data <= 20'hfff39; 
        10'b0001101110: data <= 20'hffedc; 
        10'b0001101111: data <= 20'hffca6; 
        10'b0001110000: data <= 20'hffe89; 
        10'b0001110001: data <= 20'hfff94; 
        10'b0001110010: data <= 20'hffde5; 
        10'b0001110011: data <= 20'hffca8; 
        10'b0001110100: data <= 20'hfffd1; 
        10'b0001110101: data <= 20'hfffbe; 
        10'b0001110110: data <= 20'hffe8b; 
        10'b0001110111: data <= 20'hffcf8; 
        10'b0001111000: data <= 20'hffcf4; 
        10'b0001111001: data <= 20'hffe36; 
        10'b0001111010: data <= 20'hffe6b; 
        10'b0001111011: data <= 20'hfff21; 
        10'b0001111100: data <= 20'h004dd; 
        10'b0001111101: data <= 20'h00324; 
        10'b0001111110: data <= 20'h00a98; 
        10'b0001111111: data <= 20'h0080a; 
        10'b0010000000: data <= 20'h003a8; 
        10'b0010000001: data <= 20'h00200; 
        10'b0010000010: data <= 20'h00300; 
        10'b0010000011: data <= 20'hffd55; 
        10'b0010000100: data <= 20'hffcc0; 
        10'b0010000101: data <= 20'hffe4f; 
        10'b0010000110: data <= 20'hffb19; 
        10'b0010000111: data <= 20'hffc7c; 
        10'b0010001000: data <= 20'hfffe3; 
        10'b0010001001: data <= 20'h0003c; 
        10'b0010001010: data <= 20'hffe1b; 
        10'b0010001011: data <= 20'hffe8b; 
        10'b0010001100: data <= 20'hffe9b; 
        10'b0010001101: data <= 20'hfff57; 
        10'b0010001110: data <= 20'hfff96; 
        10'b0010001111: data <= 20'hfffe0; 
        10'b0010010000: data <= 20'hffd1d; 
        10'b0010010001: data <= 20'hffe4b; 
        10'b0010010010: data <= 20'hffd82; 
        10'b0010010011: data <= 20'hff946; 
        10'b0010010100: data <= 20'hffd4c; 
        10'b0010010101: data <= 20'h00267; 
        10'b0010010110: data <= 20'hffa71; 
        10'b0010010111: data <= 20'h00767; 
        10'b0010011000: data <= 20'h00deb; 
        10'b0010011001: data <= 20'h00b94; 
        10'b0010011010: data <= 20'h00c0d; 
        10'b0010011011: data <= 20'h005c0; 
        10'b0010011100: data <= 20'h004bf; 
        10'b0010011101: data <= 20'h00b27; 
        10'b0010011110: data <= 20'h0008e; 
        10'b0010011111: data <= 20'hfff7e; 
        10'b0010100000: data <= 20'h003fa; 
        10'b0010100001: data <= 20'h0020f; 
        10'b0010100010: data <= 20'hff93e; 
        10'b0010100011: data <= 20'hffa54; 
        10'b0010100100: data <= 20'hffc13; 
        10'b0010100101: data <= 20'h002fe; 
        10'b0010100110: data <= 20'hffec8; 
        10'b0010100111: data <= 20'h00083; 
        10'b0010101000: data <= 20'hffd41; 
        10'b0010101001: data <= 20'hffd07; 
        10'b0010101010: data <= 20'hffc63; 
        10'b0010101011: data <= 20'hffc79; 
        10'b0010101100: data <= 20'hffbf4; 
        10'b0010101101: data <= 20'hffc0b; 
        10'b0010101110: data <= 20'hff9a4; 
        10'b0010101111: data <= 20'hff99f; 
        10'b0010110000: data <= 20'h00072; 
        10'b0010110001: data <= 20'h001e1; 
        10'b0010110010: data <= 20'hfff82; 
        10'b0010110011: data <= 20'h00395; 
        10'b0010110100: data <= 20'h005ac; 
        10'b0010110101: data <= 20'h0048b; 
        10'b0010110110: data <= 20'h00668; 
        10'b0010110111: data <= 20'h00bfd; 
        10'b0010111000: data <= 20'h005cd; 
        10'b0010111001: data <= 20'h006d3; 
        10'b0010111010: data <= 20'h00171; 
        10'b0010111011: data <= 20'h007ca; 
        10'b0010111100: data <= 20'h002f9; 
        10'b0010111101: data <= 20'h003a8; 
        10'b0010111110: data <= 20'h0048c; 
        10'b0010111111: data <= 20'h0043e; 
        10'b0011000000: data <= 20'h00395; 
        10'b0011000001: data <= 20'h00181; 
        10'b0011000010: data <= 20'hffe89; 
        10'b0011000011: data <= 20'hfffa2; 
        10'b0011000100: data <= 20'h00087; 
        10'b0011000101: data <= 20'hffd48; 
        10'b0011000110: data <= 20'hffcd0; 
        10'b0011000111: data <= 20'hffd83; 
        10'b0011001000: data <= 20'hffbc7; 
        10'b0011001001: data <= 20'hffe76; 
        10'b0011001010: data <= 20'hffbaa; 
        10'b0011001011: data <= 20'hfffbf; 
        10'b0011001100: data <= 20'h00449; 
        10'b0011001101: data <= 20'h001c1; 
        10'b0011001110: data <= 20'h00227; 
        10'b0011001111: data <= 20'hffea7; 
        10'b0011010000: data <= 20'hffa85; 
        10'b0011010001: data <= 20'hffbe4; 
        10'b0011010010: data <= 20'hff9f3; 
        10'b0011010011: data <= 20'h003a1; 
        10'b0011010100: data <= 20'h0048e; 
        10'b0011010101: data <= 20'hfffb8; 
        10'b0011010110: data <= 20'h0031a; 
        10'b0011010111: data <= 20'hffc9d; 
        10'b0011011000: data <= 20'h004a5; 
        10'b0011011001: data <= 20'h0073d; 
        10'b0011011010: data <= 20'h0014e; 
        10'b0011011011: data <= 20'h00f02; 
        10'b0011011100: data <= 20'h00932; 
        10'b0011011101: data <= 20'hfffa6; 
        10'b0011011110: data <= 20'h00038; 
        10'b0011011111: data <= 20'hfff5f; 
        10'b0011100000: data <= 20'hfff5d; 
        10'b0011100001: data <= 20'h00034; 
        10'b0011100010: data <= 20'hfff42; 
        10'b0011100011: data <= 20'hffd09; 
        10'b0011100100: data <= 20'hfff36; 
        10'b0011100101: data <= 20'hffe9b; 
        10'b0011100110: data <= 20'h00638; 
        10'b0011100111: data <= 20'h003d7; 
        10'b0011101000: data <= 20'h00163; 
        10'b0011101001: data <= 20'h00aca; 
        10'b0011101010: data <= 20'h0009e; 
        10'b0011101011: data <= 20'h0005d; 
        10'b0011101100: data <= 20'h00735; 
        10'b0011101101: data <= 20'h00956; 
        10'b0011101110: data <= 20'hff8a1; 
        10'b0011101111: data <= 20'hff9bd; 
        10'b0011110000: data <= 20'h0051b; 
        10'b0011110001: data <= 20'hffc62; 
        10'b0011110010: data <= 20'h001b3; 
        10'b0011110011: data <= 20'h004e3; 
        10'b0011110100: data <= 20'h00339; 
        10'b0011110101: data <= 20'h009f3; 
        10'b0011110110: data <= 20'h006ac; 
        10'b0011110111: data <= 20'h00b56; 
        10'b0011111000: data <= 20'h00a50; 
        10'b0011111001: data <= 20'hffec5; 
        10'b0011111010: data <= 20'hfff20; 
        10'b0011111011: data <= 20'h00105; 
        10'b0011111100: data <= 20'h00010; 
        10'b0011111101: data <= 20'h00034; 
        10'b0011111110: data <= 20'hffe63; 
        10'b0011111111: data <= 20'hffe01; 
        10'b0100000000: data <= 20'hffee9; 
        10'b0100000001: data <= 20'h0064c; 
        10'b0100000010: data <= 20'h004ac; 
        10'b0100000011: data <= 20'h009a0; 
        10'b0100000100: data <= 20'h00cea; 
        10'b0100000101: data <= 20'h00ae4; 
        10'b0100000110: data <= 20'h006e6; 
        10'b0100000111: data <= 20'h00c20; 
        10'b0100001000: data <= 20'h0034a; 
        10'b0100001001: data <= 20'h00382; 
        10'b0100001010: data <= 20'hff1d1; 
        10'b0100001011: data <= 20'hfec46; 
        10'b0100001100: data <= 20'hff91f; 
        10'b0100001101: data <= 20'h0010d; 
        10'b0100001110: data <= 20'h00223; 
        10'b0100001111: data <= 20'h003d4; 
        10'b0100010000: data <= 20'h0050f; 
        10'b0100010001: data <= 20'h0045d; 
        10'b0100010010: data <= 20'h00a6b; 
        10'b0100010011: data <= 20'h00ab4; 
        10'b0100010100: data <= 20'hffe42; 
        10'b0100010101: data <= 20'hffe88; 
        10'b0100010110: data <= 20'h00262; 
        10'b0100010111: data <= 20'hffcbb; 
        10'b0100011000: data <= 20'hffd68; 
        10'b0100011001: data <= 20'h0001b; 
        10'b0100011010: data <= 20'hffd3d; 
        10'b0100011011: data <= 20'h00046; 
        10'b0100011100: data <= 20'h0026d; 
        10'b0100011101: data <= 20'h007bd; 
        10'b0100011110: data <= 20'h007b1; 
        10'b0100011111: data <= 20'h00e19; 
        10'b0100100000: data <= 20'h00a77; 
        10'b0100100001: data <= 20'h00c3a; 
        10'b0100100010: data <= 20'h011de; 
        10'b0100100011: data <= 20'h00890; 
        10'b0100100100: data <= 20'h008f4; 
        10'b0100100101: data <= 20'h0074d; 
        10'b0100100110: data <= 20'hffda1; 
        10'b0100100111: data <= 20'hfed39; 
        10'b0100101000: data <= 20'hff09c; 
        10'b0100101001: data <= 20'hffb4f; 
        10'b0100101010: data <= 20'h0055a; 
        10'b0100101011: data <= 20'h00554; 
        10'b0100101100: data <= 20'h00577; 
        10'b0100101101: data <= 20'h00cb5; 
        10'b0100101110: data <= 20'h00e0f; 
        10'b0100101111: data <= 20'h00b79; 
        10'b0100110000: data <= 20'h00025; 
        10'b0100110001: data <= 20'hfff2a; 
        10'b0100110010: data <= 20'hffe82; 
        10'b0100110011: data <= 20'hffd86; 
        10'b0100110100: data <= 20'hffd3d; 
        10'b0100110101: data <= 20'h000a0; 
        10'b0100110110: data <= 20'hfffc0; 
        10'b0100110111: data <= 20'hffba5; 
        10'b0100111000: data <= 20'h003b1; 
        10'b0100111001: data <= 20'h0088b; 
        10'b0100111010: data <= 20'h01044; 
        10'b0100111011: data <= 20'h0151d; 
        10'b0100111100: data <= 20'h01098; 
        10'b0100111101: data <= 20'h014f8; 
        10'b0100111110: data <= 20'h00e5b; 
        10'b0100111111: data <= 20'h006c9; 
        10'b0101000000: data <= 20'h008bf; 
        10'b0101000001: data <= 20'h014e0; 
        10'b0101000010: data <= 20'h0196c; 
        10'b0101000011: data <= 20'hffce0; 
        10'b0101000100: data <= 20'hff0df; 
        10'b0101000101: data <= 20'hffacc; 
        10'b0101000110: data <= 20'hffb0c; 
        10'b0101000111: data <= 20'h00215; 
        10'b0101001000: data <= 20'h00b80; 
        10'b0101001001: data <= 20'h00dc7; 
        10'b0101001010: data <= 20'h0124c; 
        10'b0101001011: data <= 20'h01145; 
        10'b0101001100: data <= 20'h00c05; 
        10'b0101001101: data <= 20'h001f3; 
        10'b0101001110: data <= 20'h0010f; 
        10'b0101001111: data <= 20'hfff04; 
        10'b0101010000: data <= 20'hffd99; 
        10'b0101010001: data <= 20'hfff30; 
        10'b0101010010: data <= 20'hffdf9; 
        10'b0101010011: data <= 20'hfff0e; 
        10'b0101010100: data <= 20'hfff3a; 
        10'b0101010101: data <= 20'h00a37; 
        10'b0101010110: data <= 20'h00878; 
        10'b0101010111: data <= 20'h00cef; 
        10'b0101011000: data <= 20'h00c35; 
        10'b0101011001: data <= 20'h00f55; 
        10'b0101011010: data <= 20'h0029d; 
        10'b0101011011: data <= 20'h003a9; 
        10'b0101011100: data <= 20'h00207; 
        10'b0101011101: data <= 20'h01935; 
        10'b0101011110: data <= 20'h01956; 
        10'b0101011111: data <= 20'h005ae; 
        10'b0101100000: data <= 20'h000f6; 
        10'b0101100001: data <= 20'hffdc9; 
        10'b0101100010: data <= 20'hffe2d; 
        10'b0101100011: data <= 20'h00658; 
        10'b0101100100: data <= 20'h00ac8; 
        10'b0101100101: data <= 20'h01287; 
        10'b0101100110: data <= 20'h01593; 
        10'b0101100111: data <= 20'h01200; 
        10'b0101101000: data <= 20'h00b4c; 
        10'b0101101001: data <= 20'h00485; 
        10'b0101101010: data <= 20'h0023e; 
        10'b0101101011: data <= 20'hffcd1; 
        10'b0101101100: data <= 20'hffc7e; 
        10'b0101101101: data <= 20'hffebb; 
        10'b0101101110: data <= 20'h000b7; 
        10'b0101101111: data <= 20'hffcfd; 
        10'b0101110000: data <= 20'hffdb9; 
        10'b0101110001: data <= 20'hffff2; 
        10'b0101110010: data <= 20'hffe5d; 
        10'b0101110011: data <= 20'hffe75; 
        10'b0101110100: data <= 20'h00164; 
        10'b0101110101: data <= 20'hffe23; 
        10'b0101110110: data <= 20'hffa79; 
        10'b0101110111: data <= 20'h0021b; 
        10'b0101111000: data <= 20'h00943; 
        10'b0101111001: data <= 20'h0179e; 
        10'b0101111010: data <= 20'h00711; 
        10'b0101111011: data <= 20'h0115e; 
        10'b0101111100: data <= 20'h006ea; 
        10'b0101111101: data <= 20'hffb9c; 
        10'b0101111110: data <= 20'h0006a; 
        10'b0101111111: data <= 20'h00094; 
        10'b0110000000: data <= 20'h007b1; 
        10'b0110000001: data <= 20'h006fb; 
        10'b0110000010: data <= 20'h003f5; 
        10'b0110000011: data <= 20'h005a0; 
        10'b0110000100: data <= 20'h002fe; 
        10'b0110000101: data <= 20'h000aa; 
        10'b0110000110: data <= 20'h000af; 
        10'b0110000111: data <= 20'hfff6c; 
        10'b0110001000: data <= 20'hffddc; 
        10'b0110001001: data <= 20'hffc6e; 
        10'b0110001010: data <= 20'hfff84; 
        10'b0110001011: data <= 20'hffe83; 
        10'b0110001100: data <= 20'hffcd9; 
        10'b0110001101: data <= 20'hff923; 
        10'b0110001110: data <= 20'hff3c1; 
        10'b0110001111: data <= 20'hff04c; 
        10'b0110010000: data <= 20'hfed76; 
        10'b0110010001: data <= 20'hff126; 
        10'b0110010010: data <= 20'hffded; 
        10'b0110010011: data <= 20'h0097e; 
        10'b0110010100: data <= 20'h00922; 
        10'b0110010101: data <= 20'h0134e; 
        10'b0110010110: data <= 20'h00f70; 
        10'b0110010111: data <= 20'h00a70; 
        10'b0110011000: data <= 20'hffebb; 
        10'b0110011001: data <= 20'h0014c; 
        10'b0110011010: data <= 20'hffd4a; 
        10'b0110011011: data <= 20'hff9b5; 
        10'b0110011100: data <= 20'hff5c1; 
        10'b0110011101: data <= 20'hff6d5; 
        10'b0110011110: data <= 20'hff81d; 
        10'b0110011111: data <= 20'hff6ae; 
        10'b0110100000: data <= 20'hffbc7; 
        10'b0110100001: data <= 20'hfff63; 
        10'b0110100010: data <= 20'hffc3b; 
        10'b0110100011: data <= 20'h0001c; 
        10'b0110100100: data <= 20'h0004c; 
        10'b0110100101: data <= 20'hffdb6; 
        10'b0110100110: data <= 20'hffd5f; 
        10'b0110100111: data <= 20'hffee7; 
        10'b0110101000: data <= 20'hffc8d; 
        10'b0110101001: data <= 20'hff930; 
        10'b0110101010: data <= 20'hff0be; 
        10'b0110101011: data <= 20'hfed4c; 
        10'b0110101100: data <= 20'hfeef3; 
        10'b0110101101: data <= 20'hffbd7; 
        10'b0110101110: data <= 20'h000a4; 
        10'b0110101111: data <= 20'h0006b; 
        10'b0110110000: data <= 20'h00d30; 
        10'b0110110001: data <= 20'h00f97; 
        10'b0110110010: data <= 20'h00da3; 
        10'b0110110011: data <= 20'h007dd; 
        10'b0110110100: data <= 20'hffc0f; 
        10'b0110110101: data <= 20'hffc90; 
        10'b0110110110: data <= 20'hffd98; 
        10'b0110110111: data <= 20'hff231; 
        10'b0110111000: data <= 20'hfeecd; 
        10'b0110111001: data <= 20'hff2cf; 
        10'b0110111010: data <= 20'hff7a3; 
        10'b0110111011: data <= 20'hff809; 
        10'b0110111100: data <= 20'hff9fe; 
        10'b0110111101: data <= 20'hffef6; 
        10'b0110111110: data <= 20'hffbd9; 
        10'b0110111111: data <= 20'h00056; 
        10'b0111000000: data <= 20'hffe28; 
        10'b0111000001: data <= 20'hffc98; 
        10'b0111000010: data <= 20'hffda5; 
        10'b0111000011: data <= 20'hffec3; 
        10'b0111000100: data <= 20'hffa7c; 
        10'b0111000101: data <= 20'hff623; 
        10'b0111000110: data <= 20'hff026; 
        10'b0111000111: data <= 20'hff6a5; 
        10'b0111001000: data <= 20'h00649; 
        10'b0111001001: data <= 20'h006fb; 
        10'b0111001010: data <= 20'h002db; 
        10'b0111001011: data <= 20'h00666; 
        10'b0111001100: data <= 20'h00cbf; 
        10'b0111001101: data <= 20'h00b2c; 
        10'b0111001110: data <= 20'h00402; 
        10'b0111001111: data <= 20'h006aa; 
        10'b0111010000: data <= 20'h00243; 
        10'b0111010001: data <= 20'hffac8; 
        10'b0111010010: data <= 20'hff4db; 
        10'b0111010011: data <= 20'hff013; 
        10'b0111010100: data <= 20'hff013; 
        10'b0111010101: data <= 20'hfefd2; 
        10'b0111010110: data <= 20'hff305; 
        10'b0111010111: data <= 20'hffbb2; 
        10'b0111011000: data <= 20'hffa53; 
        10'b0111011001: data <= 20'hffe10; 
        10'b0111011010: data <= 20'hffdfd; 
        10'b0111011011: data <= 20'hffc80; 
        10'b0111011100: data <= 20'h000c7; 
        10'b0111011101: data <= 20'h0008a; 
        10'b0111011110: data <= 20'hffd45; 
        10'b0111011111: data <= 20'hffca8; 
        10'b0111100000: data <= 20'hffc59; 
        10'b0111100001: data <= 20'hff5cb; 
        10'b0111100010: data <= 20'hff201; 
        10'b0111100011: data <= 20'h00279; 
        10'b0111100100: data <= 20'h00d02; 
        10'b0111100101: data <= 20'h0101e; 
        10'b0111100110: data <= 20'h00529; 
        10'b0111100111: data <= 20'h00c32; 
        10'b0111101000: data <= 20'h013d9; 
        10'b0111101001: data <= 20'h00c0a; 
        10'b0111101010: data <= 20'h00105; 
        10'b0111101011: data <= 20'hffcc7; 
        10'b0111101100: data <= 20'h00171; 
        10'b0111101101: data <= 20'hff9d2; 
        10'b0111101110: data <= 20'hfefa2; 
        10'b0111101111: data <= 20'hff840; 
        10'b0111110000: data <= 20'hff84e; 
        10'b0111110001: data <= 20'hff521; 
        10'b0111110010: data <= 20'hff7f2; 
        10'b0111110011: data <= 20'hffaee; 
        10'b0111110100: data <= 20'hffd1c; 
        10'b0111110101: data <= 20'hffbe0; 
        10'b0111110110: data <= 20'hfff51; 
        10'b0111110111: data <= 20'hffddd; 
        10'b0111111000: data <= 20'hffd86; 
        10'b0111111001: data <= 20'h00028; 
        10'b0111111010: data <= 20'hffc76; 
        10'b0111111011: data <= 20'hffb76; 
        10'b0111111100: data <= 20'hff9c7; 
        10'b0111111101: data <= 20'hff99f; 
        10'b0111111110: data <= 20'hffc0e; 
        10'b0111111111: data <= 20'h003d8; 
        10'b1000000000: data <= 20'h00ab2; 
        10'b1000000001: data <= 20'h0134e; 
        10'b1000000010: data <= 20'h00d7d; 
        10'b1000000011: data <= 20'h01267; 
        10'b1000000100: data <= 20'h00bfc; 
        10'b1000000101: data <= 20'h006e7; 
        10'b1000000110: data <= 20'hff7a2; 
        10'b1000000111: data <= 20'hffdd7; 
        10'b1000001000: data <= 20'hffb49; 
        10'b1000001001: data <= 20'hff370; 
        10'b1000001010: data <= 20'hffcf9; 
        10'b1000001011: data <= 20'hffda2; 
        10'b1000001100: data <= 20'h000ed; 
        10'b1000001101: data <= 20'hff916; 
        10'b1000001110: data <= 20'hffef3; 
        10'b1000001111: data <= 20'hffa21; 
        10'b1000010000: data <= 20'hff804; 
        10'b1000010001: data <= 20'hffbe5; 
        10'b1000010010: data <= 20'hfff57; 
        10'b1000010011: data <= 20'h00081; 
        10'b1000010100: data <= 20'hffd94; 
        10'b1000010101: data <= 20'hffecd; 
        10'b1000010110: data <= 20'hfff19; 
        10'b1000010111: data <= 20'hffa97; 
        10'b1000011000: data <= 20'hff919; 
        10'b1000011001: data <= 20'hffd38; 
        10'b1000011010: data <= 20'h001d8; 
        10'b1000011011: data <= 20'h0051a; 
        10'b1000011100: data <= 20'h0054f; 
        10'b1000011101: data <= 20'h00d13; 
        10'b1000011110: data <= 20'h006b7; 
        10'b1000011111: data <= 20'hfff13; 
        10'b1000100000: data <= 20'h00331; 
        10'b1000100001: data <= 20'hff73f; 
        10'b1000100010: data <= 20'hff5c0; 
        10'b1000100011: data <= 20'hffc15; 
        10'b1000100100: data <= 20'hffcc9; 
        10'b1000100101: data <= 20'hffbcd; 
        10'b1000100110: data <= 20'h00339; 
        10'b1000100111: data <= 20'h000ed; 
        10'b1000101000: data <= 20'h00426; 
        10'b1000101001: data <= 20'h00059; 
        10'b1000101010: data <= 20'h002b1; 
        10'b1000101011: data <= 20'hffdb5; 
        10'b1000101100: data <= 20'hff9e9; 
        10'b1000101101: data <= 20'hffc5c; 
        10'b1000101110: data <= 20'hffce7; 
        10'b1000101111: data <= 20'h0005f; 
        10'b1000110000: data <= 20'hffd06; 
        10'b1000110001: data <= 20'hfff5b; 
        10'b1000110010: data <= 20'hffd46; 
        10'b1000110011: data <= 20'hffc07; 
        10'b1000110100: data <= 20'hff807; 
        10'b1000110101: data <= 20'hffea8; 
        10'b1000110110: data <= 20'h00145; 
        10'b1000110111: data <= 20'h00b50; 
        10'b1000111000: data <= 20'h0035f; 
        10'b1000111001: data <= 20'hffe8a; 
        10'b1000111010: data <= 20'hfffef; 
        10'b1000111011: data <= 20'hff670; 
        10'b1000111100: data <= 20'h0009b; 
        10'b1000111101: data <= 20'hfffc0; 
        10'b1000111110: data <= 20'hff6ec; 
        10'b1000111111: data <= 20'hffe59; 
        10'b1001000000: data <= 20'hff566; 
        10'b1001000001: data <= 20'hffca5; 
        10'b1001000010: data <= 20'h001e0; 
        10'b1001000011: data <= 20'h00129; 
        10'b1001000100: data <= 20'h0035b; 
        10'b1001000101: data <= 20'h005b2; 
        10'b1001000110: data <= 20'h005ae; 
        10'b1001000111: data <= 20'hffe99; 
        10'b1001001000: data <= 20'hffc43; 
        10'b1001001001: data <= 20'hffb16; 
        10'b1001001010: data <= 20'hffe8b; 
        10'b1001001011: data <= 20'hffd22; 
        10'b1001001100: data <= 20'h00042; 
        10'b1001001101: data <= 20'hffe6a; 
        10'b1001001110: data <= 20'h0008f; 
        10'b1001001111: data <= 20'hff9bd; 
        10'b1001010000: data <= 20'hff6b3; 
        10'b1001010001: data <= 20'hfff13; 
        10'b1001010010: data <= 20'h004e6; 
        10'b1001010011: data <= 20'h00a77; 
        10'b1001010100: data <= 20'h00231; 
        10'b1001010101: data <= 20'h0047c; 
        10'b1001010110: data <= 20'hfff2d; 
        10'b1001010111: data <= 20'hff917; 
        10'b1001011000: data <= 20'hffc22; 
        10'b1001011001: data <= 20'h00262; 
        10'b1001011010: data <= 20'hfffc9; 
        10'b1001011011: data <= 20'hffee8; 
        10'b1001011100: data <= 20'hff7e2; 
        10'b1001011101: data <= 20'hffc98; 
        10'b1001011110: data <= 20'hffdbd; 
        10'b1001011111: data <= 20'hfffad; 
        10'b1001100000: data <= 20'hfffcf; 
        10'b1001100001: data <= 20'h001f2; 
        10'b1001100010: data <= 20'h001af; 
        10'b1001100011: data <= 20'hffd8f; 
        10'b1001100100: data <= 20'hffd0f; 
        10'b1001100101: data <= 20'hfffd1; 
        10'b1001100110: data <= 20'hfff64; 
        10'b1001100111: data <= 20'hffe1e; 
        10'b1001101000: data <= 20'hfff0e; 
        10'b1001101001: data <= 20'hffc72; 
        10'b1001101010: data <= 20'hffdba; 
        10'b1001101011: data <= 20'hffc05; 
        10'b1001101100: data <= 20'hff895; 
        10'b1001101101: data <= 20'hff4ef; 
        10'b1001101110: data <= 20'h00150; 
        10'b1001101111: data <= 20'h002fb; 
        10'b1001110000: data <= 20'hfff52; 
        10'b1001110001: data <= 20'hffc76; 
        10'b1001110010: data <= 20'h0023e; 
        10'b1001110011: data <= 20'h000cc; 
        10'b1001110100: data <= 20'h00d38; 
        10'b1001110101: data <= 20'h00ddc; 
        10'b1001110110: data <= 20'h009cc; 
        10'b1001110111: data <= 20'h007a8; 
        10'b1001111000: data <= 20'hfff58; 
        10'b1001111001: data <= 20'hfff47; 
        10'b1001111010: data <= 20'h0034f; 
        10'b1001111011: data <= 20'hffbe2; 
        10'b1001111100: data <= 20'hffb8c; 
        10'b1001111101: data <= 20'h001e5; 
        10'b1001111110: data <= 20'hfff34; 
        10'b1001111111: data <= 20'hffd2a; 
        10'b1010000000: data <= 20'hfff4a; 
        10'b1010000001: data <= 20'hfff45; 
        10'b1010000010: data <= 20'hfff2d; 
        10'b1010000011: data <= 20'hffd42; 
        10'b1010000100: data <= 20'hffd39; 
        10'b1010000101: data <= 20'hfffa6; 
        10'b1010000110: data <= 20'hffebe; 
        10'b1010000111: data <= 20'hffc75; 
        10'b1010001000: data <= 20'hff83d; 
        10'b1010001001: data <= 20'hfed7d; 
        10'b1010001010: data <= 20'hff17c; 
        10'b1010001011: data <= 20'hff8b1; 
        10'b1010001100: data <= 20'h00286; 
        10'b1010001101: data <= 20'h0027e; 
        10'b1010001110: data <= 20'h0055e; 
        10'b1010001111: data <= 20'h00702; 
        10'b1010010000: data <= 20'h00fa6; 
        10'b1010010001: data <= 20'h01680; 
        10'b1010010010: data <= 20'h01327; 
        10'b1010010011: data <= 20'h00f44; 
        10'b1010010100: data <= 20'h00c5d; 
        10'b1010010101: data <= 20'h008db; 
        10'b1010010110: data <= 20'h00708; 
        10'b1010010111: data <= 20'h008fe; 
        10'b1010011000: data <= 20'h006a2; 
        10'b1010011001: data <= 20'h00198; 
        10'b1010011010: data <= 20'hfff29; 
        10'b1010011011: data <= 20'hffde8; 
        10'b1010011100: data <= 20'hffbe9; 
        10'b1010011101: data <= 20'hfff9d; 
        10'b1010011110: data <= 20'hffc60; 
        10'b1010011111: data <= 20'hfff48; 
        10'b1010100000: data <= 20'hfff8e; 
        10'b1010100001: data <= 20'hfff49; 
        10'b1010100010: data <= 20'h000b0; 
        10'b1010100011: data <= 20'hffcd2; 
        10'b1010100100: data <= 20'hffcc8; 
        10'b1010100101: data <= 20'hff3c1; 
        10'b1010100110: data <= 20'hfef01; 
        10'b1010100111: data <= 20'hff1bb; 
        10'b1010101000: data <= 20'hfff1f; 
        10'b1010101001: data <= 20'h00356; 
        10'b1010101010: data <= 20'hffebc; 
        10'b1010101011: data <= 20'h00610; 
        10'b1010101100: data <= 20'h00477; 
        10'b1010101101: data <= 20'h002f2; 
        10'b1010101110: data <= 20'h0076b; 
        10'b1010101111: data <= 20'h0101f; 
        10'b1010110000: data <= 20'h0111e; 
        10'b1010110001: data <= 20'h00b7f; 
        10'b1010110010: data <= 20'h01019; 
        10'b1010110011: data <= 20'h00f1c; 
        10'b1010110100: data <= 20'h004fb; 
        10'b1010110101: data <= 20'h00049; 
        10'b1010110110: data <= 20'hffc95; 
        10'b1010110111: data <= 20'h00059; 
        10'b1010111000: data <= 20'hffe99; 
        10'b1010111001: data <= 20'hffda6; 
        10'b1010111010: data <= 20'h0008e; 
        10'b1010111011: data <= 20'hfff10; 
        10'b1010111100: data <= 20'h000bf; 
        10'b1010111101: data <= 20'hfff76; 
        10'b1010111110: data <= 20'h0005c; 
        10'b1010111111: data <= 20'hffcca; 
        10'b1011000000: data <= 20'hffd92; 
        10'b1011000001: data <= 20'hffb74; 
        10'b1011000010: data <= 20'hff996; 
        10'b1011000011: data <= 20'hff807; 
        10'b1011000100: data <= 20'hff71c; 
        10'b1011000101: data <= 20'hff715; 
        10'b1011000110: data <= 20'hffcaa; 
        10'b1011000111: data <= 20'hff9b2; 
        10'b1011001000: data <= 20'hffc44; 
        10'b1011001001: data <= 20'hffc35; 
        10'b1011001010: data <= 20'hfff9f; 
        10'b1011001011: data <= 20'h005aa; 
        10'b1011001100: data <= 20'h00409; 
        10'b1011001101: data <= 20'h0051f; 
        10'b1011001110: data <= 20'h005d7; 
        10'b1011001111: data <= 20'h000ec; 
        10'b1011010000: data <= 20'hffec2; 
        10'b1011010001: data <= 20'hfffd7; 
        10'b1011010010: data <= 20'hffc22; 
        10'b1011010011: data <= 20'hffc49; 
        10'b1011010100: data <= 20'hfffaf; 
        10'b1011010101: data <= 20'hffef8; 
        10'b1011010110: data <= 20'hffd9b; 
        10'b1011010111: data <= 20'hffee4; 
        10'b1011011000: data <= 20'hfff67; 
        10'b1011011001: data <= 20'h00016; 
        10'b1011011010: data <= 20'hffe39; 
        10'b1011011011: data <= 20'hffd68; 
        10'b1011011100: data <= 20'hffc38; 
        10'b1011011101: data <= 20'hffcd4; 
        10'b1011011110: data <= 20'hffb24; 
        10'b1011011111: data <= 20'hffea1; 
        10'b1011100000: data <= 20'hffb9a; 
        10'b1011100001: data <= 20'hffc40; 
        10'b1011100010: data <= 20'hffb79; 
        10'b1011100011: data <= 20'hffd6a; 
        10'b1011100100: data <= 20'hffd26; 
        10'b1011100101: data <= 20'hffd92; 
        10'b1011100110: data <= 20'hffc68; 
        10'b1011100111: data <= 20'hffd66; 
        10'b1011101000: data <= 20'hffcdc; 
        10'b1011101001: data <= 20'hffbd4; 
        10'b1011101010: data <= 20'hffb59; 
        10'b1011101011: data <= 20'hffd13; 
        10'b1011101100: data <= 20'hffdf9; 
        10'b1011101101: data <= 20'hfff5e; 
        10'b1011101110: data <= 20'hffe2c; 
        10'b1011101111: data <= 20'h000d4; 
        10'b1011110000: data <= 20'h000c1; 
        10'b1011110001: data <= 20'hffc81; 
        10'b1011110010: data <= 20'hffee4; 
        10'b1011110011: data <= 20'hffe86; 
        10'b1011110100: data <= 20'hfff35; 
        10'b1011110101: data <= 20'hffd4f; 
        10'b1011110110: data <= 20'hffe51; 
        10'b1011110111: data <= 20'hffeef; 
        10'b1011111000: data <= 20'hfff15; 
        10'b1011111001: data <= 20'hffc69; 
        10'b1011111010: data <= 20'hfffdf; 
        10'b1011111011: data <= 20'hffd95; 
        10'b1011111100: data <= 20'h00097; 
        10'b1011111101: data <= 20'hffe3a; 
        10'b1011111110: data <= 20'hffce7; 
        10'b1011111111: data <= 20'hfffac; 
        10'b1100000000: data <= 20'hffd7a; 
        10'b1100000001: data <= 20'hffcf5; 
        10'b1100000010: data <= 20'hffe1b; 
        10'b1100000011: data <= 20'hfff30; 
        10'b1100000100: data <= 20'hffedf; 
        10'b1100000101: data <= 20'h00010; 
        10'b1100000110: data <= 20'h0007f; 
        10'b1100000111: data <= 20'h000b4; 
        10'b1100001000: data <= 20'hfff66; 
        10'b1100001001: data <= 20'hffefb; 
        10'b1100001010: data <= 20'hfff5b; 
        10'b1100001011: data <= 20'hffd3c; 
        10'b1100001100: data <= 20'hffeb8; 
        10'b1100001101: data <= 20'h00085; 
        10'b1100001110: data <= 20'hffcaf; 
        10'b1100001111: data <= 20'hffebf; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 15) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 21'h1ffc68; 
        10'b0000000001: data <= 21'h1ffd22; 
        10'b0000000010: data <= 21'h1ffc86; 
        10'b0000000011: data <= 21'h1ffe58; 
        10'b0000000100: data <= 21'h1ffde7; 
        10'b0000000101: data <= 21'h0000b7; 
        10'b0000000110: data <= 21'h1ff8a9; 
        10'b0000000111: data <= 21'h1ffe6d; 
        10'b0000001000: data <= 21'h1ffb10; 
        10'b0000001001: data <= 21'h1ffbd1; 
        10'b0000001010: data <= 21'h1ffa1a; 
        10'b0000001011: data <= 21'h00009d; 
        10'b0000001100: data <= 21'h1ffda8; 
        10'b0000001101: data <= 21'h1fff9b; 
        10'b0000001110: data <= 21'h1ff9e2; 
        10'b0000001111: data <= 21'h1fffab; 
        10'b0000010000: data <= 21'h1ffe1c; 
        10'b0000010001: data <= 21'h1ff96a; 
        10'b0000010010: data <= 21'h0000a8; 
        10'b0000010011: data <= 21'h1ffd1b; 
        10'b0000010100: data <= 21'h1ffc8a; 
        10'b0000010101: data <= 21'h1ffc53; 
        10'b0000010110: data <= 21'h1ffcd7; 
        10'b0000010111: data <= 21'h00015c; 
        10'b0000011000: data <= 21'h000009; 
        10'b0000011001: data <= 21'h1ffbca; 
        10'b0000011010: data <= 21'h1ffac1; 
        10'b0000011011: data <= 21'h1ffcb4; 
        10'b0000011100: data <= 21'h1ffc88; 
        10'b0000011101: data <= 21'h1ff8b1; 
        10'b0000011110: data <= 21'h00013b; 
        10'b0000011111: data <= 21'h000002; 
        10'b0000100000: data <= 21'h1ff956; 
        10'b0000100001: data <= 21'h1ff988; 
        10'b0000100010: data <= 21'h1ff8ef; 
        10'b0000100011: data <= 21'h1ff98c; 
        10'b0000100100: data <= 21'h0000e9; 
        10'b0000100101: data <= 21'h1ffd4c; 
        10'b0000100110: data <= 21'h1ffd03; 
        10'b0000100111: data <= 21'h1ff8bd; 
        10'b0000101000: data <= 21'h0000cc; 
        10'b0000101001: data <= 21'h1ffed8; 
        10'b0000101010: data <= 21'h1ffb0c; 
        10'b0000101011: data <= 21'h1ffc3e; 
        10'b0000101100: data <= 21'h1ffee0; 
        10'b0000101101: data <= 21'h1ffda5; 
        10'b0000101110: data <= 21'h1ffa5e; 
        10'b0000101111: data <= 21'h1ffddb; 
        10'b0000110000: data <= 21'h0000b3; 
        10'b0000110001: data <= 21'h1ff92d; 
        10'b0000110010: data <= 21'h1ffec7; 
        10'b0000110011: data <= 21'h1ffa6e; 
        10'b0000110100: data <= 21'h1fff79; 
        10'b0000110101: data <= 21'h000183; 
        10'b0000110110: data <= 21'h1ffb0c; 
        10'b0000110111: data <= 21'h1ffa63; 
        10'b0000111000: data <= 21'h1ff9e4; 
        10'b0000111001: data <= 21'h1fffe3; 
        10'b0000111010: data <= 21'h1ffd8e; 
        10'b0000111011: data <= 21'h1ffcf6; 
        10'b0000111100: data <= 21'h1ffa2c; 
        10'b0000111101: data <= 21'h1ff8d5; 
        10'b0000111110: data <= 21'h1ffd98; 
        10'b0000111111: data <= 21'h1ff8a1; 
        10'b0001000000: data <= 21'h00014f; 
        10'b0001000001: data <= 21'h1ff89a; 
        10'b0001000010: data <= 21'h1ff8f2; 
        10'b0001000011: data <= 21'h1ffe8d; 
        10'b0001000100: data <= 21'h1ffd87; 
        10'b0001000101: data <= 21'h1ff86e; 
        10'b0001000110: data <= 21'h1ffe7a; 
        10'b0001000111: data <= 21'h1ffdf7; 
        10'b0001001000: data <= 21'h1ff7f9; 
        10'b0001001001: data <= 21'h1ffb46; 
        10'b0001001010: data <= 21'h1ffb4e; 
        10'b0001001011: data <= 21'h1ffeff; 
        10'b0001001100: data <= 21'h1fffc3; 
        10'b0001001101: data <= 21'h1fff9f; 
        10'b0001001110: data <= 21'h1ffe3a; 
        10'b0001001111: data <= 21'h1ffcc0; 
        10'b0001010000: data <= 21'h0000b2; 
        10'b0001010001: data <= 21'h1ffb08; 
        10'b0001010010: data <= 21'h1ffedf; 
        10'b0001010011: data <= 21'h0000f1; 
        10'b0001010100: data <= 21'h1ffa85; 
        10'b0001010101: data <= 21'h1ffcd6; 
        10'b0001010110: data <= 21'h1ffce7; 
        10'b0001010111: data <= 21'h1ff9a3; 
        10'b0001011000: data <= 21'h000148; 
        10'b0001011001: data <= 21'h1ff9fd; 
        10'b0001011010: data <= 21'h1ff91d; 
        10'b0001011011: data <= 21'h1ffbda; 
        10'b0001011100: data <= 21'h1ff8ca; 
        10'b0001011101: data <= 21'h1ffd7d; 
        10'b0001011110: data <= 21'h1ffa95; 
        10'b0001011111: data <= 21'h1ff5f2; 
        10'b0001100000: data <= 21'h1ff4d1; 
        10'b0001100001: data <= 21'h1ff271; 
        10'b0001100010: data <= 21'h1ff4c0; 
        10'b0001100011: data <= 21'h1ff954; 
        10'b0001100100: data <= 21'h1ff4b6; 
        10'b0001100101: data <= 21'h1ff73c; 
        10'b0001100110: data <= 21'h1ff9e4; 
        10'b0001100111: data <= 21'h1ffc41; 
        10'b0001101000: data <= 21'h1ff776; 
        10'b0001101001: data <= 21'h000088; 
        10'b0001101010: data <= 21'h1ffb87; 
        10'b0001101011: data <= 21'h1fff8e; 
        10'b0001101100: data <= 21'h1ffb21; 
        10'b0001101101: data <= 21'h1ffe71; 
        10'b0001101110: data <= 21'h1ffdb8; 
        10'b0001101111: data <= 21'h1ff94c; 
        10'b0001110000: data <= 21'h1ffd12; 
        10'b0001110001: data <= 21'h1fff28; 
        10'b0001110010: data <= 21'h1ffbca; 
        10'b0001110011: data <= 21'h1ff950; 
        10'b0001110100: data <= 21'h1fffa2; 
        10'b0001110101: data <= 21'h1fff7d; 
        10'b0001110110: data <= 21'h1ffd16; 
        10'b0001110111: data <= 21'h1ff9ef; 
        10'b0001111000: data <= 21'h1ff9e8; 
        10'b0001111001: data <= 21'h1ffc6c; 
        10'b0001111010: data <= 21'h1ffcd6; 
        10'b0001111011: data <= 21'h1ffe41; 
        10'b0001111100: data <= 21'h0009bb; 
        10'b0001111101: data <= 21'h000648; 
        10'b0001111110: data <= 21'h001531; 
        10'b0001111111: data <= 21'h001014; 
        10'b0010000000: data <= 21'h00074f; 
        10'b0010000001: data <= 21'h000400; 
        10'b0010000010: data <= 21'h000600; 
        10'b0010000011: data <= 21'h1ffaaa; 
        10'b0010000100: data <= 21'h1ff980; 
        10'b0010000101: data <= 21'h1ffc9f; 
        10'b0010000110: data <= 21'h1ff632; 
        10'b0010000111: data <= 21'h1ff8f9; 
        10'b0010001000: data <= 21'h1fffc7; 
        10'b0010001001: data <= 21'h000078; 
        10'b0010001010: data <= 21'h1ffc36; 
        10'b0010001011: data <= 21'h1ffd15; 
        10'b0010001100: data <= 21'h1ffd36; 
        10'b0010001101: data <= 21'h1ffeaf; 
        10'b0010001110: data <= 21'h1fff2c; 
        10'b0010001111: data <= 21'h1fffc0; 
        10'b0010010000: data <= 21'h1ffa39; 
        10'b0010010001: data <= 21'h1ffc96; 
        10'b0010010010: data <= 21'h1ffb04; 
        10'b0010010011: data <= 21'h1ff28b; 
        10'b0010010100: data <= 21'h1ffa98; 
        10'b0010010101: data <= 21'h0004ce; 
        10'b0010010110: data <= 21'h1ff4e2; 
        10'b0010010111: data <= 21'h000ece; 
        10'b0010011000: data <= 21'h001bd6; 
        10'b0010011001: data <= 21'h001729; 
        10'b0010011010: data <= 21'h00181a; 
        10'b0010011011: data <= 21'h000b80; 
        10'b0010011100: data <= 21'h00097d; 
        10'b0010011101: data <= 21'h00164d; 
        10'b0010011110: data <= 21'h00011d; 
        10'b0010011111: data <= 21'h1ffefc; 
        10'b0010100000: data <= 21'h0007f5; 
        10'b0010100001: data <= 21'h00041e; 
        10'b0010100010: data <= 21'h1ff27c; 
        10'b0010100011: data <= 21'h1ff4a8; 
        10'b0010100100: data <= 21'h1ff826; 
        10'b0010100101: data <= 21'h0005fc; 
        10'b0010100110: data <= 21'h1ffd8f; 
        10'b0010100111: data <= 21'h000107; 
        10'b0010101000: data <= 21'h1ffa82; 
        10'b0010101001: data <= 21'h1ffa0e; 
        10'b0010101010: data <= 21'h1ff8c6; 
        10'b0010101011: data <= 21'h1ff8f2; 
        10'b0010101100: data <= 21'h1ff7e8; 
        10'b0010101101: data <= 21'h1ff816; 
        10'b0010101110: data <= 21'h1ff349; 
        10'b0010101111: data <= 21'h1ff33d; 
        10'b0010110000: data <= 21'h0000e4; 
        10'b0010110001: data <= 21'h0003c2; 
        10'b0010110010: data <= 21'h1fff04; 
        10'b0010110011: data <= 21'h00072a; 
        10'b0010110100: data <= 21'h000b57; 
        10'b0010110101: data <= 21'h000917; 
        10'b0010110110: data <= 21'h000cd0; 
        10'b0010110111: data <= 21'h0017fa; 
        10'b0010111000: data <= 21'h000b9b; 
        10'b0010111001: data <= 21'h000da5; 
        10'b0010111010: data <= 21'h0002e1; 
        10'b0010111011: data <= 21'h000f93; 
        10'b0010111100: data <= 21'h0005f2; 
        10'b0010111101: data <= 21'h000750; 
        10'b0010111110: data <= 21'h000918; 
        10'b0010111111: data <= 21'h00087d; 
        10'b0011000000: data <= 21'h00072a; 
        10'b0011000001: data <= 21'h000303; 
        10'b0011000010: data <= 21'h1ffd13; 
        10'b0011000011: data <= 21'h1fff45; 
        10'b0011000100: data <= 21'h00010e; 
        10'b0011000101: data <= 21'h1ffa91; 
        10'b0011000110: data <= 21'h1ff99f; 
        10'b0011000111: data <= 21'h1ffb07; 
        10'b0011001000: data <= 21'h1ff78e; 
        10'b0011001001: data <= 21'h1ffcec; 
        10'b0011001010: data <= 21'h1ff754; 
        10'b0011001011: data <= 21'h1fff7d; 
        10'b0011001100: data <= 21'h000892; 
        10'b0011001101: data <= 21'h000381; 
        10'b0011001110: data <= 21'h00044f; 
        10'b0011001111: data <= 21'h1ffd4d; 
        10'b0011010000: data <= 21'h1ff50a; 
        10'b0011010001: data <= 21'h1ff7c9; 
        10'b0011010010: data <= 21'h1ff3e6; 
        10'b0011010011: data <= 21'h000742; 
        10'b0011010100: data <= 21'h00091c; 
        10'b0011010101: data <= 21'h1fff70; 
        10'b0011010110: data <= 21'h000634; 
        10'b0011010111: data <= 21'h1ff939; 
        10'b0011011000: data <= 21'h00094a; 
        10'b0011011001: data <= 21'h000e7b; 
        10'b0011011010: data <= 21'h00029b; 
        10'b0011011011: data <= 21'h001e04; 
        10'b0011011100: data <= 21'h001263; 
        10'b0011011101: data <= 21'h1fff4c; 
        10'b0011011110: data <= 21'h000071; 
        10'b0011011111: data <= 21'h1ffebd; 
        10'b0011100000: data <= 21'h1ffeb9; 
        10'b0011100001: data <= 21'h000067; 
        10'b0011100010: data <= 21'h1ffe84; 
        10'b0011100011: data <= 21'h1ffa13; 
        10'b0011100100: data <= 21'h1ffe6d; 
        10'b0011100101: data <= 21'h1ffd36; 
        10'b0011100110: data <= 21'h000c70; 
        10'b0011100111: data <= 21'h0007af; 
        10'b0011101000: data <= 21'h0002c6; 
        10'b0011101001: data <= 21'h001593; 
        10'b0011101010: data <= 21'h00013c; 
        10'b0011101011: data <= 21'h0000ba; 
        10'b0011101100: data <= 21'h000e6a; 
        10'b0011101101: data <= 21'h0012ac; 
        10'b0011101110: data <= 21'h1ff143; 
        10'b0011101111: data <= 21'h1ff37a; 
        10'b0011110000: data <= 21'h000a35; 
        10'b0011110001: data <= 21'h1ff8c4; 
        10'b0011110010: data <= 21'h000365; 
        10'b0011110011: data <= 21'h0009c6; 
        10'b0011110100: data <= 21'h000673; 
        10'b0011110101: data <= 21'h0013e6; 
        10'b0011110110: data <= 21'h000d57; 
        10'b0011110111: data <= 21'h0016ad; 
        10'b0011111000: data <= 21'h0014a1; 
        10'b0011111001: data <= 21'h1ffd8b; 
        10'b0011111010: data <= 21'h1ffe3f; 
        10'b0011111011: data <= 21'h00020a; 
        10'b0011111100: data <= 21'h00001f; 
        10'b0011111101: data <= 21'h000068; 
        10'b0011111110: data <= 21'h1ffcc5; 
        10'b0011111111: data <= 21'h1ffc03; 
        10'b0100000000: data <= 21'h1ffdd3; 
        10'b0100000001: data <= 21'h000c99; 
        10'b0100000010: data <= 21'h000959; 
        10'b0100000011: data <= 21'h001341; 
        10'b0100000100: data <= 21'h0019d4; 
        10'b0100000101: data <= 21'h0015c7; 
        10'b0100000110: data <= 21'h000dcd; 
        10'b0100000111: data <= 21'h001840; 
        10'b0100001000: data <= 21'h000694; 
        10'b0100001001: data <= 21'h000704; 
        10'b0100001010: data <= 21'h1fe3a2; 
        10'b0100001011: data <= 21'h1fd88c; 
        10'b0100001100: data <= 21'h1ff23e; 
        10'b0100001101: data <= 21'h00021a; 
        10'b0100001110: data <= 21'h000446; 
        10'b0100001111: data <= 21'h0007a8; 
        10'b0100010000: data <= 21'h000a1d; 
        10'b0100010001: data <= 21'h0008ba; 
        10'b0100010010: data <= 21'h0014d7; 
        10'b0100010011: data <= 21'h001567; 
        10'b0100010100: data <= 21'h1ffc84; 
        10'b0100010101: data <= 21'h1ffd10; 
        10'b0100010110: data <= 21'h0004c4; 
        10'b0100010111: data <= 21'h1ff976; 
        10'b0100011000: data <= 21'h1ffad0; 
        10'b0100011001: data <= 21'h000035; 
        10'b0100011010: data <= 21'h1ffa7a; 
        10'b0100011011: data <= 21'h00008d; 
        10'b0100011100: data <= 21'h0004db; 
        10'b0100011101: data <= 21'h000f7b; 
        10'b0100011110: data <= 21'h000f62; 
        10'b0100011111: data <= 21'h001c32; 
        10'b0100100000: data <= 21'h0014ed; 
        10'b0100100001: data <= 21'h001874; 
        10'b0100100010: data <= 21'h0023bc; 
        10'b0100100011: data <= 21'h001121; 
        10'b0100100100: data <= 21'h0011e7; 
        10'b0100100101: data <= 21'h000e99; 
        10'b0100100110: data <= 21'h1ffb42; 
        10'b0100100111: data <= 21'h1fda71; 
        10'b0100101000: data <= 21'h1fe139; 
        10'b0100101001: data <= 21'h1ff69e; 
        10'b0100101010: data <= 21'h000ab5; 
        10'b0100101011: data <= 21'h000aa8; 
        10'b0100101100: data <= 21'h000aed; 
        10'b0100101101: data <= 21'h00196a; 
        10'b0100101110: data <= 21'h001c1f; 
        10'b0100101111: data <= 21'h0016f1; 
        10'b0100110000: data <= 21'h00004b; 
        10'b0100110001: data <= 21'h1ffe54; 
        10'b0100110010: data <= 21'h1ffd05; 
        10'b0100110011: data <= 21'h1ffb0c; 
        10'b0100110100: data <= 21'h1ffa7a; 
        10'b0100110101: data <= 21'h000140; 
        10'b0100110110: data <= 21'h1fff80; 
        10'b0100110111: data <= 21'h1ff74a; 
        10'b0100111000: data <= 21'h000761; 
        10'b0100111001: data <= 21'h001115; 
        10'b0100111010: data <= 21'h002088; 
        10'b0100111011: data <= 21'h002a39; 
        10'b0100111100: data <= 21'h002130; 
        10'b0100111101: data <= 21'h0029f0; 
        10'b0100111110: data <= 21'h001cb7; 
        10'b0100111111: data <= 21'h000d93; 
        10'b0101000000: data <= 21'h00117d; 
        10'b0101000001: data <= 21'h0029c0; 
        10'b0101000010: data <= 21'h0032d8; 
        10'b0101000011: data <= 21'h1ff9c0; 
        10'b0101000100: data <= 21'h1fe1be; 
        10'b0101000101: data <= 21'h1ff598; 
        10'b0101000110: data <= 21'h1ff617; 
        10'b0101000111: data <= 21'h00042a; 
        10'b0101001000: data <= 21'h0016ff; 
        10'b0101001001: data <= 21'h001b8e; 
        10'b0101001010: data <= 21'h002499; 
        10'b0101001011: data <= 21'h00228b; 
        10'b0101001100: data <= 21'h00180a; 
        10'b0101001101: data <= 21'h0003e7; 
        10'b0101001110: data <= 21'h00021d; 
        10'b0101001111: data <= 21'h1ffe07; 
        10'b0101010000: data <= 21'h1ffb33; 
        10'b0101010001: data <= 21'h1ffe61; 
        10'b0101010010: data <= 21'h1ffbf1; 
        10'b0101010011: data <= 21'h1ffe1d; 
        10'b0101010100: data <= 21'h1ffe74; 
        10'b0101010101: data <= 21'h00146e; 
        10'b0101010110: data <= 21'h0010ef; 
        10'b0101010111: data <= 21'h0019de; 
        10'b0101011000: data <= 21'h001869; 
        10'b0101011001: data <= 21'h001eab; 
        10'b0101011010: data <= 21'h000539; 
        10'b0101011011: data <= 21'h000752; 
        10'b0101011100: data <= 21'h00040e; 
        10'b0101011101: data <= 21'h00326b; 
        10'b0101011110: data <= 21'h0032ab; 
        10'b0101011111: data <= 21'h000b5c; 
        10'b0101100000: data <= 21'h0001ed; 
        10'b0101100001: data <= 21'h1ffb92; 
        10'b0101100010: data <= 21'h1ffc5a; 
        10'b0101100011: data <= 21'h000cb1; 
        10'b0101100100: data <= 21'h00158f; 
        10'b0101100101: data <= 21'h00250e; 
        10'b0101100110: data <= 21'h002b26; 
        10'b0101100111: data <= 21'h0023ff; 
        10'b0101101000: data <= 21'h001698; 
        10'b0101101001: data <= 21'h00090b; 
        10'b0101101010: data <= 21'h00047b; 
        10'b0101101011: data <= 21'h1ff9a2; 
        10'b0101101100: data <= 21'h1ff8fb; 
        10'b0101101101: data <= 21'h1ffd76; 
        10'b0101101110: data <= 21'h00016e; 
        10'b0101101111: data <= 21'h1ff9fb; 
        10'b0101110000: data <= 21'h1ffb71; 
        10'b0101110001: data <= 21'h1fffe4; 
        10'b0101110010: data <= 21'h1ffcba; 
        10'b0101110011: data <= 21'h1ffcea; 
        10'b0101110100: data <= 21'h0002c8; 
        10'b0101110101: data <= 21'h1ffc46; 
        10'b0101110110: data <= 21'h1ff4f3; 
        10'b0101110111: data <= 21'h000436; 
        10'b0101111000: data <= 21'h001285; 
        10'b0101111001: data <= 21'h002f3b; 
        10'b0101111010: data <= 21'h000e22; 
        10'b0101111011: data <= 21'h0022bc; 
        10'b0101111100: data <= 21'h000dd3; 
        10'b0101111101: data <= 21'h1ff738; 
        10'b0101111110: data <= 21'h0000d3; 
        10'b0101111111: data <= 21'h000128; 
        10'b0110000000: data <= 21'h000f62; 
        10'b0110000001: data <= 21'h000df6; 
        10'b0110000010: data <= 21'h0007ea; 
        10'b0110000011: data <= 21'h000b41; 
        10'b0110000100: data <= 21'h0005fc; 
        10'b0110000101: data <= 21'h000154; 
        10'b0110000110: data <= 21'h00015d; 
        10'b0110000111: data <= 21'h1ffed7; 
        10'b0110001000: data <= 21'h1ffbb8; 
        10'b0110001001: data <= 21'h1ff8dc; 
        10'b0110001010: data <= 21'h1fff07; 
        10'b0110001011: data <= 21'h1ffd07; 
        10'b0110001100: data <= 21'h1ff9b3; 
        10'b0110001101: data <= 21'h1ff247; 
        10'b0110001110: data <= 21'h1fe781; 
        10'b0110001111: data <= 21'h1fe098; 
        10'b0110010000: data <= 21'h1fdaec; 
        10'b0110010001: data <= 21'h1fe24d; 
        10'b0110010010: data <= 21'h1ffbda; 
        10'b0110010011: data <= 21'h0012fd; 
        10'b0110010100: data <= 21'h001244; 
        10'b0110010101: data <= 21'h00269b; 
        10'b0110010110: data <= 21'h001ee0; 
        10'b0110010111: data <= 21'h0014e1; 
        10'b0110011000: data <= 21'h1ffd76; 
        10'b0110011001: data <= 21'h000299; 
        10'b0110011010: data <= 21'h1ffa94; 
        10'b0110011011: data <= 21'h1ff369; 
        10'b0110011100: data <= 21'h1feb81; 
        10'b0110011101: data <= 21'h1fedaa; 
        10'b0110011110: data <= 21'h1ff03b; 
        10'b0110011111: data <= 21'h1fed5c; 
        10'b0110100000: data <= 21'h1ff78e; 
        10'b0110100001: data <= 21'h1ffec6; 
        10'b0110100010: data <= 21'h1ff875; 
        10'b0110100011: data <= 21'h000038; 
        10'b0110100100: data <= 21'h000098; 
        10'b0110100101: data <= 21'h1ffb6c; 
        10'b0110100110: data <= 21'h1ffabe; 
        10'b0110100111: data <= 21'h1ffdce; 
        10'b0110101000: data <= 21'h1ff91a; 
        10'b0110101001: data <= 21'h1ff25f; 
        10'b0110101010: data <= 21'h1fe17b; 
        10'b0110101011: data <= 21'h1fda99; 
        10'b0110101100: data <= 21'h1fdde6; 
        10'b0110101101: data <= 21'h1ff7af; 
        10'b0110101110: data <= 21'h000149; 
        10'b0110101111: data <= 21'h0000d6; 
        10'b0110110000: data <= 21'h001a5f; 
        10'b0110110001: data <= 21'h001f2d; 
        10'b0110110010: data <= 21'h001b46; 
        10'b0110110011: data <= 21'h000fba; 
        10'b0110110100: data <= 21'h1ff81d; 
        10'b0110110101: data <= 21'h1ff921; 
        10'b0110110110: data <= 21'h1ffb2f; 
        10'b0110110111: data <= 21'h1fe462; 
        10'b0110111000: data <= 21'h1fdd9a; 
        10'b0110111001: data <= 21'h1fe59e; 
        10'b0110111010: data <= 21'h1fef46; 
        10'b0110111011: data <= 21'h1ff012; 
        10'b0110111100: data <= 21'h1ff3fc; 
        10'b0110111101: data <= 21'h1ffdec; 
        10'b0110111110: data <= 21'h1ff7b2; 
        10'b0110111111: data <= 21'h0000ad; 
        10'b0111000000: data <= 21'h1ffc50; 
        10'b0111000001: data <= 21'h1ff930; 
        10'b0111000010: data <= 21'h1ffb4a; 
        10'b0111000011: data <= 21'h1ffd86; 
        10'b0111000100: data <= 21'h1ff4f8; 
        10'b0111000101: data <= 21'h1fec47; 
        10'b0111000110: data <= 21'h1fe04d; 
        10'b0111000111: data <= 21'h1fed49; 
        10'b0111001000: data <= 21'h000c92; 
        10'b0111001001: data <= 21'h000df6; 
        10'b0111001010: data <= 21'h0005b6; 
        10'b0111001011: data <= 21'h000ccd; 
        10'b0111001100: data <= 21'h00197f; 
        10'b0111001101: data <= 21'h001658; 
        10'b0111001110: data <= 21'h000804; 
        10'b0111001111: data <= 21'h000d55; 
        10'b0111010000: data <= 21'h000485; 
        10'b0111010001: data <= 21'h1ff58f; 
        10'b0111010010: data <= 21'h1fe9b6; 
        10'b0111010011: data <= 21'h1fe026; 
        10'b0111010100: data <= 21'h1fe026; 
        10'b0111010101: data <= 21'h1fdfa3; 
        10'b0111010110: data <= 21'h1fe60b; 
        10'b0111010111: data <= 21'h1ff764; 
        10'b0111011000: data <= 21'h1ff4a7; 
        10'b0111011001: data <= 21'h1ffc1f; 
        10'b0111011010: data <= 21'h1ffbf9; 
        10'b0111011011: data <= 21'h1ff900; 
        10'b0111011100: data <= 21'h00018e; 
        10'b0111011101: data <= 21'h000114; 
        10'b0111011110: data <= 21'h1ffa8a; 
        10'b0111011111: data <= 21'h1ff950; 
        10'b0111100000: data <= 21'h1ff8b3; 
        10'b0111100001: data <= 21'h1feb95; 
        10'b0111100010: data <= 21'h1fe403; 
        10'b0111100011: data <= 21'h0004f3; 
        10'b0111100100: data <= 21'h001a04; 
        10'b0111100101: data <= 21'h00203c; 
        10'b0111100110: data <= 21'h000a51; 
        10'b0111100111: data <= 21'h001864; 
        10'b0111101000: data <= 21'h0027b2; 
        10'b0111101001: data <= 21'h001814; 
        10'b0111101010: data <= 21'h000209; 
        10'b0111101011: data <= 21'h1ff98d; 
        10'b0111101100: data <= 21'h0002e3; 
        10'b0111101101: data <= 21'h1ff3a3; 
        10'b0111101110: data <= 21'h1fdf45; 
        10'b0111101111: data <= 21'h1ff07f; 
        10'b0111110000: data <= 21'h1ff09d; 
        10'b0111110001: data <= 21'h1fea41; 
        10'b0111110010: data <= 21'h1fefe5; 
        10'b0111110011: data <= 21'h1ff5db; 
        10'b0111110100: data <= 21'h1ffa39; 
        10'b0111110101: data <= 21'h1ff7c0; 
        10'b0111110110: data <= 21'h1ffea2; 
        10'b0111110111: data <= 21'h1ffbba; 
        10'b0111111000: data <= 21'h1ffb0c; 
        10'b0111111001: data <= 21'h000050; 
        10'b0111111010: data <= 21'h1ff8ec; 
        10'b0111111011: data <= 21'h1ff6ed; 
        10'b0111111100: data <= 21'h1ff38d; 
        10'b0111111101: data <= 21'h1ff33e; 
        10'b0111111110: data <= 21'h1ff81d; 
        10'b0111111111: data <= 21'h0007b0; 
        10'b1000000000: data <= 21'h001564; 
        10'b1000000001: data <= 21'h00269b; 
        10'b1000000010: data <= 21'h001afa; 
        10'b1000000011: data <= 21'h0024ce; 
        10'b1000000100: data <= 21'h0017f7; 
        10'b1000000101: data <= 21'h000dcf; 
        10'b1000000110: data <= 21'h1fef44; 
        10'b1000000111: data <= 21'h1ffbae; 
        10'b1000001000: data <= 21'h1ff692; 
        10'b1000001001: data <= 21'h1fe6e1; 
        10'b1000001010: data <= 21'h1ff9f2; 
        10'b1000001011: data <= 21'h1ffb45; 
        10'b1000001100: data <= 21'h0001da; 
        10'b1000001101: data <= 21'h1ff22b; 
        10'b1000001110: data <= 21'h1ffde6; 
        10'b1000001111: data <= 21'h1ff441; 
        10'b1000010000: data <= 21'h1ff007; 
        10'b1000010001: data <= 21'h1ff7cb; 
        10'b1000010010: data <= 21'h1ffeaf; 
        10'b1000010011: data <= 21'h000103; 
        10'b1000010100: data <= 21'h1ffb27; 
        10'b1000010101: data <= 21'h1ffd9a; 
        10'b1000010110: data <= 21'h1ffe33; 
        10'b1000010111: data <= 21'h1ff52f; 
        10'b1000011000: data <= 21'h1ff233; 
        10'b1000011001: data <= 21'h1ffa71; 
        10'b1000011010: data <= 21'h0003af; 
        10'b1000011011: data <= 21'h000a33; 
        10'b1000011100: data <= 21'h000a9e; 
        10'b1000011101: data <= 21'h001a25; 
        10'b1000011110: data <= 21'h000d6e; 
        10'b1000011111: data <= 21'h1ffe25; 
        10'b1000100000: data <= 21'h000662; 
        10'b1000100001: data <= 21'h1fee7f; 
        10'b1000100010: data <= 21'h1feb81; 
        10'b1000100011: data <= 21'h1ff82a; 
        10'b1000100100: data <= 21'h1ff991; 
        10'b1000100101: data <= 21'h1ff79a; 
        10'b1000100110: data <= 21'h000672; 
        10'b1000100111: data <= 21'h0001da; 
        10'b1000101000: data <= 21'h00084b; 
        10'b1000101001: data <= 21'h0000b3; 
        10'b1000101010: data <= 21'h000562; 
        10'b1000101011: data <= 21'h1ffb6a; 
        10'b1000101100: data <= 21'h1ff3d1; 
        10'b1000101101: data <= 21'h1ff8b8; 
        10'b1000101110: data <= 21'h1ff9ce; 
        10'b1000101111: data <= 21'h0000bd; 
        10'b1000110000: data <= 21'h1ffa0c; 
        10'b1000110001: data <= 21'h1ffeb5; 
        10'b1000110010: data <= 21'h1ffa8c; 
        10'b1000110011: data <= 21'h1ff80e; 
        10'b1000110100: data <= 21'h1ff00e; 
        10'b1000110101: data <= 21'h1ffd50; 
        10'b1000110110: data <= 21'h00028b; 
        10'b1000110111: data <= 21'h00169f; 
        10'b1000111000: data <= 21'h0006be; 
        10'b1000111001: data <= 21'h1ffd15; 
        10'b1000111010: data <= 21'h1fffdf; 
        10'b1000111011: data <= 21'h1fecdf; 
        10'b1000111100: data <= 21'h000136; 
        10'b1000111101: data <= 21'h1fff7f; 
        10'b1000111110: data <= 21'h1fedd8; 
        10'b1000111111: data <= 21'h1ffcb3; 
        10'b1001000000: data <= 21'h1feacc; 
        10'b1001000001: data <= 21'h1ff94a; 
        10'b1001000010: data <= 21'h0003c0; 
        10'b1001000011: data <= 21'h000252; 
        10'b1001000100: data <= 21'h0006b6; 
        10'b1001000101: data <= 21'h000b65; 
        10'b1001000110: data <= 21'h000b5c; 
        10'b1001000111: data <= 21'h1ffd32; 
        10'b1001001000: data <= 21'h1ff886; 
        10'b1001001001: data <= 21'h1ff62d; 
        10'b1001001010: data <= 21'h1ffd17; 
        10'b1001001011: data <= 21'h1ffa44; 
        10'b1001001100: data <= 21'h000084; 
        10'b1001001101: data <= 21'h1ffcd4; 
        10'b1001001110: data <= 21'h00011f; 
        10'b1001001111: data <= 21'h1ff37a; 
        10'b1001010000: data <= 21'h1fed67; 
        10'b1001010001: data <= 21'h1ffe25; 
        10'b1001010010: data <= 21'h0009cc; 
        10'b1001010011: data <= 21'h0014ee; 
        10'b1001010100: data <= 21'h000461; 
        10'b1001010101: data <= 21'h0008f8; 
        10'b1001010110: data <= 21'h1ffe5a; 
        10'b1001010111: data <= 21'h1ff22e; 
        10'b1001011000: data <= 21'h1ff844; 
        10'b1001011001: data <= 21'h0004c4; 
        10'b1001011010: data <= 21'h1fff93; 
        10'b1001011011: data <= 21'h1ffdd0; 
        10'b1001011100: data <= 21'h1fefc3; 
        10'b1001011101: data <= 21'h1ff930; 
        10'b1001011110: data <= 21'h1ffb7a; 
        10'b1001011111: data <= 21'h1fff59; 
        10'b1001100000: data <= 21'h1fff9f; 
        10'b1001100001: data <= 21'h0003e4; 
        10'b1001100010: data <= 21'h00035e; 
        10'b1001100011: data <= 21'h1ffb1e; 
        10'b1001100100: data <= 21'h1ffa1d; 
        10'b1001100101: data <= 21'h1fffa2; 
        10'b1001100110: data <= 21'h1ffec8; 
        10'b1001100111: data <= 21'h1ffc3b; 
        10'b1001101000: data <= 21'h1ffe1c; 
        10'b1001101001: data <= 21'h1ff8e3; 
        10'b1001101010: data <= 21'h1ffb75; 
        10'b1001101011: data <= 21'h1ff80a; 
        10'b1001101100: data <= 21'h1ff129; 
        10'b1001101101: data <= 21'h1fe9dd; 
        10'b1001101110: data <= 21'h0002a0; 
        10'b1001101111: data <= 21'h0005f5; 
        10'b1001110000: data <= 21'h1ffea3; 
        10'b1001110001: data <= 21'h1ff8ec; 
        10'b1001110010: data <= 21'h00047c; 
        10'b1001110011: data <= 21'h000199; 
        10'b1001110100: data <= 21'h001a6f; 
        10'b1001110101: data <= 21'h001bb8; 
        10'b1001110110: data <= 21'h001398; 
        10'b1001110111: data <= 21'h000f50; 
        10'b1001111000: data <= 21'h1ffeaf; 
        10'b1001111001: data <= 21'h1ffe8e; 
        10'b1001111010: data <= 21'h00069f; 
        10'b1001111011: data <= 21'h1ff7c4; 
        10'b1001111100: data <= 21'h1ff719; 
        10'b1001111101: data <= 21'h0003cb; 
        10'b1001111110: data <= 21'h1ffe68; 
        10'b1001111111: data <= 21'h1ffa53; 
        10'b1010000000: data <= 21'h1ffe94; 
        10'b1010000001: data <= 21'h1ffe8a; 
        10'b1010000010: data <= 21'h1ffe5b; 
        10'b1010000011: data <= 21'h1ffa83; 
        10'b1010000100: data <= 21'h1ffa71; 
        10'b1010000101: data <= 21'h1fff4d; 
        10'b1010000110: data <= 21'h1ffd7c; 
        10'b1010000111: data <= 21'h1ff8ea; 
        10'b1010001000: data <= 21'h1ff079; 
        10'b1010001001: data <= 21'h1fdafa; 
        10'b1010001010: data <= 21'h1fe2f9; 
        10'b1010001011: data <= 21'h1ff161; 
        10'b1010001100: data <= 21'h00050d; 
        10'b1010001101: data <= 21'h0004fd; 
        10'b1010001110: data <= 21'h000abc; 
        10'b1010001111: data <= 21'h000e04; 
        10'b1010010000: data <= 21'h001f4d; 
        10'b1010010001: data <= 21'h002d01; 
        10'b1010010010: data <= 21'h00264e; 
        10'b1010010011: data <= 21'h001e89; 
        10'b1010010100: data <= 21'h0018ba; 
        10'b1010010101: data <= 21'h0011b6; 
        10'b1010010110: data <= 21'h000e10; 
        10'b1010010111: data <= 21'h0011fb; 
        10'b1010011000: data <= 21'h000d44; 
        10'b1010011001: data <= 21'h00032f; 
        10'b1010011010: data <= 21'h1ffe53; 
        10'b1010011011: data <= 21'h1ffbd0; 
        10'b1010011100: data <= 21'h1ff7d2; 
        10'b1010011101: data <= 21'h1fff3b; 
        10'b1010011110: data <= 21'h1ff8c1; 
        10'b1010011111: data <= 21'h1ffe90; 
        10'b1010100000: data <= 21'h1fff1d; 
        10'b1010100001: data <= 21'h1ffe92; 
        10'b1010100010: data <= 21'h000161; 
        10'b1010100011: data <= 21'h1ff9a3; 
        10'b1010100100: data <= 21'h1ff991; 
        10'b1010100101: data <= 21'h1fe782; 
        10'b1010100110: data <= 21'h1fde02; 
        10'b1010100111: data <= 21'h1fe376; 
        10'b1010101000: data <= 21'h1ffe3e; 
        10'b1010101001: data <= 21'h0006ab; 
        10'b1010101010: data <= 21'h1ffd78; 
        10'b1010101011: data <= 21'h000c1f; 
        10'b1010101100: data <= 21'h0008ef; 
        10'b1010101101: data <= 21'h0005e4; 
        10'b1010101110: data <= 21'h000ed7; 
        10'b1010101111: data <= 21'h00203f; 
        10'b1010110000: data <= 21'h00223c; 
        10'b1010110001: data <= 21'h0016fe; 
        10'b1010110010: data <= 21'h002032; 
        10'b1010110011: data <= 21'h001e38; 
        10'b1010110100: data <= 21'h0009f6; 
        10'b1010110101: data <= 21'h000093; 
        10'b1010110110: data <= 21'h1ff929; 
        10'b1010110111: data <= 21'h0000b1; 
        10'b1010111000: data <= 21'h1ffd32; 
        10'b1010111001: data <= 21'h1ffb4d; 
        10'b1010111010: data <= 21'h00011b; 
        10'b1010111011: data <= 21'h1ffe21; 
        10'b1010111100: data <= 21'h00017e; 
        10'b1010111101: data <= 21'h1ffeeb; 
        10'b1010111110: data <= 21'h0000b7; 
        10'b1010111111: data <= 21'h1ff993; 
        10'b1011000000: data <= 21'h1ffb25; 
        10'b1011000001: data <= 21'h1ff6e8; 
        10'b1011000010: data <= 21'h1ff32d; 
        10'b1011000011: data <= 21'h1ff00e; 
        10'b1011000100: data <= 21'h1fee37; 
        10'b1011000101: data <= 21'h1fee2a; 
        10'b1011000110: data <= 21'h1ff954; 
        10'b1011000111: data <= 21'h1ff363; 
        10'b1011001000: data <= 21'h1ff888; 
        10'b1011001001: data <= 21'h1ff86b; 
        10'b1011001010: data <= 21'h1fff3e; 
        10'b1011001011: data <= 21'h000b53; 
        10'b1011001100: data <= 21'h000812; 
        10'b1011001101: data <= 21'h000a3e; 
        10'b1011001110: data <= 21'h000bae; 
        10'b1011001111: data <= 21'h0001d9; 
        10'b1011010000: data <= 21'h1ffd84; 
        10'b1011010001: data <= 21'h1fffae; 
        10'b1011010010: data <= 21'h1ff844; 
        10'b1011010011: data <= 21'h1ff891; 
        10'b1011010100: data <= 21'h1fff5e; 
        10'b1011010101: data <= 21'h1ffdf0; 
        10'b1011010110: data <= 21'h1ffb37; 
        10'b1011010111: data <= 21'h1ffdc8; 
        10'b1011011000: data <= 21'h1ffece; 
        10'b1011011001: data <= 21'h00002b; 
        10'b1011011010: data <= 21'h1ffc71; 
        10'b1011011011: data <= 21'h1ffad0; 
        10'b1011011100: data <= 21'h1ff870; 
        10'b1011011101: data <= 21'h1ff9a8; 
        10'b1011011110: data <= 21'h1ff647; 
        10'b1011011111: data <= 21'h1ffd43; 
        10'b1011100000: data <= 21'h1ff733; 
        10'b1011100001: data <= 21'h1ff87f; 
        10'b1011100010: data <= 21'h1ff6f1; 
        10'b1011100011: data <= 21'h1ffad4; 
        10'b1011100100: data <= 21'h1ffa4c; 
        10'b1011100101: data <= 21'h1ffb24; 
        10'b1011100110: data <= 21'h1ff8d0; 
        10'b1011100111: data <= 21'h1ffacc; 
        10'b1011101000: data <= 21'h1ff9b8; 
        10'b1011101001: data <= 21'h1ff7a9; 
        10'b1011101010: data <= 21'h1ff6b2; 
        10'b1011101011: data <= 21'h1ffa26; 
        10'b1011101100: data <= 21'h1ffbf3; 
        10'b1011101101: data <= 21'h1ffebc; 
        10'b1011101110: data <= 21'h1ffc57; 
        10'b1011101111: data <= 21'h0001a8; 
        10'b1011110000: data <= 21'h000182; 
        10'b1011110001: data <= 21'h1ff902; 
        10'b1011110010: data <= 21'h1ffdc9; 
        10'b1011110011: data <= 21'h1ffd0d; 
        10'b1011110100: data <= 21'h1ffe6b; 
        10'b1011110101: data <= 21'h1ffa9e; 
        10'b1011110110: data <= 21'h1ffca3; 
        10'b1011110111: data <= 21'h1ffddf; 
        10'b1011111000: data <= 21'h1ffe2a; 
        10'b1011111001: data <= 21'h1ff8d2; 
        10'b1011111010: data <= 21'h1fffbe; 
        10'b1011111011: data <= 21'h1ffb2a; 
        10'b1011111100: data <= 21'h00012f; 
        10'b1011111101: data <= 21'h1ffc74; 
        10'b1011111110: data <= 21'h1ff9cd; 
        10'b1011111111: data <= 21'h1fff58; 
        10'b1100000000: data <= 21'h1ffaf5; 
        10'b1100000001: data <= 21'h1ff9e9; 
        10'b1100000010: data <= 21'h1ffc36; 
        10'b1100000011: data <= 21'h1ffe61; 
        10'b1100000100: data <= 21'h1ffdbd; 
        10'b1100000101: data <= 21'h000021; 
        10'b1100000110: data <= 21'h0000fe; 
        10'b1100000111: data <= 21'h000169; 
        10'b1100001000: data <= 21'h1ffecc; 
        10'b1100001001: data <= 21'h1ffdf6; 
        10'b1100001010: data <= 21'h1ffeb6; 
        10'b1100001011: data <= 21'h1ffa77; 
        10'b1100001100: data <= 21'h1ffd71; 
        10'b1100001101: data <= 21'h00010a; 
        10'b1100001110: data <= 21'h1ff95d; 
        10'b1100001111: data <= 21'h1ffd7e; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 16) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 22'h3ff8d1; 
        10'b0000000001: data <= 22'h3ffa44; 
        10'b0000000010: data <= 22'h3ff90c; 
        10'b0000000011: data <= 22'h3ffcb0; 
        10'b0000000100: data <= 22'h3ffbce; 
        10'b0000000101: data <= 22'h00016f; 
        10'b0000000110: data <= 22'h3ff153; 
        10'b0000000111: data <= 22'h3ffcda; 
        10'b0000001000: data <= 22'h3ff620; 
        10'b0000001001: data <= 22'h3ff7a2; 
        10'b0000001010: data <= 22'h3ff434; 
        10'b0000001011: data <= 22'h00013a; 
        10'b0000001100: data <= 22'h3ffb50; 
        10'b0000001101: data <= 22'h3fff35; 
        10'b0000001110: data <= 22'h3ff3c4; 
        10'b0000001111: data <= 22'h3fff57; 
        10'b0000010000: data <= 22'h3ffc39; 
        10'b0000010001: data <= 22'h3ff2d4; 
        10'b0000010010: data <= 22'h000150; 
        10'b0000010011: data <= 22'h3ffa36; 
        10'b0000010100: data <= 22'h3ff914; 
        10'b0000010101: data <= 22'h3ff8a5; 
        10'b0000010110: data <= 22'h3ff9ae; 
        10'b0000010111: data <= 22'h0002b9; 
        10'b0000011000: data <= 22'h000011; 
        10'b0000011001: data <= 22'h3ff793; 
        10'b0000011010: data <= 22'h3ff582; 
        10'b0000011011: data <= 22'h3ff968; 
        10'b0000011100: data <= 22'h3ff90f; 
        10'b0000011101: data <= 22'h3ff162; 
        10'b0000011110: data <= 22'h000276; 
        10'b0000011111: data <= 22'h000004; 
        10'b0000100000: data <= 22'h3ff2ab; 
        10'b0000100001: data <= 22'h3ff310; 
        10'b0000100010: data <= 22'h3ff1dd; 
        10'b0000100011: data <= 22'h3ff318; 
        10'b0000100100: data <= 22'h0001d1; 
        10'b0000100101: data <= 22'h3ffa98; 
        10'b0000100110: data <= 22'h3ffa06; 
        10'b0000100111: data <= 22'h3ff179; 
        10'b0000101000: data <= 22'h000199; 
        10'b0000101001: data <= 22'h3ffdb0; 
        10'b0000101010: data <= 22'h3ff618; 
        10'b0000101011: data <= 22'h3ff87c; 
        10'b0000101100: data <= 22'h3ffdc1; 
        10'b0000101101: data <= 22'h3ffb4a; 
        10'b0000101110: data <= 22'h3ff4bc; 
        10'b0000101111: data <= 22'h3ffbb6; 
        10'b0000110000: data <= 22'h000165; 
        10'b0000110001: data <= 22'h3ff25a; 
        10'b0000110010: data <= 22'h3ffd8d; 
        10'b0000110011: data <= 22'h3ff4dc; 
        10'b0000110100: data <= 22'h3ffef3; 
        10'b0000110101: data <= 22'h000306; 
        10'b0000110110: data <= 22'h3ff618; 
        10'b0000110111: data <= 22'h3ff4c6; 
        10'b0000111000: data <= 22'h3ff3c9; 
        10'b0000111001: data <= 22'h3fffc6; 
        10'b0000111010: data <= 22'h3ffb1c; 
        10'b0000111011: data <= 22'h3ff9ed; 
        10'b0000111100: data <= 22'h3ff458; 
        10'b0000111101: data <= 22'h3ff1aa; 
        10'b0000111110: data <= 22'h3ffb30; 
        10'b0000111111: data <= 22'h3ff141; 
        10'b0001000000: data <= 22'h00029e; 
        10'b0001000001: data <= 22'h3ff134; 
        10'b0001000010: data <= 22'h3ff1e5; 
        10'b0001000011: data <= 22'h3ffd1b; 
        10'b0001000100: data <= 22'h3ffb0d; 
        10'b0001000101: data <= 22'h3ff0dc; 
        10'b0001000110: data <= 22'h3ffcf3; 
        10'b0001000111: data <= 22'h3ffbee; 
        10'b0001001000: data <= 22'h3feff2; 
        10'b0001001001: data <= 22'h3ff68c; 
        10'b0001001010: data <= 22'h3ff69c; 
        10'b0001001011: data <= 22'h3ffdfe; 
        10'b0001001100: data <= 22'h3fff86; 
        10'b0001001101: data <= 22'h3fff3f; 
        10'b0001001110: data <= 22'h3ffc74; 
        10'b0001001111: data <= 22'h3ff97f; 
        10'b0001010000: data <= 22'h000165; 
        10'b0001010001: data <= 22'h3ff610; 
        10'b0001010010: data <= 22'h3ffdbe; 
        10'b0001010011: data <= 22'h0001e1; 
        10'b0001010100: data <= 22'h3ff509; 
        10'b0001010101: data <= 22'h3ff9ab; 
        10'b0001010110: data <= 22'h3ff9cd; 
        10'b0001010111: data <= 22'h3ff345; 
        10'b0001011000: data <= 22'h00028f; 
        10'b0001011001: data <= 22'h3ff3f9; 
        10'b0001011010: data <= 22'h3ff239; 
        10'b0001011011: data <= 22'h3ff7b5; 
        10'b0001011100: data <= 22'h3ff194; 
        10'b0001011101: data <= 22'h3ffafa; 
        10'b0001011110: data <= 22'h3ff52a; 
        10'b0001011111: data <= 22'h3febe4; 
        10'b0001100000: data <= 22'h3fe9a3; 
        10'b0001100001: data <= 22'h3fe4e3; 
        10'b0001100010: data <= 22'h3fe980; 
        10'b0001100011: data <= 22'h3ff2a8; 
        10'b0001100100: data <= 22'h3fe96c; 
        10'b0001100101: data <= 22'h3fee78; 
        10'b0001100110: data <= 22'h3ff3c8; 
        10'b0001100111: data <= 22'h3ff883; 
        10'b0001101000: data <= 22'h3feeec; 
        10'b0001101001: data <= 22'h000110; 
        10'b0001101010: data <= 22'h3ff70e; 
        10'b0001101011: data <= 22'h3fff1b; 
        10'b0001101100: data <= 22'h3ff642; 
        10'b0001101101: data <= 22'h3ffce3; 
        10'b0001101110: data <= 22'h3ffb70; 
        10'b0001101111: data <= 22'h3ff298; 
        10'b0001110000: data <= 22'h3ffa24; 
        10'b0001110001: data <= 22'h3ffe50; 
        10'b0001110010: data <= 22'h3ff795; 
        10'b0001110011: data <= 22'h3ff2a0; 
        10'b0001110100: data <= 22'h3fff44; 
        10'b0001110101: data <= 22'h3ffef9; 
        10'b0001110110: data <= 22'h3ffa2d; 
        10'b0001110111: data <= 22'h3ff3de; 
        10'b0001111000: data <= 22'h3ff3d1; 
        10'b0001111001: data <= 22'h3ff8d7; 
        10'b0001111010: data <= 22'h3ff9ac; 
        10'b0001111011: data <= 22'h3ffc83; 
        10'b0001111100: data <= 22'h001375; 
        10'b0001111101: data <= 22'h000c90; 
        10'b0001111110: data <= 22'h002a61; 
        10'b0001111111: data <= 22'h002028; 
        10'b0010000000: data <= 22'h000e9e; 
        10'b0010000001: data <= 22'h000800; 
        10'b0010000010: data <= 22'h000c00; 
        10'b0010000011: data <= 22'h3ff553; 
        10'b0010000100: data <= 22'h3ff300; 
        10'b0010000101: data <= 22'h3ff93d; 
        10'b0010000110: data <= 22'h3fec64; 
        10'b0010000111: data <= 22'h3ff1f2; 
        10'b0010001000: data <= 22'h3fff8d; 
        10'b0010001001: data <= 22'h0000f0; 
        10'b0010001010: data <= 22'h3ff86b; 
        10'b0010001011: data <= 22'h3ffa2b; 
        10'b0010001100: data <= 22'h3ffa6c; 
        10'b0010001101: data <= 22'h3ffd5d; 
        10'b0010001110: data <= 22'h3ffe57; 
        10'b0010001111: data <= 22'h3fff7f; 
        10'b0010010000: data <= 22'h3ff473; 
        10'b0010010001: data <= 22'h3ff92d; 
        10'b0010010010: data <= 22'h3ff608; 
        10'b0010010011: data <= 22'h3fe517; 
        10'b0010010100: data <= 22'h3ff530; 
        10'b0010010101: data <= 22'h00099c; 
        10'b0010010110: data <= 22'h3fe9c4; 
        10'b0010010111: data <= 22'h001d9c; 
        10'b0010011000: data <= 22'h0037ad; 
        10'b0010011001: data <= 22'h002e52; 
        10'b0010011010: data <= 22'h003033; 
        10'b0010011011: data <= 22'h001700; 
        10'b0010011100: data <= 22'h0012fa; 
        10'b0010011101: data <= 22'h002c9b; 
        10'b0010011110: data <= 22'h00023a; 
        10'b0010011111: data <= 22'h3ffdf8; 
        10'b0010100000: data <= 22'h000fea; 
        10'b0010100001: data <= 22'h00083d; 
        10'b0010100010: data <= 22'h3fe4f9; 
        10'b0010100011: data <= 22'h3fe94f; 
        10'b0010100100: data <= 22'h3ff04c; 
        10'b0010100101: data <= 22'h000bf7; 
        10'b0010100110: data <= 22'h3ffb1e; 
        10'b0010100111: data <= 22'h00020d; 
        10'b0010101000: data <= 22'h3ff505; 
        10'b0010101001: data <= 22'h3ff41d; 
        10'b0010101010: data <= 22'h3ff18d; 
        10'b0010101011: data <= 22'h3ff1e4; 
        10'b0010101100: data <= 22'h3fefcf; 
        10'b0010101101: data <= 22'h3ff02b; 
        10'b0010101110: data <= 22'h3fe692; 
        10'b0010101111: data <= 22'h3fe67a; 
        10'b0010110000: data <= 22'h0001c8; 
        10'b0010110001: data <= 22'h000783; 
        10'b0010110010: data <= 22'h3ffe07; 
        10'b0010110011: data <= 22'h000e54; 
        10'b0010110100: data <= 22'h0016ae; 
        10'b0010110101: data <= 22'h00122d; 
        10'b0010110110: data <= 22'h00199f; 
        10'b0010110111: data <= 22'h002ff4; 
        10'b0010111000: data <= 22'h001736; 
        10'b0010111001: data <= 22'h001b4b; 
        10'b0010111010: data <= 22'h0005c3; 
        10'b0010111011: data <= 22'h001f26; 
        10'b0010111100: data <= 22'h000be3; 
        10'b0010111101: data <= 22'h000e9f; 
        10'b0010111110: data <= 22'h001231; 
        10'b0010111111: data <= 22'h0010f9; 
        10'b0011000000: data <= 22'h000e54; 
        10'b0011000001: data <= 22'h000605; 
        10'b0011000010: data <= 22'h3ffa25; 
        10'b0011000011: data <= 22'h3ffe89; 
        10'b0011000100: data <= 22'h00021d; 
        10'b0011000101: data <= 22'h3ff521; 
        10'b0011000110: data <= 22'h3ff33f; 
        10'b0011000111: data <= 22'h3ff60d; 
        10'b0011001000: data <= 22'h3fef1c; 
        10'b0011001001: data <= 22'h3ff9d9; 
        10'b0011001010: data <= 22'h3feea8; 
        10'b0011001011: data <= 22'h3ffefb; 
        10'b0011001100: data <= 22'h001125; 
        10'b0011001101: data <= 22'h000702; 
        10'b0011001110: data <= 22'h00089e; 
        10'b0011001111: data <= 22'h3ffa9a; 
        10'b0011010000: data <= 22'h3fea14; 
        10'b0011010001: data <= 22'h3fef92; 
        10'b0011010010: data <= 22'h3fe7cc; 
        10'b0011010011: data <= 22'h000e84; 
        10'b0011010100: data <= 22'h001238; 
        10'b0011010101: data <= 22'h3ffee0; 
        10'b0011010110: data <= 22'h000c69; 
        10'b0011010111: data <= 22'h3ff273; 
        10'b0011011000: data <= 22'h001295; 
        10'b0011011001: data <= 22'h001cf5; 
        10'b0011011010: data <= 22'h000536; 
        10'b0011011011: data <= 22'h003c08; 
        10'b0011011100: data <= 22'h0024c7; 
        10'b0011011101: data <= 22'h3ffe98; 
        10'b0011011110: data <= 22'h0000e2; 
        10'b0011011111: data <= 22'h3ffd7a; 
        10'b0011100000: data <= 22'h3ffd72; 
        10'b0011100001: data <= 22'h0000cf; 
        10'b0011100010: data <= 22'h3ffd09; 
        10'b0011100011: data <= 22'h3ff425; 
        10'b0011100100: data <= 22'h3ffcda; 
        10'b0011100101: data <= 22'h3ffa6c; 
        10'b0011100110: data <= 22'h0018e1; 
        10'b0011100111: data <= 22'h000f5e; 
        10'b0011101000: data <= 22'h00058b; 
        10'b0011101001: data <= 22'h002b27; 
        10'b0011101010: data <= 22'h000277; 
        10'b0011101011: data <= 22'h000173; 
        10'b0011101100: data <= 22'h001cd4; 
        10'b0011101101: data <= 22'h002558; 
        10'b0011101110: data <= 22'h3fe285; 
        10'b0011101111: data <= 22'h3fe6f5; 
        10'b0011110000: data <= 22'h00146b; 
        10'b0011110001: data <= 22'h3ff188; 
        10'b0011110010: data <= 22'h0006ca; 
        10'b0011110011: data <= 22'h00138b; 
        10'b0011110100: data <= 22'h000ce6; 
        10'b0011110101: data <= 22'h0027cc; 
        10'b0011110110: data <= 22'h001aae; 
        10'b0011110111: data <= 22'h002d5a; 
        10'b0011111000: data <= 22'h002941; 
        10'b0011111001: data <= 22'h3ffb16; 
        10'b0011111010: data <= 22'h3ffc7f; 
        10'b0011111011: data <= 22'h000413; 
        10'b0011111100: data <= 22'h00003f; 
        10'b0011111101: data <= 22'h0000d1; 
        10'b0011111110: data <= 22'h3ff98a; 
        10'b0011111111: data <= 22'h3ff805; 
        10'b0100000000: data <= 22'h3ffba5; 
        10'b0100000001: data <= 22'h001932; 
        10'b0100000010: data <= 22'h0012b1; 
        10'b0100000011: data <= 22'h002682; 
        10'b0100000100: data <= 22'h0033a9; 
        10'b0100000101: data <= 22'h002b8f; 
        10'b0100000110: data <= 22'h001b99; 
        10'b0100000111: data <= 22'h003081; 
        10'b0100001000: data <= 22'h000d28; 
        10'b0100001001: data <= 22'h000e08; 
        10'b0100001010: data <= 22'h3fc744; 
        10'b0100001011: data <= 22'h3fb117; 
        10'b0100001100: data <= 22'h3fe47c; 
        10'b0100001101: data <= 22'h000434; 
        10'b0100001110: data <= 22'h00088d; 
        10'b0100001111: data <= 22'h000f50; 
        10'b0100010000: data <= 22'h00143b; 
        10'b0100010001: data <= 22'h001173; 
        10'b0100010010: data <= 22'h0029ad; 
        10'b0100010011: data <= 22'h002acf; 
        10'b0100010100: data <= 22'h3ff908; 
        10'b0100010101: data <= 22'h3ffa20; 
        10'b0100010110: data <= 22'h000987; 
        10'b0100010111: data <= 22'h3ff2ec; 
        10'b0100011000: data <= 22'h3ff5a0; 
        10'b0100011001: data <= 22'h00006a; 
        10'b0100011010: data <= 22'h3ff4f4; 
        10'b0100011011: data <= 22'h00011a; 
        10'b0100011100: data <= 22'h0009b5; 
        10'b0100011101: data <= 22'h001ef6; 
        10'b0100011110: data <= 22'h001ec3; 
        10'b0100011111: data <= 22'h003863; 
        10'b0100100000: data <= 22'h0029db; 
        10'b0100100001: data <= 22'h0030e9; 
        10'b0100100010: data <= 22'h004778; 
        10'b0100100011: data <= 22'h002242; 
        10'b0100100100: data <= 22'h0023cf; 
        10'b0100100101: data <= 22'h001d32; 
        10'b0100100110: data <= 22'h3ff684; 
        10'b0100100111: data <= 22'h3fb4e3; 
        10'b0100101000: data <= 22'h3fc271; 
        10'b0100101001: data <= 22'h3fed3c; 
        10'b0100101010: data <= 22'h00156a; 
        10'b0100101011: data <= 22'h001550; 
        10'b0100101100: data <= 22'h0015db; 
        10'b0100101101: data <= 22'h0032d4; 
        10'b0100101110: data <= 22'h00383d; 
        10'b0100101111: data <= 22'h002de3; 
        10'b0100110000: data <= 22'h000096; 
        10'b0100110001: data <= 22'h3ffca8; 
        10'b0100110010: data <= 22'h3ffa09; 
        10'b0100110011: data <= 22'h3ff618; 
        10'b0100110100: data <= 22'h3ff4f5; 
        10'b0100110101: data <= 22'h000280; 
        10'b0100110110: data <= 22'h3fff01; 
        10'b0100110111: data <= 22'h3fee94; 
        10'b0100111000: data <= 22'h000ec2; 
        10'b0100111001: data <= 22'h00222a; 
        10'b0100111010: data <= 22'h004110; 
        10'b0100111011: data <= 22'h005472; 
        10'b0100111100: data <= 22'h004261; 
        10'b0100111101: data <= 22'h0053e0; 
        10'b0100111110: data <= 22'h00396e; 
        10'b0100111111: data <= 22'h001b25; 
        10'b0101000000: data <= 22'h0022fb; 
        10'b0101000001: data <= 22'h00537f; 
        10'b0101000010: data <= 22'h0065b0; 
        10'b0101000011: data <= 22'h3ff37f; 
        10'b0101000100: data <= 22'h3fc37c; 
        10'b0101000101: data <= 22'h3feb2f; 
        10'b0101000110: data <= 22'h3fec2f; 
        10'b0101000111: data <= 22'h000854; 
        10'b0101001000: data <= 22'h002dff; 
        10'b0101001001: data <= 22'h00371b; 
        10'b0101001010: data <= 22'h004932; 
        10'b0101001011: data <= 22'h004516; 
        10'b0101001100: data <= 22'h003013; 
        10'b0101001101: data <= 22'h0007ce; 
        10'b0101001110: data <= 22'h00043b; 
        10'b0101001111: data <= 22'h3ffc0f; 
        10'b0101010000: data <= 22'h3ff666; 
        10'b0101010001: data <= 22'h3ffcc1; 
        10'b0101010010: data <= 22'h3ff7e3; 
        10'b0101010011: data <= 22'h3ffc3a; 
        10'b0101010100: data <= 22'h3ffce7; 
        10'b0101010101: data <= 22'h0028dc; 
        10'b0101010110: data <= 22'h0021de; 
        10'b0101010111: data <= 22'h0033bb; 
        10'b0101011000: data <= 22'h0030d2; 
        10'b0101011001: data <= 22'h003d55; 
        10'b0101011010: data <= 22'h000a72; 
        10'b0101011011: data <= 22'h000ea4; 
        10'b0101011100: data <= 22'h00081d; 
        10'b0101011101: data <= 22'h0064d6; 
        10'b0101011110: data <= 22'h006556; 
        10'b0101011111: data <= 22'h0016b7; 
        10'b0101100000: data <= 22'h0003d9; 
        10'b0101100001: data <= 22'h3ff724; 
        10'b0101100010: data <= 22'h3ff8b4; 
        10'b0101100011: data <= 22'h001962; 
        10'b0101100100: data <= 22'h002b1e; 
        10'b0101100101: data <= 22'h004a1b; 
        10'b0101100110: data <= 22'h00564c; 
        10'b0101100111: data <= 22'h0047fe; 
        10'b0101101000: data <= 22'h002d30; 
        10'b0101101001: data <= 22'h001216; 
        10'b0101101010: data <= 22'h0008f6; 
        10'b0101101011: data <= 22'h3ff345; 
        10'b0101101100: data <= 22'h3ff1f7; 
        10'b0101101101: data <= 22'h3ffaec; 
        10'b0101101110: data <= 22'h0002db; 
        10'b0101101111: data <= 22'h3ff3f6; 
        10'b0101110000: data <= 22'h3ff6e2; 
        10'b0101110001: data <= 22'h3fffc8; 
        10'b0101110010: data <= 22'h3ff974; 
        10'b0101110011: data <= 22'h3ff9d4; 
        10'b0101110100: data <= 22'h00058f; 
        10'b0101110101: data <= 22'h3ff88c; 
        10'b0101110110: data <= 22'h3fe9e5; 
        10'b0101110111: data <= 22'h00086b; 
        10'b0101111000: data <= 22'h00250a; 
        10'b0101111001: data <= 22'h005e76; 
        10'b0101111010: data <= 22'h001c44; 
        10'b0101111011: data <= 22'h004578; 
        10'b0101111100: data <= 22'h001ba6; 
        10'b0101111101: data <= 22'h3fee70; 
        10'b0101111110: data <= 22'h0001a7; 
        10'b0101111111: data <= 22'h00024f; 
        10'b0110000000: data <= 22'h001ec4; 
        10'b0110000001: data <= 22'h001bec; 
        10'b0110000010: data <= 22'h000fd5; 
        10'b0110000011: data <= 22'h001682; 
        10'b0110000100: data <= 22'h000bf9; 
        10'b0110000101: data <= 22'h0002a8; 
        10'b0110000110: data <= 22'h0002bb; 
        10'b0110000111: data <= 22'h3ffdaf; 
        10'b0110001000: data <= 22'h3ff770; 
        10'b0110001001: data <= 22'h3ff1b9; 
        10'b0110001010: data <= 22'h3ffe0e; 
        10'b0110001011: data <= 22'h3ffa0d; 
        10'b0110001100: data <= 22'h3ff366; 
        10'b0110001101: data <= 22'h3fe48d; 
        10'b0110001110: data <= 22'h3fcf03; 
        10'b0110001111: data <= 22'h3fc130; 
        10'b0110010000: data <= 22'h3fb5d8; 
        10'b0110010001: data <= 22'h3fc49a; 
        10'b0110010010: data <= 22'h3ff7b3; 
        10'b0110010011: data <= 22'h0025f9; 
        10'b0110010100: data <= 22'h002489; 
        10'b0110010101: data <= 22'h004d36; 
        10'b0110010110: data <= 22'h003dc0; 
        10'b0110010111: data <= 22'h0029c1; 
        10'b0110011000: data <= 22'h3ffaeb; 
        10'b0110011001: data <= 22'h000532; 
        10'b0110011010: data <= 22'h3ff527; 
        10'b0110011011: data <= 22'h3fe6d3; 
        10'b0110011100: data <= 22'h3fd702; 
        10'b0110011101: data <= 22'h3fdb54; 
        10'b0110011110: data <= 22'h3fe075; 
        10'b0110011111: data <= 22'h3fdab9; 
        10'b0110100000: data <= 22'h3fef1b; 
        10'b0110100001: data <= 22'h3ffd8c; 
        10'b0110100010: data <= 22'h3ff0ea; 
        10'b0110100011: data <= 22'h00006f; 
        10'b0110100100: data <= 22'h000130; 
        10'b0110100101: data <= 22'h3ff6d8; 
        10'b0110100110: data <= 22'h3ff57b; 
        10'b0110100111: data <= 22'h3ffb9b; 
        10'b0110101000: data <= 22'h3ff235; 
        10'b0110101001: data <= 22'h3fe4be; 
        10'b0110101010: data <= 22'h3fc2f6; 
        10'b0110101011: data <= 22'h3fb531; 
        10'b0110101100: data <= 22'h3fbbcd; 
        10'b0110101101: data <= 22'h3fef5d; 
        10'b0110101110: data <= 22'h000291; 
        10'b0110101111: data <= 22'h0001ac; 
        10'b0110110000: data <= 22'h0034be; 
        10'b0110110001: data <= 22'h003e5a; 
        10'b0110110010: data <= 22'h00368d; 
        10'b0110110011: data <= 22'h001f75; 
        10'b0110110100: data <= 22'h3ff03b; 
        10'b0110110101: data <= 22'h3ff241; 
        10'b0110110110: data <= 22'h3ff65f; 
        10'b0110110111: data <= 22'h3fc8c4; 
        10'b0110111000: data <= 22'h3fbb35; 
        10'b0110111001: data <= 22'h3fcb3c; 
        10'b0110111010: data <= 22'h3fde8c; 
        10'b0110111011: data <= 22'h3fe025; 
        10'b0110111100: data <= 22'h3fe7f8; 
        10'b0110111101: data <= 22'h3ffbd7; 
        10'b0110111110: data <= 22'h3fef63; 
        10'b0110111111: data <= 22'h00015a; 
        10'b0111000000: data <= 22'h3ff89f; 
        10'b0111000001: data <= 22'h3ff260; 
        10'b0111000010: data <= 22'h3ff694; 
        10'b0111000011: data <= 22'h3ffb0b; 
        10'b0111000100: data <= 22'h3fe9f1; 
        10'b0111000101: data <= 22'h3fd88e; 
        10'b0111000110: data <= 22'h3fc09a; 
        10'b0111000111: data <= 22'h3fda92; 
        10'b0111001000: data <= 22'h001924; 
        10'b0111001001: data <= 22'h001bec; 
        10'b0111001010: data <= 22'h000b6c; 
        10'b0111001011: data <= 22'h001999; 
        10'b0111001100: data <= 22'h0032fe; 
        10'b0111001101: data <= 22'h002caf; 
        10'b0111001110: data <= 22'h001007; 
        10'b0111001111: data <= 22'h001aaa; 
        10'b0111010000: data <= 22'h00090a; 
        10'b0111010001: data <= 22'h3feb1e; 
        10'b0111010010: data <= 22'h3fd36d; 
        10'b0111010011: data <= 22'h3fc04c; 
        10'b0111010100: data <= 22'h3fc04c; 
        10'b0111010101: data <= 22'h3fbf46; 
        10'b0111010110: data <= 22'h3fcc16; 
        10'b0111010111: data <= 22'h3feec8; 
        10'b0111011000: data <= 22'h3fe94d; 
        10'b0111011001: data <= 22'h3ff83f; 
        10'b0111011010: data <= 22'h3ff7f2; 
        10'b0111011011: data <= 22'h3ff200; 
        10'b0111011100: data <= 22'h00031d; 
        10'b0111011101: data <= 22'h000228; 
        10'b0111011110: data <= 22'h3ff514; 
        10'b0111011111: data <= 22'h3ff2a0; 
        10'b0111100000: data <= 22'h3ff166; 
        10'b0111100001: data <= 22'h3fd72a; 
        10'b0111100010: data <= 22'h3fc805; 
        10'b0111100011: data <= 22'h0009e6; 
        10'b0111100100: data <= 22'h003409; 
        10'b0111100101: data <= 22'h004079; 
        10'b0111100110: data <= 22'h0014a2; 
        10'b0111100111: data <= 22'h0030c9; 
        10'b0111101000: data <= 22'h004f64; 
        10'b0111101001: data <= 22'h003028; 
        10'b0111101010: data <= 22'h000412; 
        10'b0111101011: data <= 22'h3ff31b; 
        10'b0111101100: data <= 22'h0005c5; 
        10'b0111101101: data <= 22'h3fe747; 
        10'b0111101110: data <= 22'h3fbe89; 
        10'b0111101111: data <= 22'h3fe0fe; 
        10'b0111110000: data <= 22'h3fe13a; 
        10'b0111110001: data <= 22'h3fd482; 
        10'b0111110010: data <= 22'h3fdfc9; 
        10'b0111110011: data <= 22'h3febb7; 
        10'b0111110100: data <= 22'h3ff472; 
        10'b0111110101: data <= 22'h3fef7f; 
        10'b0111110110: data <= 22'h3ffd45; 
        10'b0111110111: data <= 22'h3ff774; 
        10'b0111111000: data <= 22'h3ff617; 
        10'b0111111001: data <= 22'h0000a1; 
        10'b0111111010: data <= 22'h3ff1d7; 
        10'b0111111011: data <= 22'h3fedda; 
        10'b0111111100: data <= 22'h3fe71b; 
        10'b0111111101: data <= 22'h3fe67d; 
        10'b0111111110: data <= 22'h3ff039; 
        10'b0111111111: data <= 22'h000f60; 
        10'b1000000000: data <= 22'h002ac9; 
        10'b1000000001: data <= 22'h004d36; 
        10'b1000000010: data <= 22'h0035f5; 
        10'b1000000011: data <= 22'h00499c; 
        10'b1000000100: data <= 22'h002fee; 
        10'b1000000101: data <= 22'h001b9e; 
        10'b1000000110: data <= 22'h3fde88; 
        10'b1000000111: data <= 22'h3ff75c; 
        10'b1000001000: data <= 22'h3fed24; 
        10'b1000001001: data <= 22'h3fcdc2; 
        10'b1000001010: data <= 22'h3ff3e4; 
        10'b1000001011: data <= 22'h3ff689; 
        10'b1000001100: data <= 22'h0003b5; 
        10'b1000001101: data <= 22'h3fe457; 
        10'b1000001110: data <= 22'h3ffbcc; 
        10'b1000001111: data <= 22'h3fe882; 
        10'b1000010000: data <= 22'h3fe00f; 
        10'b1000010001: data <= 22'h3fef96; 
        10'b1000010010: data <= 22'h3ffd5d; 
        10'b1000010011: data <= 22'h000205; 
        10'b1000010100: data <= 22'h3ff64e; 
        10'b1000010101: data <= 22'h3ffb33; 
        10'b1000010110: data <= 22'h3ffc65; 
        10'b1000010111: data <= 22'h3fea5e; 
        10'b1000011000: data <= 22'h3fe466; 
        10'b1000011001: data <= 22'h3ff4e1; 
        10'b1000011010: data <= 22'h00075f; 
        10'b1000011011: data <= 22'h001467; 
        10'b1000011100: data <= 22'h00153c; 
        10'b1000011101: data <= 22'h00344a; 
        10'b1000011110: data <= 22'h001adc; 
        10'b1000011111: data <= 22'h3ffc4b; 
        10'b1000100000: data <= 22'h000cc5; 
        10'b1000100001: data <= 22'h3fdcfd; 
        10'b1000100010: data <= 22'h3fd702; 
        10'b1000100011: data <= 22'h3ff054; 
        10'b1000100100: data <= 22'h3ff323; 
        10'b1000100101: data <= 22'h3fef34; 
        10'b1000100110: data <= 22'h000ce4; 
        10'b1000100111: data <= 22'h0003b5; 
        10'b1000101000: data <= 22'h001096; 
        10'b1000101001: data <= 22'h000166; 
        10'b1000101010: data <= 22'h000ac3; 
        10'b1000101011: data <= 22'h3ff6d4; 
        10'b1000101100: data <= 22'h3fe7a2; 
        10'b1000101101: data <= 22'h3ff16f; 
        10'b1000101110: data <= 22'h3ff39b; 
        10'b1000101111: data <= 22'h00017b; 
        10'b1000110000: data <= 22'h3ff419; 
        10'b1000110001: data <= 22'h3ffd6b; 
        10'b1000110010: data <= 22'h3ff518; 
        10'b1000110011: data <= 22'h3ff01c; 
        10'b1000110100: data <= 22'h3fe01c; 
        10'b1000110101: data <= 22'h3ffa9f; 
        10'b1000110110: data <= 22'h000515; 
        10'b1000110111: data <= 22'h002d3e; 
        10'b1000111000: data <= 22'h000d7d; 
        10'b1000111001: data <= 22'h3ffa29; 
        10'b1000111010: data <= 22'h3fffbd; 
        10'b1000111011: data <= 22'h3fd9bf; 
        10'b1000111100: data <= 22'h00026b; 
        10'b1000111101: data <= 22'h3ffefe; 
        10'b1000111110: data <= 22'h3fdbb1; 
        10'b1000111111: data <= 22'h3ff965; 
        10'b1001000000: data <= 22'h3fd597; 
        10'b1001000001: data <= 22'h3ff294; 
        10'b1001000010: data <= 22'h00077f; 
        10'b1001000011: data <= 22'h0004a4; 
        10'b1001000100: data <= 22'h000d6c; 
        10'b1001000101: data <= 22'h0016ca; 
        10'b1001000110: data <= 22'h0016b9; 
        10'b1001000111: data <= 22'h3ffa63; 
        10'b1001001000: data <= 22'h3ff10c; 
        10'b1001001001: data <= 22'h3fec59; 
        10'b1001001010: data <= 22'h3ffa2e; 
        10'b1001001011: data <= 22'h3ff488; 
        10'b1001001100: data <= 22'h000109; 
        10'b1001001101: data <= 22'h3ff9a7; 
        10'b1001001110: data <= 22'h00023d; 
        10'b1001001111: data <= 22'h3fe6f5; 
        10'b1001010000: data <= 22'h3fdace; 
        10'b1001010001: data <= 22'h3ffc4b; 
        10'b1001010010: data <= 22'h001398; 
        10'b1001010011: data <= 22'h0029dd; 
        10'b1001010100: data <= 22'h0008c2; 
        10'b1001010101: data <= 22'h0011f0; 
        10'b1001010110: data <= 22'h3ffcb4; 
        10'b1001010111: data <= 22'h3fe45c; 
        10'b1001011000: data <= 22'h3ff088; 
        10'b1001011001: data <= 22'h000988; 
        10'b1001011010: data <= 22'h3fff26; 
        10'b1001011011: data <= 22'h3ffba0; 
        10'b1001011100: data <= 22'h3fdf86; 
        10'b1001011101: data <= 22'h3ff260; 
        10'b1001011110: data <= 22'h3ff6f4; 
        10'b1001011111: data <= 22'h3ffeb2; 
        10'b1001100000: data <= 22'h3fff3e; 
        10'b1001100001: data <= 22'h0007c9; 
        10'b1001100010: data <= 22'h0006bc; 
        10'b1001100011: data <= 22'h3ff63c; 
        10'b1001100100: data <= 22'h3ff43a; 
        10'b1001100101: data <= 22'h3fff44; 
        10'b1001100110: data <= 22'h3ffd90; 
        10'b1001100111: data <= 22'h3ff876; 
        10'b1001101000: data <= 22'h3ffc38; 
        10'b1001101001: data <= 22'h3ff1c7; 
        10'b1001101010: data <= 22'h3ff6ea; 
        10'b1001101011: data <= 22'h3ff014; 
        10'b1001101100: data <= 22'h3fe252; 
        10'b1001101101: data <= 22'h3fd3ba; 
        10'b1001101110: data <= 22'h000541; 
        10'b1001101111: data <= 22'h000bea; 
        10'b1001110000: data <= 22'h3ffd46; 
        10'b1001110001: data <= 22'h3ff1d9; 
        10'b1001110010: data <= 22'h0008f7; 
        10'b1001110011: data <= 22'h000331; 
        10'b1001110100: data <= 22'h0034de; 
        10'b1001110101: data <= 22'h003770; 
        10'b1001110110: data <= 22'h002730; 
        10'b1001110111: data <= 22'h001ea1; 
        10'b1001111000: data <= 22'h3ffd5e; 
        10'b1001111001: data <= 22'h3ffd1c; 
        10'b1001111010: data <= 22'h000d3d; 
        10'b1001111011: data <= 22'h3fef87; 
        10'b1001111100: data <= 22'h3fee31; 
        10'b1001111101: data <= 22'h000796; 
        10'b1001111110: data <= 22'h3ffcd0; 
        10'b1001111111: data <= 22'h3ff4a7; 
        10'b1010000000: data <= 22'h3ffd29; 
        10'b1010000001: data <= 22'h3ffd15; 
        10'b1010000010: data <= 22'h3ffcb6; 
        10'b1010000011: data <= 22'h3ff506; 
        10'b1010000100: data <= 22'h3ff4e2; 
        10'b1010000101: data <= 22'h3ffe99; 
        10'b1010000110: data <= 22'h3ffaf8; 
        10'b1010000111: data <= 22'h3ff1d5; 
        10'b1010001000: data <= 22'h3fe0f3; 
        10'b1010001001: data <= 22'h3fb5f5; 
        10'b1010001010: data <= 22'h3fc5f1; 
        10'b1010001011: data <= 22'h3fe2c2; 
        10'b1010001100: data <= 22'h000a1a; 
        10'b1010001101: data <= 22'h0009fa; 
        10'b1010001110: data <= 22'h001578; 
        10'b1010001111: data <= 22'h001c09; 
        10'b1010010000: data <= 22'h003e9a; 
        10'b1010010001: data <= 22'h005a02; 
        10'b1010010010: data <= 22'h004c9b; 
        10'b1010010011: data <= 22'h003d12; 
        10'b1010010100: data <= 22'h003174; 
        10'b1010010101: data <= 22'h00236c; 
        10'b1010010110: data <= 22'h001c20; 
        10'b1010010111: data <= 22'h0023f7; 
        10'b1010011000: data <= 22'h001a88; 
        10'b1010011001: data <= 22'h00065e; 
        10'b1010011010: data <= 22'h3ffca6; 
        10'b1010011011: data <= 22'h3ff7a0; 
        10'b1010011100: data <= 22'h3fefa4; 
        10'b1010011101: data <= 22'h3ffe76; 
        10'b1010011110: data <= 22'h3ff182; 
        10'b1010011111: data <= 22'h3ffd20; 
        10'b1010100000: data <= 22'h3ffe3a; 
        10'b1010100001: data <= 22'h3ffd24; 
        10'b1010100010: data <= 22'h0002c2; 
        10'b1010100011: data <= 22'h3ff346; 
        10'b1010100100: data <= 22'h3ff322; 
        10'b1010100101: data <= 22'h3fcf04; 
        10'b1010100110: data <= 22'h3fbc05; 
        10'b1010100111: data <= 22'h3fc6eb; 
        10'b1010101000: data <= 22'h3ffc7d; 
        10'b1010101001: data <= 22'h000d56; 
        10'b1010101010: data <= 22'h3ffaf1; 
        10'b1010101011: data <= 22'h00183e; 
        10'b1010101100: data <= 22'h0011de; 
        10'b1010101101: data <= 22'h000bc9; 
        10'b1010101110: data <= 22'h001dad; 
        10'b1010101111: data <= 22'h00407d; 
        10'b1010110000: data <= 22'h004478; 
        10'b1010110001: data <= 22'h002dfb; 
        10'b1010110010: data <= 22'h004064; 
        10'b1010110011: data <= 22'h003c70; 
        10'b1010110100: data <= 22'h0013ec; 
        10'b1010110101: data <= 22'h000125; 
        10'b1010110110: data <= 22'h3ff252; 
        10'b1010110111: data <= 22'h000163; 
        10'b1010111000: data <= 22'h3ffa63; 
        10'b1010111001: data <= 22'h3ff69a; 
        10'b1010111010: data <= 22'h000237; 
        10'b1010111011: data <= 22'h3ffc42; 
        10'b1010111100: data <= 22'h0002fb; 
        10'b1010111101: data <= 22'h3ffdd7; 
        10'b1010111110: data <= 22'h00016e; 
        10'b1010111111: data <= 22'h3ff326; 
        10'b1011000000: data <= 22'h3ff649; 
        10'b1011000001: data <= 22'h3fedcf; 
        10'b1011000010: data <= 22'h3fe65a; 
        10'b1011000011: data <= 22'h3fe01c; 
        10'b1011000100: data <= 22'h3fdc6e; 
        10'b1011000101: data <= 22'h3fdc53; 
        10'b1011000110: data <= 22'h3ff2a8; 
        10'b1011000111: data <= 22'h3fe6c6; 
        10'b1011001000: data <= 22'h3ff110; 
        10'b1011001001: data <= 22'h3ff0d5; 
        10'b1011001010: data <= 22'h3ffe7d; 
        10'b1011001011: data <= 22'h0016a6; 
        10'b1011001100: data <= 22'h001024; 
        10'b1011001101: data <= 22'h00147d; 
        10'b1011001110: data <= 22'h00175b; 
        10'b1011001111: data <= 22'h0003b2; 
        10'b1011010000: data <= 22'h3ffb08; 
        10'b1011010001: data <= 22'h3fff5d; 
        10'b1011010010: data <= 22'h3ff088; 
        10'b1011010011: data <= 22'h3ff123; 
        10'b1011010100: data <= 22'h3ffebc; 
        10'b1011010101: data <= 22'h3ffbe1; 
        10'b1011010110: data <= 22'h3ff66e; 
        10'b1011010111: data <= 22'h3ffb8f; 
        10'b1011011000: data <= 22'h3ffd9c; 
        10'b1011011001: data <= 22'h000056; 
        10'b1011011010: data <= 22'h3ff8e3; 
        10'b1011011011: data <= 22'h3ff59f; 
        10'b1011011100: data <= 22'h3ff0e0; 
        10'b1011011101: data <= 22'h3ff350; 
        10'b1011011110: data <= 22'h3fec8e; 
        10'b1011011111: data <= 22'h3ffa85; 
        10'b1011100000: data <= 22'h3fee66; 
        10'b1011100001: data <= 22'h3ff0ff; 
        10'b1011100010: data <= 22'h3fede2; 
        10'b1011100011: data <= 22'h3ff5a8; 
        10'b1011100100: data <= 22'h3ff498; 
        10'b1011100101: data <= 22'h3ff649; 
        10'b1011100110: data <= 22'h3ff1a1; 
        10'b1011100111: data <= 22'h3ff597; 
        10'b1011101000: data <= 22'h3ff36f; 
        10'b1011101001: data <= 22'h3fef51; 
        10'b1011101010: data <= 22'h3fed63; 
        10'b1011101011: data <= 22'h3ff44d; 
        10'b1011101100: data <= 22'h3ff7e5; 
        10'b1011101101: data <= 22'h3ffd78; 
        10'b1011101110: data <= 22'h3ff8af; 
        10'b1011101111: data <= 22'h00034f; 
        10'b1011110000: data <= 22'h000304; 
        10'b1011110001: data <= 22'h3ff204; 
        10'b1011110010: data <= 22'h3ffb92; 
        10'b1011110011: data <= 22'h3ffa1a; 
        10'b1011110100: data <= 22'h3ffcd5; 
        10'b1011110101: data <= 22'h3ff53d; 
        10'b1011110110: data <= 22'h3ff946; 
        10'b1011110111: data <= 22'h3ffbbe; 
        10'b1011111000: data <= 22'h3ffc53; 
        10'b1011111001: data <= 22'h3ff1a3; 
        10'b1011111010: data <= 22'h3fff7c; 
        10'b1011111011: data <= 22'h3ff654; 
        10'b1011111100: data <= 22'h00025e; 
        10'b1011111101: data <= 22'h3ff8e7; 
        10'b1011111110: data <= 22'h3ff39a; 
        10'b1011111111: data <= 22'h3ffeaf; 
        10'b1100000000: data <= 22'h3ff5ea; 
        10'b1100000001: data <= 22'h3ff3d2; 
        10'b1100000010: data <= 22'h3ff86c; 
        10'b1100000011: data <= 22'h3ffcc2; 
        10'b1100000100: data <= 22'h3ffb7a; 
        10'b1100000101: data <= 22'h000042; 
        10'b1100000110: data <= 22'h0001fc; 
        10'b1100000111: data <= 22'h0002d1; 
        10'b1100001000: data <= 22'h3ffd99; 
        10'b1100001001: data <= 22'h3ffbed; 
        10'b1100001010: data <= 22'h3ffd6c; 
        10'b1100001011: data <= 22'h3ff4ef; 
        10'b1100001100: data <= 22'h3ffae1; 
        10'b1100001101: data <= 22'h000214; 
        10'b1100001110: data <= 22'h3ff2ba; 
        10'b1100001111: data <= 22'h3ffafc; 
      endcase 
    end 
  end 
endgenerate 
assign dout = data; 
endmodule
