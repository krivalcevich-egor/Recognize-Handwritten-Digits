`timescale 1ns / 1ps 
 
////////////////////////////////////////////////////////////////////////////////// 
// WEIGHT MEMORY (ROM) 
////////////////////////////////////////////////////////////////////////////////// 
module ROM_weights_7 #( 
    parameter int WGHT_INT = 6, // integer part 
    parameter int WGHT_FRC = 16 // fractional part 
)( 
    input logic clk, // clock 
    input logic [9:0] address,
    output [WGHT_INT + WGHT_FRC-1:0] dout 
); 

(* rom_style = "block" *) reg [WGHT_INT + WGHT_FRC-1:0] data;
generate 
  if (WGHT_FRC == 1) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 7'h00; 
        10'b0000000001: data <= 7'h00; 
        10'b0000000010: data <= 7'h00; 
        10'b0000000011: data <= 7'h00; 
        10'b0000000100: data <= 7'h00; 
        10'b0000000101: data <= 7'h00; 
        10'b0000000110: data <= 7'h00; 
        10'b0000000111: data <= 7'h00; 
        10'b0000001000: data <= 7'h00; 
        10'b0000001001: data <= 7'h00; 
        10'b0000001010: data <= 7'h00; 
        10'b0000001011: data <= 7'h00; 
        10'b0000001100: data <= 7'h00; 
        10'b0000001101: data <= 7'h00; 
        10'b0000001110: data <= 7'h00; 
        10'b0000001111: data <= 7'h00; 
        10'b0000010000: data <= 7'h00; 
        10'b0000010001: data <= 7'h00; 
        10'b0000010010: data <= 7'h00; 
        10'b0000010011: data <= 7'h00; 
        10'b0000010100: data <= 7'h00; 
        10'b0000010101: data <= 7'h00; 
        10'b0000010110: data <= 7'h00; 
        10'b0000010111: data <= 7'h00; 
        10'b0000011000: data <= 7'h00; 
        10'b0000011001: data <= 7'h00; 
        10'b0000011010: data <= 7'h00; 
        10'b0000011011: data <= 7'h00; 
        10'b0000011100: data <= 7'h00; 
        10'b0000011101: data <= 7'h00; 
        10'b0000011110: data <= 7'h00; 
        10'b0000011111: data <= 7'h00; 
        10'b0000100000: data <= 7'h00; 
        10'b0000100001: data <= 7'h00; 
        10'b0000100010: data <= 7'h00; 
        10'b0000100011: data <= 7'h00; 
        10'b0000100100: data <= 7'h00; 
        10'b0000100101: data <= 7'h00; 
        10'b0000100110: data <= 7'h00; 
        10'b0000100111: data <= 7'h00; 
        10'b0000101000: data <= 7'h00; 
        10'b0000101001: data <= 7'h00; 
        10'b0000101010: data <= 7'h00; 
        10'b0000101011: data <= 7'h00; 
        10'b0000101100: data <= 7'h00; 
        10'b0000101101: data <= 7'h00; 
        10'b0000101110: data <= 7'h00; 
        10'b0000101111: data <= 7'h00; 
        10'b0000110000: data <= 7'h00; 
        10'b0000110001: data <= 7'h00; 
        10'b0000110010: data <= 7'h00; 
        10'b0000110011: data <= 7'h00; 
        10'b0000110100: data <= 7'h00; 
        10'b0000110101: data <= 7'h00; 
        10'b0000110110: data <= 7'h00; 
        10'b0000110111: data <= 7'h00; 
        10'b0000111000: data <= 7'h00; 
        10'b0000111001: data <= 7'h00; 
        10'b0000111010: data <= 7'h00; 
        10'b0000111011: data <= 7'h00; 
        10'b0000111100: data <= 7'h00; 
        10'b0000111101: data <= 7'h00; 
        10'b0000111110: data <= 7'h00; 
        10'b0000111111: data <= 7'h00; 
        10'b0001000000: data <= 7'h00; 
        10'b0001000001: data <= 7'h00; 
        10'b0001000010: data <= 7'h00; 
        10'b0001000011: data <= 7'h00; 
        10'b0001000100: data <= 7'h00; 
        10'b0001000101: data <= 7'h00; 
        10'b0001000110: data <= 7'h00; 
        10'b0001000111: data <= 7'h00; 
        10'b0001001000: data <= 7'h00; 
        10'b0001001001: data <= 7'h00; 
        10'b0001001010: data <= 7'h00; 
        10'b0001001011: data <= 7'h00; 
        10'b0001001100: data <= 7'h00; 
        10'b0001001101: data <= 7'h00; 
        10'b0001001110: data <= 7'h00; 
        10'b0001001111: data <= 7'h00; 
        10'b0001010000: data <= 7'h00; 
        10'b0001010001: data <= 7'h00; 
        10'b0001010010: data <= 7'h00; 
        10'b0001010011: data <= 7'h00; 
        10'b0001010100: data <= 7'h00; 
        10'b0001010101: data <= 7'h00; 
        10'b0001010110: data <= 7'h00; 
        10'b0001010111: data <= 7'h00; 
        10'b0001011000: data <= 7'h00; 
        10'b0001011001: data <= 7'h00; 
        10'b0001011010: data <= 7'h00; 
        10'b0001011011: data <= 7'h00; 
        10'b0001011100: data <= 7'h00; 
        10'b0001011101: data <= 7'h00; 
        10'b0001011110: data <= 7'h00; 
        10'b0001011111: data <= 7'h00; 
        10'b0001100000: data <= 7'h00; 
        10'b0001100001: data <= 7'h00; 
        10'b0001100010: data <= 7'h00; 
        10'b0001100011: data <= 7'h00; 
        10'b0001100100: data <= 7'h00; 
        10'b0001100101: data <= 7'h00; 
        10'b0001100110: data <= 7'h00; 
        10'b0001100111: data <= 7'h00; 
        10'b0001101000: data <= 7'h00; 
        10'b0001101001: data <= 7'h00; 
        10'b0001101010: data <= 7'h00; 
        10'b0001101011: data <= 7'h00; 
        10'b0001101100: data <= 7'h00; 
        10'b0001101101: data <= 7'h00; 
        10'b0001101110: data <= 7'h00; 
        10'b0001101111: data <= 7'h00; 
        10'b0001110000: data <= 7'h00; 
        10'b0001110001: data <= 7'h00; 
        10'b0001110010: data <= 7'h00; 
        10'b0001110011: data <= 7'h00; 
        10'b0001110100: data <= 7'h00; 
        10'b0001110101: data <= 7'h00; 
        10'b0001110110: data <= 7'h00; 
        10'b0001110111: data <= 7'h00; 
        10'b0001111000: data <= 7'h00; 
        10'b0001111001: data <= 7'h00; 
        10'b0001111010: data <= 7'h00; 
        10'b0001111011: data <= 7'h00; 
        10'b0001111100: data <= 7'h00; 
        10'b0001111101: data <= 7'h00; 
        10'b0001111110: data <= 7'h00; 
        10'b0001111111: data <= 7'h00; 
        10'b0010000000: data <= 7'h00; 
        10'b0010000001: data <= 7'h00; 
        10'b0010000010: data <= 7'h00; 
        10'b0010000011: data <= 7'h00; 
        10'b0010000100: data <= 7'h00; 
        10'b0010000101: data <= 7'h00; 
        10'b0010000110: data <= 7'h00; 
        10'b0010000111: data <= 7'h00; 
        10'b0010001000: data <= 7'h00; 
        10'b0010001001: data <= 7'h00; 
        10'b0010001010: data <= 7'h00; 
        10'b0010001011: data <= 7'h00; 
        10'b0010001100: data <= 7'h00; 
        10'b0010001101: data <= 7'h00; 
        10'b0010001110: data <= 7'h00; 
        10'b0010001111: data <= 7'h00; 
        10'b0010010000: data <= 7'h00; 
        10'b0010010001: data <= 7'h00; 
        10'b0010010010: data <= 7'h00; 
        10'b0010010011: data <= 7'h00; 
        10'b0010010100: data <= 7'h00; 
        10'b0010010101: data <= 7'h00; 
        10'b0010010110: data <= 7'h00; 
        10'b0010010111: data <= 7'h00; 
        10'b0010011000: data <= 7'h00; 
        10'b0010011001: data <= 7'h7f; 
        10'b0010011010: data <= 7'h7f; 
        10'b0010011011: data <= 7'h7f; 
        10'b0010011100: data <= 7'h7f; 
        10'b0010011101: data <= 7'h7f; 
        10'b0010011110: data <= 7'h7f; 
        10'b0010011111: data <= 7'h00; 
        10'b0010100000: data <= 7'h00; 
        10'b0010100001: data <= 7'h00; 
        10'b0010100010: data <= 7'h00; 
        10'b0010100011: data <= 7'h00; 
        10'b0010100100: data <= 7'h00; 
        10'b0010100101: data <= 7'h00; 
        10'b0010100110: data <= 7'h00; 
        10'b0010100111: data <= 7'h00; 
        10'b0010101000: data <= 7'h00; 
        10'b0010101001: data <= 7'h00; 
        10'b0010101010: data <= 7'h00; 
        10'b0010101011: data <= 7'h00; 
        10'b0010101100: data <= 7'h00; 
        10'b0010101101: data <= 7'h00; 
        10'b0010101110: data <= 7'h00; 
        10'b0010101111: data <= 7'h00; 
        10'b0010110000: data <= 7'h00; 
        10'b0010110001: data <= 7'h00; 
        10'b0010110010: data <= 7'h00; 
        10'b0010110011: data <= 7'h00; 
        10'b0010110100: data <= 7'h00; 
        10'b0010110101: data <= 7'h00; 
        10'b0010110110: data <= 7'h00; 
        10'b0010110111: data <= 7'h00; 
        10'b0010111000: data <= 7'h00; 
        10'b0010111001: data <= 7'h00; 
        10'b0010111010: data <= 7'h00; 
        10'b0010111011: data <= 7'h00; 
        10'b0010111100: data <= 7'h00; 
        10'b0010111101: data <= 7'h00; 
        10'b0010111110: data <= 7'h00; 
        10'b0010111111: data <= 7'h00; 
        10'b0011000000: data <= 7'h00; 
        10'b0011000001: data <= 7'h00; 
        10'b0011000010: data <= 7'h00; 
        10'b0011000011: data <= 7'h00; 
        10'b0011000100: data <= 7'h00; 
        10'b0011000101: data <= 7'h00; 
        10'b0011000110: data <= 7'h00; 
        10'b0011000111: data <= 7'h00; 
        10'b0011001000: data <= 7'h00; 
        10'b0011001001: data <= 7'h00; 
        10'b0011001010: data <= 7'h00; 
        10'b0011001011: data <= 7'h00; 
        10'b0011001100: data <= 7'h01; 
        10'b0011001101: data <= 7'h00; 
        10'b0011001110: data <= 7'h00; 
        10'b0011001111: data <= 7'h00; 
        10'b0011010000: data <= 7'h00; 
        10'b0011010001: data <= 7'h00; 
        10'b0011010010: data <= 7'h00; 
        10'b0011010011: data <= 7'h00; 
        10'b0011010100: data <= 7'h00; 
        10'b0011010101: data <= 7'h00; 
        10'b0011010110: data <= 7'h00; 
        10'b0011010111: data <= 7'h00; 
        10'b0011011000: data <= 7'h00; 
        10'b0011011001: data <= 7'h00; 
        10'b0011011010: data <= 7'h00; 
        10'b0011011011: data <= 7'h00; 
        10'b0011011100: data <= 7'h00; 
        10'b0011011101: data <= 7'h00; 
        10'b0011011110: data <= 7'h00; 
        10'b0011011111: data <= 7'h00; 
        10'b0011100000: data <= 7'h00; 
        10'b0011100001: data <= 7'h00; 
        10'b0011100010: data <= 7'h00; 
        10'b0011100011: data <= 7'h00; 
        10'b0011100100: data <= 7'h00; 
        10'b0011100101: data <= 7'h00; 
        10'b0011100110: data <= 7'h00; 
        10'b0011100111: data <= 7'h01; 
        10'b0011101000: data <= 7'h00; 
        10'b0011101001: data <= 7'h00; 
        10'b0011101010: data <= 7'h00; 
        10'b0011101011: data <= 7'h01; 
        10'b0011101100: data <= 7'h00; 
        10'b0011101101: data <= 7'h00; 
        10'b0011101110: data <= 7'h00; 
        10'b0011101111: data <= 7'h00; 
        10'b0011110000: data <= 7'h00; 
        10'b0011110001: data <= 7'h01; 
        10'b0011110010: data <= 7'h00; 
        10'b0011110011: data <= 7'h00; 
        10'b0011110100: data <= 7'h00; 
        10'b0011110101: data <= 7'h00; 
        10'b0011110110: data <= 7'h00; 
        10'b0011110111: data <= 7'h00; 
        10'b0011111000: data <= 7'h00; 
        10'b0011111001: data <= 7'h00; 
        10'b0011111010: data <= 7'h00; 
        10'b0011111011: data <= 7'h00; 
        10'b0011111100: data <= 7'h00; 
        10'b0011111101: data <= 7'h00; 
        10'b0011111110: data <= 7'h00; 
        10'b0011111111: data <= 7'h00; 
        10'b0100000000: data <= 7'h00; 
        10'b0100000001: data <= 7'h00; 
        10'b0100000010: data <= 7'h00; 
        10'b0100000011: data <= 7'h00; 
        10'b0100000100: data <= 7'h00; 
        10'b0100000101: data <= 7'h00; 
        10'b0100000110: data <= 7'h00; 
        10'b0100000111: data <= 7'h00; 
        10'b0100001000: data <= 7'h00; 
        10'b0100001001: data <= 7'h00; 
        10'b0100001010: data <= 7'h01; 
        10'b0100001011: data <= 7'h01; 
        10'b0100001100: data <= 7'h01; 
        10'b0100001101: data <= 7'h01; 
        10'b0100001110: data <= 7'h00; 
        10'b0100001111: data <= 7'h00; 
        10'b0100010000: data <= 7'h00; 
        10'b0100010001: data <= 7'h00; 
        10'b0100010010: data <= 7'h00; 
        10'b0100010011: data <= 7'h00; 
        10'b0100010100: data <= 7'h00; 
        10'b0100010101: data <= 7'h00; 
        10'b0100010110: data <= 7'h00; 
        10'b0100010111: data <= 7'h00; 
        10'b0100011000: data <= 7'h00; 
        10'b0100011001: data <= 7'h00; 
        10'b0100011010: data <= 7'h00; 
        10'b0100011011: data <= 7'h00; 
        10'b0100011100: data <= 7'h00; 
        10'b0100011101: data <= 7'h00; 
        10'b0100011110: data <= 7'h00; 
        10'b0100011111: data <= 7'h00; 
        10'b0100100000: data <= 7'h00; 
        10'b0100100001: data <= 7'h00; 
        10'b0100100010: data <= 7'h00; 
        10'b0100100011: data <= 7'h00; 
        10'b0100100100: data <= 7'h00; 
        10'b0100100101: data <= 7'h01; 
        10'b0100100110: data <= 7'h01; 
        10'b0100100111: data <= 7'h01; 
        10'b0100101000: data <= 7'h01; 
        10'b0100101001: data <= 7'h01; 
        10'b0100101010: data <= 7'h01; 
        10'b0100101011: data <= 7'h01; 
        10'b0100101100: data <= 7'h01; 
        10'b0100101101: data <= 7'h00; 
        10'b0100101110: data <= 7'h00; 
        10'b0100101111: data <= 7'h00; 
        10'b0100110000: data <= 7'h00; 
        10'b0100110001: data <= 7'h00; 
        10'b0100110010: data <= 7'h00; 
        10'b0100110011: data <= 7'h00; 
        10'b0100110100: data <= 7'h00; 
        10'b0100110101: data <= 7'h00; 
        10'b0100110110: data <= 7'h00; 
        10'b0100110111: data <= 7'h00; 
        10'b0100111000: data <= 7'h00; 
        10'b0100111001: data <= 7'h00; 
        10'b0100111010: data <= 7'h00; 
        10'b0100111011: data <= 7'h00; 
        10'b0100111100: data <= 7'h00; 
        10'b0100111101: data <= 7'h00; 
        10'b0100111110: data <= 7'h00; 
        10'b0100111111: data <= 7'h00; 
        10'b0101000000: data <= 7'h00; 
        10'b0101000001: data <= 7'h00; 
        10'b0101000010: data <= 7'h00; 
        10'b0101000011: data <= 7'h01; 
        10'b0101000100: data <= 7'h01; 
        10'b0101000101: data <= 7'h01; 
        10'b0101000110: data <= 7'h01; 
        10'b0101000111: data <= 7'h00; 
        10'b0101001000: data <= 7'h00; 
        10'b0101001001: data <= 7'h00; 
        10'b0101001010: data <= 7'h00; 
        10'b0101001011: data <= 7'h00; 
        10'b0101001100: data <= 7'h00; 
        10'b0101001101: data <= 7'h00; 
        10'b0101001110: data <= 7'h00; 
        10'b0101001111: data <= 7'h00; 
        10'b0101010000: data <= 7'h00; 
        10'b0101010001: data <= 7'h00; 
        10'b0101010010: data <= 7'h00; 
        10'b0101010011: data <= 7'h00; 
        10'b0101010100: data <= 7'h00; 
        10'b0101010101: data <= 7'h00; 
        10'b0101010110: data <= 7'h00; 
        10'b0101010111: data <= 7'h00; 
        10'b0101011000: data <= 7'h00; 
        10'b0101011001: data <= 7'h00; 
        10'b0101011010: data <= 7'h00; 
        10'b0101011011: data <= 7'h00; 
        10'b0101011100: data <= 7'h7f; 
        10'b0101011101: data <= 7'h7f; 
        10'b0101011110: data <= 7'h7f; 
        10'b0101011111: data <= 7'h00; 
        10'b0101100000: data <= 7'h01; 
        10'b0101100001: data <= 7'h01; 
        10'b0101100010: data <= 7'h00; 
        10'b0101100011: data <= 7'h00; 
        10'b0101100100: data <= 7'h00; 
        10'b0101100101: data <= 7'h00; 
        10'b0101100110: data <= 7'h00; 
        10'b0101100111: data <= 7'h00; 
        10'b0101101000: data <= 7'h00; 
        10'b0101101001: data <= 7'h00; 
        10'b0101101010: data <= 7'h00; 
        10'b0101101011: data <= 7'h00; 
        10'b0101101100: data <= 7'h00; 
        10'b0101101101: data <= 7'h00; 
        10'b0101101110: data <= 7'h00; 
        10'b0101101111: data <= 7'h00; 
        10'b0101110000: data <= 7'h00; 
        10'b0101110001: data <= 7'h00; 
        10'b0101110010: data <= 7'h00; 
        10'b0101110011: data <= 7'h00; 
        10'b0101110100: data <= 7'h00; 
        10'b0101110101: data <= 7'h00; 
        10'b0101110110: data <= 7'h00; 
        10'b0101110111: data <= 7'h7f; 
        10'b0101111000: data <= 7'h7e; 
        10'b0101111001: data <= 7'h7e; 
        10'b0101111010: data <= 7'h7f; 
        10'b0101111011: data <= 7'h00; 
        10'b0101111100: data <= 7'h00; 
        10'b0101111101: data <= 7'h00; 
        10'b0101111110: data <= 7'h00; 
        10'b0101111111: data <= 7'h00; 
        10'b0110000000: data <= 7'h00; 
        10'b0110000001: data <= 7'h00; 
        10'b0110000010: data <= 7'h00; 
        10'b0110000011: data <= 7'h00; 
        10'b0110000100: data <= 7'h00; 
        10'b0110000101: data <= 7'h00; 
        10'b0110000110: data <= 7'h00; 
        10'b0110000111: data <= 7'h00; 
        10'b0110001000: data <= 7'h00; 
        10'b0110001001: data <= 7'h00; 
        10'b0110001010: data <= 7'h00; 
        10'b0110001011: data <= 7'h00; 
        10'b0110001100: data <= 7'h00; 
        10'b0110001101: data <= 7'h00; 
        10'b0110001110: data <= 7'h00; 
        10'b0110001111: data <= 7'h00; 
        10'b0110010000: data <= 7'h00; 
        10'b0110010001: data <= 7'h00; 
        10'b0110010010: data <= 7'h7f; 
        10'b0110010011: data <= 7'h7f; 
        10'b0110010100: data <= 7'h7f; 
        10'b0110010101: data <= 7'h7f; 
        10'b0110010110: data <= 7'h00; 
        10'b0110010111: data <= 7'h00; 
        10'b0110011000: data <= 7'h00; 
        10'b0110011001: data <= 7'h00; 
        10'b0110011010: data <= 7'h01; 
        10'b0110011011: data <= 7'h01; 
        10'b0110011100: data <= 7'h00; 
        10'b0110011101: data <= 7'h00; 
        10'b0110011110: data <= 7'h00; 
        10'b0110011111: data <= 7'h00; 
        10'b0110100000: data <= 7'h00; 
        10'b0110100001: data <= 7'h00; 
        10'b0110100010: data <= 7'h00; 
        10'b0110100011: data <= 7'h00; 
        10'b0110100100: data <= 7'h00; 
        10'b0110100101: data <= 7'h00; 
        10'b0110100110: data <= 7'h00; 
        10'b0110100111: data <= 7'h00; 
        10'b0110101000: data <= 7'h00; 
        10'b0110101001: data <= 7'h00; 
        10'b0110101010: data <= 7'h00; 
        10'b0110101011: data <= 7'h00; 
        10'b0110101100: data <= 7'h00; 
        10'b0110101101: data <= 7'h7f; 
        10'b0110101110: data <= 7'h7f; 
        10'b0110101111: data <= 7'h7f; 
        10'b0110110000: data <= 7'h7f; 
        10'b0110110001: data <= 7'h7f; 
        10'b0110110010: data <= 7'h00; 
        10'b0110110011: data <= 7'h00; 
        10'b0110110100: data <= 7'h00; 
        10'b0110110101: data <= 7'h01; 
        10'b0110110110: data <= 7'h01; 
        10'b0110110111: data <= 7'h01; 
        10'b0110111000: data <= 7'h01; 
        10'b0110111001: data <= 7'h01; 
        10'b0110111010: data <= 7'h00; 
        10'b0110111011: data <= 7'h00; 
        10'b0110111100: data <= 7'h00; 
        10'b0110111101: data <= 7'h00; 
        10'b0110111110: data <= 7'h00; 
        10'b0110111111: data <= 7'h00; 
        10'b0111000000: data <= 7'h00; 
        10'b0111000001: data <= 7'h00; 
        10'b0111000010: data <= 7'h00; 
        10'b0111000011: data <= 7'h00; 
        10'b0111000100: data <= 7'h00; 
        10'b0111000101: data <= 7'h00; 
        10'b0111000110: data <= 7'h00; 
        10'b0111000111: data <= 7'h00; 
        10'b0111001000: data <= 7'h00; 
        10'b0111001001: data <= 7'h00; 
        10'b0111001010: data <= 7'h7f; 
        10'b0111001011: data <= 7'h7f; 
        10'b0111001100: data <= 7'h7f; 
        10'b0111001101: data <= 7'h00; 
        10'b0111001110: data <= 7'h00; 
        10'b0111001111: data <= 7'h00; 
        10'b0111010000: data <= 7'h00; 
        10'b0111010001: data <= 7'h01; 
        10'b0111010010: data <= 7'h01; 
        10'b0111010011: data <= 7'h01; 
        10'b0111010100: data <= 7'h00; 
        10'b0111010101: data <= 7'h00; 
        10'b0111010110: data <= 7'h00; 
        10'b0111010111: data <= 7'h00; 
        10'b0111011000: data <= 7'h00; 
        10'b0111011001: data <= 7'h00; 
        10'b0111011010: data <= 7'h00; 
        10'b0111011011: data <= 7'h00; 
        10'b0111011100: data <= 7'h00; 
        10'b0111011101: data <= 7'h00; 
        10'b0111011110: data <= 7'h00; 
        10'b0111011111: data <= 7'h00; 
        10'b0111100000: data <= 7'h00; 
        10'b0111100001: data <= 7'h00; 
        10'b0111100010: data <= 7'h00; 
        10'b0111100011: data <= 7'h00; 
        10'b0111100100: data <= 7'h00; 
        10'b0111100101: data <= 7'h00; 
        10'b0111100110: data <= 7'h00; 
        10'b0111100111: data <= 7'h00; 
        10'b0111101000: data <= 7'h00; 
        10'b0111101001: data <= 7'h00; 
        10'b0111101010: data <= 7'h00; 
        10'b0111101011: data <= 7'h00; 
        10'b0111101100: data <= 7'h00; 
        10'b0111101101: data <= 7'h00; 
        10'b0111101110: data <= 7'h00; 
        10'b0111101111: data <= 7'h00; 
        10'b0111110000: data <= 7'h00; 
        10'b0111110001: data <= 7'h00; 
        10'b0111110010: data <= 7'h00; 
        10'b0111110011: data <= 7'h00; 
        10'b0111110100: data <= 7'h00; 
        10'b0111110101: data <= 7'h00; 
        10'b0111110110: data <= 7'h00; 
        10'b0111110111: data <= 7'h00; 
        10'b0111111000: data <= 7'h00; 
        10'b0111111001: data <= 7'h00; 
        10'b0111111010: data <= 7'h00; 
        10'b0111111011: data <= 7'h00; 
        10'b0111111100: data <= 7'h00; 
        10'b0111111101: data <= 7'h00; 
        10'b0111111110: data <= 7'h00; 
        10'b0111111111: data <= 7'h7f; 
        10'b1000000000: data <= 7'h00; 
        10'b1000000001: data <= 7'h00; 
        10'b1000000010: data <= 7'h7f; 
        10'b1000000011: data <= 7'h00; 
        10'b1000000100: data <= 7'h00; 
        10'b1000000101: data <= 7'h00; 
        10'b1000000110: data <= 7'h00; 
        10'b1000000111: data <= 7'h00; 
        10'b1000001000: data <= 7'h00; 
        10'b1000001001: data <= 7'h00; 
        10'b1000001010: data <= 7'h00; 
        10'b1000001011: data <= 7'h00; 
        10'b1000001100: data <= 7'h00; 
        10'b1000001101: data <= 7'h00; 
        10'b1000001110: data <= 7'h00; 
        10'b1000001111: data <= 7'h00; 
        10'b1000010000: data <= 7'h00; 
        10'b1000010001: data <= 7'h00; 
        10'b1000010010: data <= 7'h00; 
        10'b1000010011: data <= 7'h00; 
        10'b1000010100: data <= 7'h00; 
        10'b1000010101: data <= 7'h00; 
        10'b1000010110: data <= 7'h00; 
        10'b1000010111: data <= 7'h00; 
        10'b1000011000: data <= 7'h00; 
        10'b1000011001: data <= 7'h00; 
        10'b1000011010: data <= 7'h7f; 
        10'b1000011011: data <= 7'h7f; 
        10'b1000011100: data <= 7'h7f; 
        10'b1000011101: data <= 7'h7f; 
        10'b1000011110: data <= 7'h00; 
        10'b1000011111: data <= 7'h00; 
        10'b1000100000: data <= 7'h00; 
        10'b1000100001: data <= 7'h00; 
        10'b1000100010: data <= 7'h00; 
        10'b1000100011: data <= 7'h00; 
        10'b1000100100: data <= 7'h00; 
        10'b1000100101: data <= 7'h00; 
        10'b1000100110: data <= 7'h00; 
        10'b1000100111: data <= 7'h00; 
        10'b1000101000: data <= 7'h7f; 
        10'b1000101001: data <= 7'h7f; 
        10'b1000101010: data <= 7'h00; 
        10'b1000101011: data <= 7'h00; 
        10'b1000101100: data <= 7'h00; 
        10'b1000101101: data <= 7'h00; 
        10'b1000101110: data <= 7'h00; 
        10'b1000101111: data <= 7'h00; 
        10'b1000110000: data <= 7'h00; 
        10'b1000110001: data <= 7'h00; 
        10'b1000110010: data <= 7'h00; 
        10'b1000110011: data <= 7'h00; 
        10'b1000110100: data <= 7'h00; 
        10'b1000110101: data <= 7'h00; 
        10'b1000110110: data <= 7'h7f; 
        10'b1000110111: data <= 7'h7f; 
        10'b1000111000: data <= 7'h7f; 
        10'b1000111001: data <= 7'h7f; 
        10'b1000111010: data <= 7'h00; 
        10'b1000111011: data <= 7'h00; 
        10'b1000111100: data <= 7'h00; 
        10'b1000111101: data <= 7'h00; 
        10'b1000111110: data <= 7'h00; 
        10'b1000111111: data <= 7'h00; 
        10'b1001000000: data <= 7'h00; 
        10'b1001000001: data <= 7'h7f; 
        10'b1001000010: data <= 7'h7f; 
        10'b1001000011: data <= 7'h00; 
        10'b1001000100: data <= 7'h7f; 
        10'b1001000101: data <= 7'h00; 
        10'b1001000110: data <= 7'h00; 
        10'b1001000111: data <= 7'h00; 
        10'b1001001000: data <= 7'h00; 
        10'b1001001001: data <= 7'h00; 
        10'b1001001010: data <= 7'h00; 
        10'b1001001011: data <= 7'h00; 
        10'b1001001100: data <= 7'h00; 
        10'b1001001101: data <= 7'h00; 
        10'b1001001110: data <= 7'h00; 
        10'b1001001111: data <= 7'h00; 
        10'b1001010000: data <= 7'h00; 
        10'b1001010001: data <= 7'h00; 
        10'b1001010010: data <= 7'h00; 
        10'b1001010011: data <= 7'h00; 
        10'b1001010100: data <= 7'h00; 
        10'b1001010101: data <= 7'h00; 
        10'b1001010110: data <= 7'h00; 
        10'b1001010111: data <= 7'h00; 
        10'b1001011000: data <= 7'h00; 
        10'b1001011001: data <= 7'h00; 
        10'b1001011010: data <= 7'h00; 
        10'b1001011011: data <= 7'h00; 
        10'b1001011100: data <= 7'h00; 
        10'b1001011101: data <= 7'h7f; 
        10'b1001011110: data <= 7'h7f; 
        10'b1001011111: data <= 7'h7f; 
        10'b1001100000: data <= 7'h7f; 
        10'b1001100001: data <= 7'h00; 
        10'b1001100010: data <= 7'h00; 
        10'b1001100011: data <= 7'h00; 
        10'b1001100100: data <= 7'h00; 
        10'b1001100101: data <= 7'h00; 
        10'b1001100110: data <= 7'h00; 
        10'b1001100111: data <= 7'h00; 
        10'b1001101000: data <= 7'h00; 
        10'b1001101001: data <= 7'h00; 
        10'b1001101010: data <= 7'h00; 
        10'b1001101011: data <= 7'h00; 
        10'b1001101100: data <= 7'h00; 
        10'b1001101101: data <= 7'h00; 
        10'b1001101110: data <= 7'h00; 
        10'b1001101111: data <= 7'h00; 
        10'b1001110000: data <= 7'h00; 
        10'b1001110001: data <= 7'h00; 
        10'b1001110010: data <= 7'h00; 
        10'b1001110011: data <= 7'h00; 
        10'b1001110100: data <= 7'h00; 
        10'b1001110101: data <= 7'h00; 
        10'b1001110110: data <= 7'h00; 
        10'b1001110111: data <= 7'h00; 
        10'b1001111000: data <= 7'h00; 
        10'b1001111001: data <= 7'h00; 
        10'b1001111010: data <= 7'h00; 
        10'b1001111011: data <= 7'h00; 
        10'b1001111100: data <= 7'h00; 
        10'b1001111101: data <= 7'h00; 
        10'b1001111110: data <= 7'h00; 
        10'b1001111111: data <= 7'h00; 
        10'b1010000000: data <= 7'h00; 
        10'b1010000001: data <= 7'h00; 
        10'b1010000010: data <= 7'h00; 
        10'b1010000011: data <= 7'h00; 
        10'b1010000100: data <= 7'h00; 
        10'b1010000101: data <= 7'h00; 
        10'b1010000110: data <= 7'h00; 
        10'b1010000111: data <= 7'h00; 
        10'b1010001000: data <= 7'h00; 
        10'b1010001001: data <= 7'h00; 
        10'b1010001010: data <= 7'h00; 
        10'b1010001011: data <= 7'h00; 
        10'b1010001100: data <= 7'h00; 
        10'b1010001101: data <= 7'h00; 
        10'b1010001110: data <= 7'h00; 
        10'b1010001111: data <= 7'h00; 
        10'b1010010000: data <= 7'h00; 
        10'b1010010001: data <= 7'h00; 
        10'b1010010010: data <= 7'h00; 
        10'b1010010011: data <= 7'h00; 
        10'b1010010100: data <= 7'h00; 
        10'b1010010101: data <= 7'h00; 
        10'b1010010110: data <= 7'h00; 
        10'b1010010111: data <= 7'h00; 
        10'b1010011000: data <= 7'h00; 
        10'b1010011001: data <= 7'h00; 
        10'b1010011010: data <= 7'h00; 
        10'b1010011011: data <= 7'h00; 
        10'b1010011100: data <= 7'h00; 
        10'b1010011101: data <= 7'h00; 
        10'b1010011110: data <= 7'h00; 
        10'b1010011111: data <= 7'h00; 
        10'b1010100000: data <= 7'h00; 
        10'b1010100001: data <= 7'h00; 
        10'b1010100010: data <= 7'h00; 
        10'b1010100011: data <= 7'h00; 
        10'b1010100100: data <= 7'h00; 
        10'b1010100101: data <= 7'h00; 
        10'b1010100110: data <= 7'h00; 
        10'b1010100111: data <= 7'h00; 
        10'b1010101000: data <= 7'h00; 
        10'b1010101001: data <= 7'h00; 
        10'b1010101010: data <= 7'h00; 
        10'b1010101011: data <= 7'h00; 
        10'b1010101100: data <= 7'h00; 
        10'b1010101101: data <= 7'h00; 
        10'b1010101110: data <= 7'h00; 
        10'b1010101111: data <= 7'h00; 
        10'b1010110000: data <= 7'h00; 
        10'b1010110001: data <= 7'h00; 
        10'b1010110010: data <= 7'h00; 
        10'b1010110011: data <= 7'h00; 
        10'b1010110100: data <= 7'h00; 
        10'b1010110101: data <= 7'h00; 
        10'b1010110110: data <= 7'h00; 
        10'b1010110111: data <= 7'h00; 
        10'b1010111000: data <= 7'h00; 
        10'b1010111001: data <= 7'h00; 
        10'b1010111010: data <= 7'h00; 
        10'b1010111011: data <= 7'h00; 
        10'b1010111100: data <= 7'h00; 
        10'b1010111101: data <= 7'h00; 
        10'b1010111110: data <= 7'h00; 
        10'b1010111111: data <= 7'h00; 
        10'b1011000000: data <= 7'h00; 
        10'b1011000001: data <= 7'h00; 
        10'b1011000010: data <= 7'h00; 
        10'b1011000011: data <= 7'h00; 
        10'b1011000100: data <= 7'h00; 
        10'b1011000101: data <= 7'h00; 
        10'b1011000110: data <= 7'h01; 
        10'b1011000111: data <= 7'h01; 
        10'b1011001000: data <= 7'h00; 
        10'b1011001001: data <= 7'h00; 
        10'b1011001010: data <= 7'h00; 
        10'b1011001011: data <= 7'h00; 
        10'b1011001100: data <= 7'h00; 
        10'b1011001101: data <= 7'h00; 
        10'b1011001110: data <= 7'h00; 
        10'b1011001111: data <= 7'h00; 
        10'b1011010000: data <= 7'h00; 
        10'b1011010001: data <= 7'h00; 
        10'b1011010010: data <= 7'h00; 
        10'b1011010011: data <= 7'h00; 
        10'b1011010100: data <= 7'h00; 
        10'b1011010101: data <= 7'h00; 
        10'b1011010110: data <= 7'h00; 
        10'b1011010111: data <= 7'h00; 
        10'b1011011000: data <= 7'h00; 
        10'b1011011001: data <= 7'h00; 
        10'b1011011010: data <= 7'h00; 
        10'b1011011011: data <= 7'h00; 
        10'b1011011100: data <= 7'h00; 
        10'b1011011101: data <= 7'h00; 
        10'b1011011110: data <= 7'h00; 
        10'b1011011111: data <= 7'h00; 
        10'b1011100000: data <= 7'h00; 
        10'b1011100001: data <= 7'h00; 
        10'b1011100010: data <= 7'h00; 
        10'b1011100011: data <= 7'h00; 
        10'b1011100100: data <= 7'h00; 
        10'b1011100101: data <= 7'h00; 
        10'b1011100110: data <= 7'h00; 
        10'b1011100111: data <= 7'h00; 
        10'b1011101000: data <= 7'h00; 
        10'b1011101001: data <= 7'h00; 
        10'b1011101010: data <= 7'h00; 
        10'b1011101011: data <= 7'h00; 
        10'b1011101100: data <= 7'h00; 
        10'b1011101101: data <= 7'h00; 
        10'b1011101110: data <= 7'h00; 
        10'b1011101111: data <= 7'h00; 
        10'b1011110000: data <= 7'h00; 
        10'b1011110001: data <= 7'h00; 
        10'b1011110010: data <= 7'h00; 
        10'b1011110011: data <= 7'h00; 
        10'b1011110100: data <= 7'h00; 
        10'b1011110101: data <= 7'h00; 
        10'b1011110110: data <= 7'h00; 
        10'b1011110111: data <= 7'h00; 
        10'b1011111000: data <= 7'h00; 
        10'b1011111001: data <= 7'h00; 
        10'b1011111010: data <= 7'h00; 
        10'b1011111011: data <= 7'h00; 
        10'b1011111100: data <= 7'h00; 
        10'b1011111101: data <= 7'h00; 
        10'b1011111110: data <= 7'h00; 
        10'b1011111111: data <= 7'h00; 
        10'b1100000000: data <= 7'h00; 
        10'b1100000001: data <= 7'h00; 
        10'b1100000010: data <= 7'h00; 
        10'b1100000011: data <= 7'h00; 
        10'b1100000100: data <= 7'h00; 
        10'b1100000101: data <= 7'h00; 
        10'b1100000110: data <= 7'h00; 
        10'b1100000111: data <= 7'h00; 
        10'b1100001000: data <= 7'h00; 
        10'b1100001001: data <= 7'h00; 
        10'b1100001010: data <= 7'h00; 
        10'b1100001011: data <= 7'h00; 
        10'b1100001100: data <= 7'h00; 
        10'b1100001101: data <= 7'h00; 
        10'b1100001110: data <= 7'h00; 
        10'b1100001111: data <= 7'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 2) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 8'h00; 
        10'b0000000001: data <= 8'h00; 
        10'b0000000010: data <= 8'h00; 
        10'b0000000011: data <= 8'h00; 
        10'b0000000100: data <= 8'h00; 
        10'b0000000101: data <= 8'h00; 
        10'b0000000110: data <= 8'h00; 
        10'b0000000111: data <= 8'h00; 
        10'b0000001000: data <= 8'h00; 
        10'b0000001001: data <= 8'h00; 
        10'b0000001010: data <= 8'h00; 
        10'b0000001011: data <= 8'h00; 
        10'b0000001100: data <= 8'h00; 
        10'b0000001101: data <= 8'h00; 
        10'b0000001110: data <= 8'h00; 
        10'b0000001111: data <= 8'h00; 
        10'b0000010000: data <= 8'h00; 
        10'b0000010001: data <= 8'h00; 
        10'b0000010010: data <= 8'h00; 
        10'b0000010011: data <= 8'h00; 
        10'b0000010100: data <= 8'h00; 
        10'b0000010101: data <= 8'h00; 
        10'b0000010110: data <= 8'h00; 
        10'b0000010111: data <= 8'h00; 
        10'b0000011000: data <= 8'h00; 
        10'b0000011001: data <= 8'h00; 
        10'b0000011010: data <= 8'h00; 
        10'b0000011011: data <= 8'h00; 
        10'b0000011100: data <= 8'h00; 
        10'b0000011101: data <= 8'h00; 
        10'b0000011110: data <= 8'h00; 
        10'b0000011111: data <= 8'h00; 
        10'b0000100000: data <= 8'h00; 
        10'b0000100001: data <= 8'h00; 
        10'b0000100010: data <= 8'h00; 
        10'b0000100011: data <= 8'h00; 
        10'b0000100100: data <= 8'h00; 
        10'b0000100101: data <= 8'h00; 
        10'b0000100110: data <= 8'h00; 
        10'b0000100111: data <= 8'h00; 
        10'b0000101000: data <= 8'h00; 
        10'b0000101001: data <= 8'h00; 
        10'b0000101010: data <= 8'h00; 
        10'b0000101011: data <= 8'h00; 
        10'b0000101100: data <= 8'h00; 
        10'b0000101101: data <= 8'h00; 
        10'b0000101110: data <= 8'h00; 
        10'b0000101111: data <= 8'h00; 
        10'b0000110000: data <= 8'h00; 
        10'b0000110001: data <= 8'h00; 
        10'b0000110010: data <= 8'h00; 
        10'b0000110011: data <= 8'h00; 
        10'b0000110100: data <= 8'h00; 
        10'b0000110101: data <= 8'h00; 
        10'b0000110110: data <= 8'h00; 
        10'b0000110111: data <= 8'h00; 
        10'b0000111000: data <= 8'h00; 
        10'b0000111001: data <= 8'h00; 
        10'b0000111010: data <= 8'h00; 
        10'b0000111011: data <= 8'h00; 
        10'b0000111100: data <= 8'h00; 
        10'b0000111101: data <= 8'h00; 
        10'b0000111110: data <= 8'h00; 
        10'b0000111111: data <= 8'h00; 
        10'b0001000000: data <= 8'h00; 
        10'b0001000001: data <= 8'h00; 
        10'b0001000010: data <= 8'h00; 
        10'b0001000011: data <= 8'h00; 
        10'b0001000100: data <= 8'h00; 
        10'b0001000101: data <= 8'h00; 
        10'b0001000110: data <= 8'h00; 
        10'b0001000111: data <= 8'h00; 
        10'b0001001000: data <= 8'h00; 
        10'b0001001001: data <= 8'h00; 
        10'b0001001010: data <= 8'h00; 
        10'b0001001011: data <= 8'h00; 
        10'b0001001100: data <= 8'h00; 
        10'b0001001101: data <= 8'h00; 
        10'b0001001110: data <= 8'h00; 
        10'b0001001111: data <= 8'h00; 
        10'b0001010000: data <= 8'h00; 
        10'b0001010001: data <= 8'h00; 
        10'b0001010010: data <= 8'h00; 
        10'b0001010011: data <= 8'h00; 
        10'b0001010100: data <= 8'h00; 
        10'b0001010101: data <= 8'h00; 
        10'b0001010110: data <= 8'h00; 
        10'b0001010111: data <= 8'h00; 
        10'b0001011000: data <= 8'h00; 
        10'b0001011001: data <= 8'h00; 
        10'b0001011010: data <= 8'h00; 
        10'b0001011011: data <= 8'h00; 
        10'b0001011100: data <= 8'h00; 
        10'b0001011101: data <= 8'h00; 
        10'b0001011110: data <= 8'h00; 
        10'b0001011111: data <= 8'h00; 
        10'b0001100000: data <= 8'h00; 
        10'b0001100001: data <= 8'h00; 
        10'b0001100010: data <= 8'h00; 
        10'b0001100011: data <= 8'h00; 
        10'b0001100100: data <= 8'h00; 
        10'b0001100101: data <= 8'h00; 
        10'b0001100110: data <= 8'h00; 
        10'b0001100111: data <= 8'h00; 
        10'b0001101000: data <= 8'h00; 
        10'b0001101001: data <= 8'h00; 
        10'b0001101010: data <= 8'h00; 
        10'b0001101011: data <= 8'h00; 
        10'b0001101100: data <= 8'h00; 
        10'b0001101101: data <= 8'h00; 
        10'b0001101110: data <= 8'h00; 
        10'b0001101111: data <= 8'h00; 
        10'b0001110000: data <= 8'h00; 
        10'b0001110001: data <= 8'h00; 
        10'b0001110010: data <= 8'h00; 
        10'b0001110011: data <= 8'h00; 
        10'b0001110100: data <= 8'h00; 
        10'b0001110101: data <= 8'h00; 
        10'b0001110110: data <= 8'h00; 
        10'b0001110111: data <= 8'h00; 
        10'b0001111000: data <= 8'h00; 
        10'b0001111001: data <= 8'h00; 
        10'b0001111010: data <= 8'h00; 
        10'b0001111011: data <= 8'h00; 
        10'b0001111100: data <= 8'h00; 
        10'b0001111101: data <= 8'h00; 
        10'b0001111110: data <= 8'h00; 
        10'b0001111111: data <= 8'hff; 
        10'b0010000000: data <= 8'h00; 
        10'b0010000001: data <= 8'h00; 
        10'b0010000010: data <= 8'h00; 
        10'b0010000011: data <= 8'h00; 
        10'b0010000100: data <= 8'h00; 
        10'b0010000101: data <= 8'h00; 
        10'b0010000110: data <= 8'h00; 
        10'b0010000111: data <= 8'h00; 
        10'b0010001000: data <= 8'h00; 
        10'b0010001001: data <= 8'h00; 
        10'b0010001010: data <= 8'h00; 
        10'b0010001011: data <= 8'h00; 
        10'b0010001100: data <= 8'h00; 
        10'b0010001101: data <= 8'h00; 
        10'b0010001110: data <= 8'h00; 
        10'b0010001111: data <= 8'h00; 
        10'b0010010000: data <= 8'h00; 
        10'b0010010001: data <= 8'h00; 
        10'b0010010010: data <= 8'h00; 
        10'b0010010011: data <= 8'h00; 
        10'b0010010100: data <= 8'h00; 
        10'b0010010101: data <= 8'h00; 
        10'b0010010110: data <= 8'hff; 
        10'b0010010111: data <= 8'hff; 
        10'b0010011000: data <= 8'hff; 
        10'b0010011001: data <= 8'hff; 
        10'b0010011010: data <= 8'hff; 
        10'b0010011011: data <= 8'hff; 
        10'b0010011100: data <= 8'hff; 
        10'b0010011101: data <= 8'hff; 
        10'b0010011110: data <= 8'hff; 
        10'b0010011111: data <= 8'hff; 
        10'b0010100000: data <= 8'hff; 
        10'b0010100001: data <= 8'h00; 
        10'b0010100010: data <= 8'h00; 
        10'b0010100011: data <= 8'h00; 
        10'b0010100100: data <= 8'h00; 
        10'b0010100101: data <= 8'h00; 
        10'b0010100110: data <= 8'h00; 
        10'b0010100111: data <= 8'h00; 
        10'b0010101000: data <= 8'h00; 
        10'b0010101001: data <= 8'h00; 
        10'b0010101010: data <= 8'h00; 
        10'b0010101011: data <= 8'h00; 
        10'b0010101100: data <= 8'h00; 
        10'b0010101101: data <= 8'h00; 
        10'b0010101110: data <= 8'h00; 
        10'b0010101111: data <= 8'h00; 
        10'b0010110000: data <= 8'h01; 
        10'b0010110001: data <= 8'h00; 
        10'b0010110010: data <= 8'h01; 
        10'b0010110011: data <= 8'h00; 
        10'b0010110100: data <= 8'h00; 
        10'b0010110101: data <= 8'hff; 
        10'b0010110110: data <= 8'hff; 
        10'b0010110111: data <= 8'h00; 
        10'b0010111000: data <= 8'h00; 
        10'b0010111001: data <= 8'h00; 
        10'b0010111010: data <= 8'h00; 
        10'b0010111011: data <= 8'h00; 
        10'b0010111100: data <= 8'hff; 
        10'b0010111101: data <= 8'h00; 
        10'b0010111110: data <= 8'hff; 
        10'b0010111111: data <= 8'h00; 
        10'b0011000000: data <= 8'h00; 
        10'b0011000001: data <= 8'h00; 
        10'b0011000010: data <= 8'h00; 
        10'b0011000011: data <= 8'h00; 
        10'b0011000100: data <= 8'h00; 
        10'b0011000101: data <= 8'h00; 
        10'b0011000110: data <= 8'h00; 
        10'b0011000111: data <= 8'h00; 
        10'b0011001000: data <= 8'h00; 
        10'b0011001001: data <= 8'h00; 
        10'b0011001010: data <= 8'h01; 
        10'b0011001011: data <= 8'h01; 
        10'b0011001100: data <= 8'h01; 
        10'b0011001101: data <= 8'h01; 
        10'b0011001110: data <= 8'h01; 
        10'b0011001111: data <= 8'h01; 
        10'b0011010000: data <= 8'h01; 
        10'b0011010001: data <= 8'h00; 
        10'b0011010010: data <= 8'h00; 
        10'b0011010011: data <= 8'h00; 
        10'b0011010100: data <= 8'h01; 
        10'b0011010101: data <= 8'h01; 
        10'b0011010110: data <= 8'h01; 
        10'b0011010111: data <= 8'h00; 
        10'b0011011000: data <= 8'h00; 
        10'b0011011001: data <= 8'h00; 
        10'b0011011010: data <= 8'h00; 
        10'b0011011011: data <= 8'h00; 
        10'b0011011100: data <= 8'h00; 
        10'b0011011101: data <= 8'h00; 
        10'b0011011110: data <= 8'h00; 
        10'b0011011111: data <= 8'h00; 
        10'b0011100000: data <= 8'h00; 
        10'b0011100001: data <= 8'h00; 
        10'b0011100010: data <= 8'h00; 
        10'b0011100011: data <= 8'h00; 
        10'b0011100100: data <= 8'h01; 
        10'b0011100101: data <= 8'h01; 
        10'b0011100110: data <= 8'h01; 
        10'b0011100111: data <= 8'h01; 
        10'b0011101000: data <= 8'h01; 
        10'b0011101001: data <= 8'h01; 
        10'b0011101010: data <= 8'h01; 
        10'b0011101011: data <= 8'h01; 
        10'b0011101100: data <= 8'h01; 
        10'b0011101101: data <= 8'h00; 
        10'b0011101110: data <= 8'h00; 
        10'b0011101111: data <= 8'h00; 
        10'b0011110000: data <= 8'h01; 
        10'b0011110001: data <= 8'h01; 
        10'b0011110010: data <= 8'h01; 
        10'b0011110011: data <= 8'h01; 
        10'b0011110100: data <= 8'h01; 
        10'b0011110101: data <= 8'h00; 
        10'b0011110110: data <= 8'h00; 
        10'b0011110111: data <= 8'h00; 
        10'b0011111000: data <= 8'h00; 
        10'b0011111001: data <= 8'h00; 
        10'b0011111010: data <= 8'h00; 
        10'b0011111011: data <= 8'h00; 
        10'b0011111100: data <= 8'h00; 
        10'b0011111101: data <= 8'h00; 
        10'b0011111110: data <= 8'h00; 
        10'b0011111111: data <= 8'h00; 
        10'b0100000000: data <= 8'h01; 
        10'b0100000001: data <= 8'h01; 
        10'b0100000010: data <= 8'h00; 
        10'b0100000011: data <= 8'h00; 
        10'b0100000100: data <= 8'h00; 
        10'b0100000101: data <= 8'h00; 
        10'b0100000110: data <= 8'h01; 
        10'b0100000111: data <= 8'h01; 
        10'b0100001000: data <= 8'h01; 
        10'b0100001001: data <= 8'h01; 
        10'b0100001010: data <= 8'h01; 
        10'b0100001011: data <= 8'h01; 
        10'b0100001100: data <= 8'h01; 
        10'b0100001101: data <= 8'h01; 
        10'b0100001110: data <= 8'h01; 
        10'b0100001111: data <= 8'h01; 
        10'b0100010000: data <= 8'h01; 
        10'b0100010001: data <= 8'h01; 
        10'b0100010010: data <= 8'h00; 
        10'b0100010011: data <= 8'h00; 
        10'b0100010100: data <= 8'h00; 
        10'b0100010101: data <= 8'h00; 
        10'b0100010110: data <= 8'h00; 
        10'b0100010111: data <= 8'h00; 
        10'b0100011000: data <= 8'h00; 
        10'b0100011001: data <= 8'h00; 
        10'b0100011010: data <= 8'h00; 
        10'b0100011011: data <= 8'h01; 
        10'b0100011100: data <= 8'h01; 
        10'b0100011101: data <= 8'h01; 
        10'b0100011110: data <= 8'h00; 
        10'b0100011111: data <= 8'h00; 
        10'b0100100000: data <= 8'h00; 
        10'b0100100001: data <= 8'h00; 
        10'b0100100010: data <= 8'h00; 
        10'b0100100011: data <= 8'h01; 
        10'b0100100100: data <= 8'h00; 
        10'b0100100101: data <= 8'h01; 
        10'b0100100110: data <= 8'h01; 
        10'b0100100111: data <= 8'h02; 
        10'b0100101000: data <= 8'h02; 
        10'b0100101001: data <= 8'h01; 
        10'b0100101010: data <= 8'h01; 
        10'b0100101011: data <= 8'h01; 
        10'b0100101100: data <= 8'h01; 
        10'b0100101101: data <= 8'h01; 
        10'b0100101110: data <= 8'h00; 
        10'b0100101111: data <= 8'h00; 
        10'b0100110000: data <= 8'h00; 
        10'b0100110001: data <= 8'h00; 
        10'b0100110010: data <= 8'h00; 
        10'b0100110011: data <= 8'h00; 
        10'b0100110100: data <= 8'h00; 
        10'b0100110101: data <= 8'h00; 
        10'b0100110110: data <= 8'h00; 
        10'b0100110111: data <= 8'h01; 
        10'b0100111000: data <= 8'h01; 
        10'b0100111001: data <= 8'h00; 
        10'b0100111010: data <= 8'h00; 
        10'b0100111011: data <= 8'h00; 
        10'b0100111100: data <= 8'h00; 
        10'b0100111101: data <= 8'h00; 
        10'b0100111110: data <= 8'h00; 
        10'b0100111111: data <= 8'h00; 
        10'b0101000000: data <= 8'h00; 
        10'b0101000001: data <= 8'h00; 
        10'b0101000010: data <= 8'h00; 
        10'b0101000011: data <= 8'h01; 
        10'b0101000100: data <= 8'h02; 
        10'b0101000101: data <= 8'h01; 
        10'b0101000110: data <= 8'h01; 
        10'b0101000111: data <= 8'h01; 
        10'b0101001000: data <= 8'h01; 
        10'b0101001001: data <= 8'h01; 
        10'b0101001010: data <= 8'h00; 
        10'b0101001011: data <= 8'h00; 
        10'b0101001100: data <= 8'h00; 
        10'b0101001101: data <= 8'h00; 
        10'b0101001110: data <= 8'h00; 
        10'b0101001111: data <= 8'h00; 
        10'b0101010000: data <= 8'h00; 
        10'b0101010001: data <= 8'h00; 
        10'b0101010010: data <= 8'h00; 
        10'b0101010011: data <= 8'h00; 
        10'b0101010100: data <= 8'h00; 
        10'b0101010101: data <= 8'h00; 
        10'b0101010110: data <= 8'h00; 
        10'b0101010111: data <= 8'h00; 
        10'b0101011000: data <= 8'h00; 
        10'b0101011001: data <= 8'h00; 
        10'b0101011010: data <= 8'h00; 
        10'b0101011011: data <= 8'hff; 
        10'b0101011100: data <= 8'hfe; 
        10'b0101011101: data <= 8'hfd; 
        10'b0101011110: data <= 8'hfe; 
        10'b0101011111: data <= 8'h00; 
        10'b0101100000: data <= 8'h01; 
        10'b0101100001: data <= 8'h01; 
        10'b0101100010: data <= 8'h00; 
        10'b0101100011: data <= 8'h00; 
        10'b0101100100: data <= 8'h00; 
        10'b0101100101: data <= 8'h00; 
        10'b0101100110: data <= 8'h00; 
        10'b0101100111: data <= 8'h00; 
        10'b0101101000: data <= 8'h00; 
        10'b0101101001: data <= 8'h00; 
        10'b0101101010: data <= 8'h00; 
        10'b0101101011: data <= 8'h00; 
        10'b0101101100: data <= 8'h00; 
        10'b0101101101: data <= 8'h00; 
        10'b0101101110: data <= 8'h00; 
        10'b0101101111: data <= 8'h00; 
        10'b0101110000: data <= 8'h00; 
        10'b0101110001: data <= 8'h00; 
        10'b0101110010: data <= 8'h00; 
        10'b0101110011: data <= 8'h00; 
        10'b0101110100: data <= 8'h00; 
        10'b0101110101: data <= 8'h00; 
        10'b0101110110: data <= 8'hff; 
        10'b0101110111: data <= 8'hfe; 
        10'b0101111000: data <= 8'hfd; 
        10'b0101111001: data <= 8'hfd; 
        10'b0101111010: data <= 8'hfe; 
        10'b0101111011: data <= 8'h00; 
        10'b0101111100: data <= 8'h01; 
        10'b0101111101: data <= 8'h00; 
        10'b0101111110: data <= 8'h00; 
        10'b0101111111: data <= 8'h00; 
        10'b0110000000: data <= 8'h00; 
        10'b0110000001: data <= 8'h00; 
        10'b0110000010: data <= 8'h00; 
        10'b0110000011: data <= 8'h00; 
        10'b0110000100: data <= 8'h00; 
        10'b0110000101: data <= 8'h00; 
        10'b0110000110: data <= 8'h00; 
        10'b0110000111: data <= 8'h00; 
        10'b0110001000: data <= 8'h00; 
        10'b0110001001: data <= 8'h00; 
        10'b0110001010: data <= 8'h00; 
        10'b0110001011: data <= 8'h00; 
        10'b0110001100: data <= 8'h00; 
        10'b0110001101: data <= 8'h00; 
        10'b0110001110: data <= 8'h00; 
        10'b0110001111: data <= 8'h00; 
        10'b0110010000: data <= 8'h00; 
        10'b0110010001: data <= 8'hff; 
        10'b0110010010: data <= 8'hff; 
        10'b0110010011: data <= 8'hfe; 
        10'b0110010100: data <= 8'hfd; 
        10'b0110010101: data <= 8'hfe; 
        10'b0110010110: data <= 8'hff; 
        10'b0110010111: data <= 8'h00; 
        10'b0110011000: data <= 8'h00; 
        10'b0110011001: data <= 8'h00; 
        10'b0110011010: data <= 8'h01; 
        10'b0110011011: data <= 8'h01; 
        10'b0110011100: data <= 8'h01; 
        10'b0110011101: data <= 8'h00; 
        10'b0110011110: data <= 8'h00; 
        10'b0110011111: data <= 8'h00; 
        10'b0110100000: data <= 8'h00; 
        10'b0110100001: data <= 8'h00; 
        10'b0110100010: data <= 8'h00; 
        10'b0110100011: data <= 8'h00; 
        10'b0110100100: data <= 8'h00; 
        10'b0110100101: data <= 8'h00; 
        10'b0110100110: data <= 8'h00; 
        10'b0110100111: data <= 8'h00; 
        10'b0110101000: data <= 8'h00; 
        10'b0110101001: data <= 8'h00; 
        10'b0110101010: data <= 8'h00; 
        10'b0110101011: data <= 8'h00; 
        10'b0110101100: data <= 8'hff; 
        10'b0110101101: data <= 8'hff; 
        10'b0110101110: data <= 8'hfe; 
        10'b0110101111: data <= 8'hfe; 
        10'b0110110000: data <= 8'hfe; 
        10'b0110110001: data <= 8'hff; 
        10'b0110110010: data <= 8'hff; 
        10'b0110110011: data <= 8'h00; 
        10'b0110110100: data <= 8'h00; 
        10'b0110110101: data <= 8'h01; 
        10'b0110110110: data <= 8'h02; 
        10'b0110110111: data <= 8'h01; 
        10'b0110111000: data <= 8'h01; 
        10'b0110111001: data <= 8'h01; 
        10'b0110111010: data <= 8'h01; 
        10'b0110111011: data <= 8'h00; 
        10'b0110111100: data <= 8'h00; 
        10'b0110111101: data <= 8'h00; 
        10'b0110111110: data <= 8'h00; 
        10'b0110111111: data <= 8'h00; 
        10'b0111000000: data <= 8'h00; 
        10'b0111000001: data <= 8'h00; 
        10'b0111000010: data <= 8'h00; 
        10'b0111000011: data <= 8'h00; 
        10'b0111000100: data <= 8'h00; 
        10'b0111000101: data <= 8'h00; 
        10'b0111000110: data <= 8'h00; 
        10'b0111000111: data <= 8'h00; 
        10'b0111001000: data <= 8'hff; 
        10'b0111001001: data <= 8'hff; 
        10'b0111001010: data <= 8'hff; 
        10'b0111001011: data <= 8'hfe; 
        10'b0111001100: data <= 8'hff; 
        10'b0111001101: data <= 8'hff; 
        10'b0111001110: data <= 8'hff; 
        10'b0111001111: data <= 8'h00; 
        10'b0111010000: data <= 8'h01; 
        10'b0111010001: data <= 8'h01; 
        10'b0111010010: data <= 8'h01; 
        10'b0111010011: data <= 8'h01; 
        10'b0111010100: data <= 8'h01; 
        10'b0111010101: data <= 8'h01; 
        10'b0111010110: data <= 8'h00; 
        10'b0111010111: data <= 8'h00; 
        10'b0111011000: data <= 8'h00; 
        10'b0111011001: data <= 8'h00; 
        10'b0111011010: data <= 8'h00; 
        10'b0111011011: data <= 8'h00; 
        10'b0111011100: data <= 8'h00; 
        10'b0111011101: data <= 8'h00; 
        10'b0111011110: data <= 8'h00; 
        10'b0111011111: data <= 8'h00; 
        10'b0111100000: data <= 8'h00; 
        10'b0111100001: data <= 8'h00; 
        10'b0111100010: data <= 8'hff; 
        10'b0111100011: data <= 8'hff; 
        10'b0111100100: data <= 8'hff; 
        10'b0111100101: data <= 8'hff; 
        10'b0111100110: data <= 8'hff; 
        10'b0111100111: data <= 8'hff; 
        10'b0111101000: data <= 8'h00; 
        10'b0111101001: data <= 8'h00; 
        10'b0111101010: data <= 8'h00; 
        10'b0111101011: data <= 8'h00; 
        10'b0111101100: data <= 8'h00; 
        10'b0111101101: data <= 8'h00; 
        10'b0111101110: data <= 8'h00; 
        10'b0111101111: data <= 8'h00; 
        10'b0111110000: data <= 8'h00; 
        10'b0111110001: data <= 8'h00; 
        10'b0111110010: data <= 8'h00; 
        10'b0111110011: data <= 8'h00; 
        10'b0111110100: data <= 8'h00; 
        10'b0111110101: data <= 8'h00; 
        10'b0111110110: data <= 8'h00; 
        10'b0111110111: data <= 8'h00; 
        10'b0111111000: data <= 8'h00; 
        10'b0111111001: data <= 8'h00; 
        10'b0111111010: data <= 8'h00; 
        10'b0111111011: data <= 8'h00; 
        10'b0111111100: data <= 8'h00; 
        10'b0111111101: data <= 8'hff; 
        10'b0111111110: data <= 8'hff; 
        10'b0111111111: data <= 8'hff; 
        10'b1000000000: data <= 8'hff; 
        10'b1000000001: data <= 8'hff; 
        10'b1000000010: data <= 8'hff; 
        10'b1000000011: data <= 8'h00; 
        10'b1000000100: data <= 8'h00; 
        10'b1000000101: data <= 8'h00; 
        10'b1000000110: data <= 8'h00; 
        10'b1000000111: data <= 8'h00; 
        10'b1000001000: data <= 8'h00; 
        10'b1000001001: data <= 8'h00; 
        10'b1000001010: data <= 8'hff; 
        10'b1000001011: data <= 8'h00; 
        10'b1000001100: data <= 8'hff; 
        10'b1000001101: data <= 8'hff; 
        10'b1000001110: data <= 8'hff; 
        10'b1000001111: data <= 8'h00; 
        10'b1000010000: data <= 8'h00; 
        10'b1000010001: data <= 8'h00; 
        10'b1000010010: data <= 8'h00; 
        10'b1000010011: data <= 8'h00; 
        10'b1000010100: data <= 8'h00; 
        10'b1000010101: data <= 8'h00; 
        10'b1000010110: data <= 8'h00; 
        10'b1000010111: data <= 8'h00; 
        10'b1000011000: data <= 8'h00; 
        10'b1000011001: data <= 8'hff; 
        10'b1000011010: data <= 8'hff; 
        10'b1000011011: data <= 8'hff; 
        10'b1000011100: data <= 8'hff; 
        10'b1000011101: data <= 8'hff; 
        10'b1000011110: data <= 8'hff; 
        10'b1000011111: data <= 8'hff; 
        10'b1000100000: data <= 8'h00; 
        10'b1000100001: data <= 8'h00; 
        10'b1000100010: data <= 8'h00; 
        10'b1000100011: data <= 8'h00; 
        10'b1000100100: data <= 8'h00; 
        10'b1000100101: data <= 8'hff; 
        10'b1000100110: data <= 8'hff; 
        10'b1000100111: data <= 8'hff; 
        10'b1000101000: data <= 8'hff; 
        10'b1000101001: data <= 8'hff; 
        10'b1000101010: data <= 8'hff; 
        10'b1000101011: data <= 8'hff; 
        10'b1000101100: data <= 8'h00; 
        10'b1000101101: data <= 8'h00; 
        10'b1000101110: data <= 8'h00; 
        10'b1000101111: data <= 8'h00; 
        10'b1000110000: data <= 8'h00; 
        10'b1000110001: data <= 8'h00; 
        10'b1000110010: data <= 8'h00; 
        10'b1000110011: data <= 8'h00; 
        10'b1000110100: data <= 8'h00; 
        10'b1000110101: data <= 8'hff; 
        10'b1000110110: data <= 8'hff; 
        10'b1000110111: data <= 8'hff; 
        10'b1000111000: data <= 8'hff; 
        10'b1000111001: data <= 8'hff; 
        10'b1000111010: data <= 8'hff; 
        10'b1000111011: data <= 8'hff; 
        10'b1000111100: data <= 8'h00; 
        10'b1000111101: data <= 8'h00; 
        10'b1000111110: data <= 8'h00; 
        10'b1000111111: data <= 8'hff; 
        10'b1001000000: data <= 8'hff; 
        10'b1001000001: data <= 8'hff; 
        10'b1001000010: data <= 8'hff; 
        10'b1001000011: data <= 8'hff; 
        10'b1001000100: data <= 8'hff; 
        10'b1001000101: data <= 8'hff; 
        10'b1001000110: data <= 8'hff; 
        10'b1001000111: data <= 8'h00; 
        10'b1001001000: data <= 8'h00; 
        10'b1001001001: data <= 8'h00; 
        10'b1001001010: data <= 8'h00; 
        10'b1001001011: data <= 8'h00; 
        10'b1001001100: data <= 8'h00; 
        10'b1001001101: data <= 8'h00; 
        10'b1001001110: data <= 8'h00; 
        10'b1001001111: data <= 8'h00; 
        10'b1001010000: data <= 8'h00; 
        10'b1001010001: data <= 8'h00; 
        10'b1001010010: data <= 8'hff; 
        10'b1001010011: data <= 8'hff; 
        10'b1001010100: data <= 8'hff; 
        10'b1001010101: data <= 8'h00; 
        10'b1001010110: data <= 8'hff; 
        10'b1001010111: data <= 8'h00; 
        10'b1001011000: data <= 8'h00; 
        10'b1001011001: data <= 8'h00; 
        10'b1001011010: data <= 8'h00; 
        10'b1001011011: data <= 8'h00; 
        10'b1001011100: data <= 8'hff; 
        10'b1001011101: data <= 8'hff; 
        10'b1001011110: data <= 8'hff; 
        10'b1001011111: data <= 8'hff; 
        10'b1001100000: data <= 8'hff; 
        10'b1001100001: data <= 8'hff; 
        10'b1001100010: data <= 8'hff; 
        10'b1001100011: data <= 8'h00; 
        10'b1001100100: data <= 8'h00; 
        10'b1001100101: data <= 8'h00; 
        10'b1001100110: data <= 8'h00; 
        10'b1001100111: data <= 8'h00; 
        10'b1001101000: data <= 8'h00; 
        10'b1001101001: data <= 8'h00; 
        10'b1001101010: data <= 8'h00; 
        10'b1001101011: data <= 8'h00; 
        10'b1001101100: data <= 8'h00; 
        10'b1001101101: data <= 8'h00; 
        10'b1001101110: data <= 8'h00; 
        10'b1001101111: data <= 8'h00; 
        10'b1001110000: data <= 8'h00; 
        10'b1001110001: data <= 8'h00; 
        10'b1001110010: data <= 8'h00; 
        10'b1001110011: data <= 8'hff; 
        10'b1001110100: data <= 8'hff; 
        10'b1001110101: data <= 8'h00; 
        10'b1001110110: data <= 8'h00; 
        10'b1001110111: data <= 8'h00; 
        10'b1001111000: data <= 8'h00; 
        10'b1001111001: data <= 8'h00; 
        10'b1001111010: data <= 8'hff; 
        10'b1001111011: data <= 8'hff; 
        10'b1001111100: data <= 8'hff; 
        10'b1001111101: data <= 8'hff; 
        10'b1001111110: data <= 8'h00; 
        10'b1001111111: data <= 8'h00; 
        10'b1010000000: data <= 8'h00; 
        10'b1010000001: data <= 8'h00; 
        10'b1010000010: data <= 8'h00; 
        10'b1010000011: data <= 8'h00; 
        10'b1010000100: data <= 8'h00; 
        10'b1010000101: data <= 8'h00; 
        10'b1010000110: data <= 8'h00; 
        10'b1010000111: data <= 8'h00; 
        10'b1010001000: data <= 8'h00; 
        10'b1010001001: data <= 8'h00; 
        10'b1010001010: data <= 8'h01; 
        10'b1010001011: data <= 8'h01; 
        10'b1010001100: data <= 8'h00; 
        10'b1010001101: data <= 8'h00; 
        10'b1010001110: data <= 8'h00; 
        10'b1010001111: data <= 8'h00; 
        10'b1010010000: data <= 8'h00; 
        10'b1010010001: data <= 8'h00; 
        10'b1010010010: data <= 8'h00; 
        10'b1010010011: data <= 8'h00; 
        10'b1010010100: data <= 8'h00; 
        10'b1010010101: data <= 8'h00; 
        10'b1010010110: data <= 8'hff; 
        10'b1010010111: data <= 8'hff; 
        10'b1010011000: data <= 8'hff; 
        10'b1010011001: data <= 8'hff; 
        10'b1010011010: data <= 8'hff; 
        10'b1010011011: data <= 8'h00; 
        10'b1010011100: data <= 8'h00; 
        10'b1010011101: data <= 8'h00; 
        10'b1010011110: data <= 8'h00; 
        10'b1010011111: data <= 8'h00; 
        10'b1010100000: data <= 8'h00; 
        10'b1010100001: data <= 8'h00; 
        10'b1010100010: data <= 8'h00; 
        10'b1010100011: data <= 8'h00; 
        10'b1010100100: data <= 8'h00; 
        10'b1010100101: data <= 8'h01; 
        10'b1010100110: data <= 8'h01; 
        10'b1010100111: data <= 8'h01; 
        10'b1010101000: data <= 8'h01; 
        10'b1010101001: data <= 8'h00; 
        10'b1010101010: data <= 8'h01; 
        10'b1010101011: data <= 8'h01; 
        10'b1010101100: data <= 8'h00; 
        10'b1010101101: data <= 8'h01; 
        10'b1010101110: data <= 8'h00; 
        10'b1010101111: data <= 8'h01; 
        10'b1010110000: data <= 8'h00; 
        10'b1010110001: data <= 8'h00; 
        10'b1010110010: data <= 8'h00; 
        10'b1010110011: data <= 8'h00; 
        10'b1010110100: data <= 8'h00; 
        10'b1010110101: data <= 8'h00; 
        10'b1010110110: data <= 8'h00; 
        10'b1010110111: data <= 8'h00; 
        10'b1010111000: data <= 8'h00; 
        10'b1010111001: data <= 8'h00; 
        10'b1010111010: data <= 8'h00; 
        10'b1010111011: data <= 8'h00; 
        10'b1010111100: data <= 8'h00; 
        10'b1010111101: data <= 8'h00; 
        10'b1010111110: data <= 8'h00; 
        10'b1010111111: data <= 8'h00; 
        10'b1011000000: data <= 8'h00; 
        10'b1011000001: data <= 8'h00; 
        10'b1011000010: data <= 8'h00; 
        10'b1011000011: data <= 8'h01; 
        10'b1011000100: data <= 8'h01; 
        10'b1011000101: data <= 8'h01; 
        10'b1011000110: data <= 8'h01; 
        10'b1011000111: data <= 8'h01; 
        10'b1011001000: data <= 8'h01; 
        10'b1011001001: data <= 8'h01; 
        10'b1011001010: data <= 8'h01; 
        10'b1011001011: data <= 8'h01; 
        10'b1011001100: data <= 8'h01; 
        10'b1011001101: data <= 8'h01; 
        10'b1011001110: data <= 8'h01; 
        10'b1011001111: data <= 8'h00; 
        10'b1011010000: data <= 8'h00; 
        10'b1011010001: data <= 8'h00; 
        10'b1011010010: data <= 8'h00; 
        10'b1011010011: data <= 8'h00; 
        10'b1011010100: data <= 8'h00; 
        10'b1011010101: data <= 8'h00; 
        10'b1011010110: data <= 8'h00; 
        10'b1011010111: data <= 8'h00; 
        10'b1011011000: data <= 8'h00; 
        10'b1011011001: data <= 8'h00; 
        10'b1011011010: data <= 8'h00; 
        10'b1011011011: data <= 8'h00; 
        10'b1011011100: data <= 8'h00; 
        10'b1011011101: data <= 8'h00; 
        10'b1011011110: data <= 8'h00; 
        10'b1011011111: data <= 8'h00; 
        10'b1011100000: data <= 8'h00; 
        10'b1011100001: data <= 8'h00; 
        10'b1011100010: data <= 8'h00; 
        10'b1011100011: data <= 8'h00; 
        10'b1011100100: data <= 8'h00; 
        10'b1011100101: data <= 8'h00; 
        10'b1011100110: data <= 8'h01; 
        10'b1011100111: data <= 8'h01; 
        10'b1011101000: data <= 8'h01; 
        10'b1011101001: data <= 8'h01; 
        10'b1011101010: data <= 8'h00; 
        10'b1011101011: data <= 8'h00; 
        10'b1011101100: data <= 8'h00; 
        10'b1011101101: data <= 8'h00; 
        10'b1011101110: data <= 8'h00; 
        10'b1011101111: data <= 8'h00; 
        10'b1011110000: data <= 8'h00; 
        10'b1011110001: data <= 8'h00; 
        10'b1011110010: data <= 8'h00; 
        10'b1011110011: data <= 8'h00; 
        10'b1011110100: data <= 8'h00; 
        10'b1011110101: data <= 8'h00; 
        10'b1011110110: data <= 8'h00; 
        10'b1011110111: data <= 8'h00; 
        10'b1011111000: data <= 8'h00; 
        10'b1011111001: data <= 8'h00; 
        10'b1011111010: data <= 8'h00; 
        10'b1011111011: data <= 8'h00; 
        10'b1011111100: data <= 8'h00; 
        10'b1011111101: data <= 8'h00; 
        10'b1011111110: data <= 8'h00; 
        10'b1011111111: data <= 8'h00; 
        10'b1100000000: data <= 8'h00; 
        10'b1100000001: data <= 8'h00; 
        10'b1100000010: data <= 8'h00; 
        10'b1100000011: data <= 8'h00; 
        10'b1100000100: data <= 8'h00; 
        10'b1100000101: data <= 8'h00; 
        10'b1100000110: data <= 8'h00; 
        10'b1100000111: data <= 8'h00; 
        10'b1100001000: data <= 8'h00; 
        10'b1100001001: data <= 8'h00; 
        10'b1100001010: data <= 8'h00; 
        10'b1100001011: data <= 8'h00; 
        10'b1100001100: data <= 8'h00; 
        10'b1100001101: data <= 8'h00; 
        10'b1100001110: data <= 8'h00; 
        10'b1100001111: data <= 8'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 3) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 9'h000; 
        10'b0000000001: data <= 9'h000; 
        10'b0000000010: data <= 9'h000; 
        10'b0000000011: data <= 9'h000; 
        10'b0000000100: data <= 9'h000; 
        10'b0000000101: data <= 9'h000; 
        10'b0000000110: data <= 9'h000; 
        10'b0000000111: data <= 9'h000; 
        10'b0000001000: data <= 9'h000; 
        10'b0000001001: data <= 9'h000; 
        10'b0000001010: data <= 9'h000; 
        10'b0000001011: data <= 9'h000; 
        10'b0000001100: data <= 9'h000; 
        10'b0000001101: data <= 9'h000; 
        10'b0000001110: data <= 9'h000; 
        10'b0000001111: data <= 9'h000; 
        10'b0000010000: data <= 9'h000; 
        10'b0000010001: data <= 9'h000; 
        10'b0000010010: data <= 9'h000; 
        10'b0000010011: data <= 9'h000; 
        10'b0000010100: data <= 9'h000; 
        10'b0000010101: data <= 9'h000; 
        10'b0000010110: data <= 9'h000; 
        10'b0000010111: data <= 9'h000; 
        10'b0000011000: data <= 9'h000; 
        10'b0000011001: data <= 9'h000; 
        10'b0000011010: data <= 9'h000; 
        10'b0000011011: data <= 9'h000; 
        10'b0000011100: data <= 9'h000; 
        10'b0000011101: data <= 9'h000; 
        10'b0000011110: data <= 9'h000; 
        10'b0000011111: data <= 9'h000; 
        10'b0000100000: data <= 9'h000; 
        10'b0000100001: data <= 9'h000; 
        10'b0000100010: data <= 9'h000; 
        10'b0000100011: data <= 9'h000; 
        10'b0000100100: data <= 9'h000; 
        10'b0000100101: data <= 9'h000; 
        10'b0000100110: data <= 9'h000; 
        10'b0000100111: data <= 9'h000; 
        10'b0000101000: data <= 9'h000; 
        10'b0000101001: data <= 9'h000; 
        10'b0000101010: data <= 9'h000; 
        10'b0000101011: data <= 9'h000; 
        10'b0000101100: data <= 9'h000; 
        10'b0000101101: data <= 9'h000; 
        10'b0000101110: data <= 9'h000; 
        10'b0000101111: data <= 9'h000; 
        10'b0000110000: data <= 9'h000; 
        10'b0000110001: data <= 9'h000; 
        10'b0000110010: data <= 9'h000; 
        10'b0000110011: data <= 9'h000; 
        10'b0000110100: data <= 9'h000; 
        10'b0000110101: data <= 9'h000; 
        10'b0000110110: data <= 9'h000; 
        10'b0000110111: data <= 9'h000; 
        10'b0000111000: data <= 9'h000; 
        10'b0000111001: data <= 9'h000; 
        10'b0000111010: data <= 9'h000; 
        10'b0000111011: data <= 9'h000; 
        10'b0000111100: data <= 9'h000; 
        10'b0000111101: data <= 9'h000; 
        10'b0000111110: data <= 9'h000; 
        10'b0000111111: data <= 9'h000; 
        10'b0001000000: data <= 9'h000; 
        10'b0001000001: data <= 9'h000; 
        10'b0001000010: data <= 9'h000; 
        10'b0001000011: data <= 9'h000; 
        10'b0001000100: data <= 9'h000; 
        10'b0001000101: data <= 9'h000; 
        10'b0001000110: data <= 9'h000; 
        10'b0001000111: data <= 9'h000; 
        10'b0001001000: data <= 9'h000; 
        10'b0001001001: data <= 9'h000; 
        10'b0001001010: data <= 9'h000; 
        10'b0001001011: data <= 9'h000; 
        10'b0001001100: data <= 9'h000; 
        10'b0001001101: data <= 9'h000; 
        10'b0001001110: data <= 9'h000; 
        10'b0001001111: data <= 9'h000; 
        10'b0001010000: data <= 9'h000; 
        10'b0001010001: data <= 9'h000; 
        10'b0001010010: data <= 9'h000; 
        10'b0001010011: data <= 9'h000; 
        10'b0001010100: data <= 9'h000; 
        10'b0001010101: data <= 9'h000; 
        10'b0001010110: data <= 9'h000; 
        10'b0001010111: data <= 9'h000; 
        10'b0001011000: data <= 9'h000; 
        10'b0001011001: data <= 9'h000; 
        10'b0001011010: data <= 9'h000; 
        10'b0001011011: data <= 9'h000; 
        10'b0001011100: data <= 9'h000; 
        10'b0001011101: data <= 9'h000; 
        10'b0001011110: data <= 9'h000; 
        10'b0001011111: data <= 9'h000; 
        10'b0001100000: data <= 9'h000; 
        10'b0001100001: data <= 9'h000; 
        10'b0001100010: data <= 9'h000; 
        10'b0001100011: data <= 9'h000; 
        10'b0001100100: data <= 9'h000; 
        10'b0001100101: data <= 9'h000; 
        10'b0001100110: data <= 9'h000; 
        10'b0001100111: data <= 9'h000; 
        10'b0001101000: data <= 9'h000; 
        10'b0001101001: data <= 9'h000; 
        10'b0001101010: data <= 9'h000; 
        10'b0001101011: data <= 9'h000; 
        10'b0001101100: data <= 9'h000; 
        10'b0001101101: data <= 9'h000; 
        10'b0001101110: data <= 9'h000; 
        10'b0001101111: data <= 9'h000; 
        10'b0001110000: data <= 9'h000; 
        10'b0001110001: data <= 9'h000; 
        10'b0001110010: data <= 9'h000; 
        10'b0001110011: data <= 9'h000; 
        10'b0001110100: data <= 9'h000; 
        10'b0001110101: data <= 9'h000; 
        10'b0001110110: data <= 9'h000; 
        10'b0001110111: data <= 9'h000; 
        10'b0001111000: data <= 9'h000; 
        10'b0001111001: data <= 9'h000; 
        10'b0001111010: data <= 9'h000; 
        10'b0001111011: data <= 9'h1ff; 
        10'b0001111100: data <= 9'h1ff; 
        10'b0001111101: data <= 9'h1ff; 
        10'b0001111110: data <= 9'h1ff; 
        10'b0001111111: data <= 9'h1ff; 
        10'b0010000000: data <= 9'h1ff; 
        10'b0010000001: data <= 9'h1ff; 
        10'b0010000010: data <= 9'h1ff; 
        10'b0010000011: data <= 9'h000; 
        10'b0010000100: data <= 9'h000; 
        10'b0010000101: data <= 9'h000; 
        10'b0010000110: data <= 9'h000; 
        10'b0010000111: data <= 9'h000; 
        10'b0010001000: data <= 9'h000; 
        10'b0010001001: data <= 9'h000; 
        10'b0010001010: data <= 9'h000; 
        10'b0010001011: data <= 9'h000; 
        10'b0010001100: data <= 9'h000; 
        10'b0010001101: data <= 9'h000; 
        10'b0010001110: data <= 9'h000; 
        10'b0010001111: data <= 9'h000; 
        10'b0010010000: data <= 9'h000; 
        10'b0010010001: data <= 9'h000; 
        10'b0010010010: data <= 9'h000; 
        10'b0010010011: data <= 9'h000; 
        10'b0010010100: data <= 9'h000; 
        10'b0010010101: data <= 9'h1ff; 
        10'b0010010110: data <= 9'h1ff; 
        10'b0010010111: data <= 9'h1fe; 
        10'b0010011000: data <= 9'h1fe; 
        10'b0010011001: data <= 9'h1fe; 
        10'b0010011010: data <= 9'h1fd; 
        10'b0010011011: data <= 9'h1fd; 
        10'b0010011100: data <= 9'h1fd; 
        10'b0010011101: data <= 9'h1fd; 
        10'b0010011110: data <= 9'h1fe; 
        10'b0010011111: data <= 9'h1fe; 
        10'b0010100000: data <= 9'h1ff; 
        10'b0010100001: data <= 9'h000; 
        10'b0010100010: data <= 9'h1ff; 
        10'b0010100011: data <= 9'h000; 
        10'b0010100100: data <= 9'h000; 
        10'b0010100101: data <= 9'h000; 
        10'b0010100110: data <= 9'h000; 
        10'b0010100111: data <= 9'h000; 
        10'b0010101000: data <= 9'h000; 
        10'b0010101001: data <= 9'h000; 
        10'b0010101010: data <= 9'h000; 
        10'b0010101011: data <= 9'h000; 
        10'b0010101100: data <= 9'h000; 
        10'b0010101101: data <= 9'h000; 
        10'b0010101110: data <= 9'h001; 
        10'b0010101111: data <= 9'h001; 
        10'b0010110000: data <= 9'h001; 
        10'b0010110001: data <= 9'h001; 
        10'b0010110010: data <= 9'h001; 
        10'b0010110011: data <= 9'h000; 
        10'b0010110100: data <= 9'h1ff; 
        10'b0010110101: data <= 9'h1fe; 
        10'b0010110110: data <= 9'h1fe; 
        10'b0010110111: data <= 9'h1ff; 
        10'b0010111000: data <= 9'h1ff; 
        10'b0010111001: data <= 9'h1ff; 
        10'b0010111010: data <= 9'h1ff; 
        10'b0010111011: data <= 9'h1ff; 
        10'b0010111100: data <= 9'h1ff; 
        10'b0010111101: data <= 9'h1ff; 
        10'b0010111110: data <= 9'h1ff; 
        10'b0010111111: data <= 9'h1ff; 
        10'b0011000000: data <= 9'h000; 
        10'b0011000001: data <= 9'h000; 
        10'b0011000010: data <= 9'h000; 
        10'b0011000011: data <= 9'h000; 
        10'b0011000100: data <= 9'h000; 
        10'b0011000101: data <= 9'h000; 
        10'b0011000110: data <= 9'h000; 
        10'b0011000111: data <= 9'h001; 
        10'b0011001000: data <= 9'h001; 
        10'b0011001001: data <= 9'h001; 
        10'b0011001010: data <= 9'h001; 
        10'b0011001011: data <= 9'h002; 
        10'b0011001100: data <= 9'h002; 
        10'b0011001101: data <= 9'h002; 
        10'b0011001110: data <= 9'h001; 
        10'b0011001111: data <= 9'h001; 
        10'b0011010000: data <= 9'h001; 
        10'b0011010001: data <= 9'h000; 
        10'b0011010010: data <= 9'h000; 
        10'b0011010011: data <= 9'h001; 
        10'b0011010100: data <= 9'h002; 
        10'b0011010101: data <= 9'h002; 
        10'b0011010110: data <= 9'h001; 
        10'b0011010111: data <= 9'h001; 
        10'b0011011000: data <= 9'h000; 
        10'b0011011001: data <= 9'h000; 
        10'b0011011010: data <= 9'h000; 
        10'b0011011011: data <= 9'h000; 
        10'b0011011100: data <= 9'h000; 
        10'b0011011101: data <= 9'h000; 
        10'b0011011110: data <= 9'h000; 
        10'b0011011111: data <= 9'h000; 
        10'b0011100000: data <= 9'h000; 
        10'b0011100001: data <= 9'h000; 
        10'b0011100010: data <= 9'h000; 
        10'b0011100011: data <= 9'h001; 
        10'b0011100100: data <= 9'h001; 
        10'b0011100101: data <= 9'h001; 
        10'b0011100110: data <= 9'h001; 
        10'b0011100111: data <= 9'h003; 
        10'b0011101000: data <= 9'h002; 
        10'b0011101001: data <= 9'h001; 
        10'b0011101010: data <= 9'h002; 
        10'b0011101011: data <= 9'h002; 
        10'b0011101100: data <= 9'h002; 
        10'b0011101101: data <= 9'h001; 
        10'b0011101110: data <= 9'h001; 
        10'b0011101111: data <= 9'h001; 
        10'b0011110000: data <= 9'h001; 
        10'b0011110001: data <= 9'h002; 
        10'b0011110010: data <= 9'h001; 
        10'b0011110011: data <= 9'h001; 
        10'b0011110100: data <= 9'h001; 
        10'b0011110101: data <= 9'h000; 
        10'b0011110110: data <= 9'h001; 
        10'b0011110111: data <= 9'h001; 
        10'b0011111000: data <= 9'h000; 
        10'b0011111001: data <= 9'h000; 
        10'b0011111010: data <= 9'h000; 
        10'b0011111011: data <= 9'h000; 
        10'b0011111100: data <= 9'h000; 
        10'b0011111101: data <= 9'h000; 
        10'b0011111110: data <= 9'h000; 
        10'b0011111111: data <= 9'h001; 
        10'b0100000000: data <= 9'h001; 
        10'b0100000001: data <= 9'h001; 
        10'b0100000010: data <= 9'h000; 
        10'b0100000011: data <= 9'h001; 
        10'b0100000100: data <= 9'h001; 
        10'b0100000101: data <= 9'h000; 
        10'b0100000110: data <= 9'h001; 
        10'b0100000111: data <= 9'h001; 
        10'b0100001000: data <= 9'h002; 
        10'b0100001001: data <= 9'h002; 
        10'b0100001010: data <= 9'h002; 
        10'b0100001011: data <= 9'h003; 
        10'b0100001100: data <= 9'h002; 
        10'b0100001101: data <= 9'h003; 
        10'b0100001110: data <= 9'h002; 
        10'b0100001111: data <= 9'h002; 
        10'b0100010000: data <= 9'h002; 
        10'b0100010001: data <= 9'h001; 
        10'b0100010010: data <= 9'h001; 
        10'b0100010011: data <= 9'h000; 
        10'b0100010100: data <= 9'h000; 
        10'b0100010101: data <= 9'h000; 
        10'b0100010110: data <= 9'h000; 
        10'b0100010111: data <= 9'h000; 
        10'b0100011000: data <= 9'h000; 
        10'b0100011001: data <= 9'h000; 
        10'b0100011010: data <= 9'h000; 
        10'b0100011011: data <= 9'h001; 
        10'b0100011100: data <= 9'h001; 
        10'b0100011101: data <= 9'h001; 
        10'b0100011110: data <= 9'h000; 
        10'b0100011111: data <= 9'h000; 
        10'b0100100000: data <= 9'h000; 
        10'b0100100001: data <= 9'h000; 
        10'b0100100010: data <= 9'h001; 
        10'b0100100011: data <= 9'h001; 
        10'b0100100100: data <= 9'h001; 
        10'b0100100101: data <= 9'h002; 
        10'b0100100110: data <= 9'h003; 
        10'b0100100111: data <= 9'h003; 
        10'b0100101000: data <= 9'h004; 
        10'b0100101001: data <= 9'h003; 
        10'b0100101010: data <= 9'h002; 
        10'b0100101011: data <= 9'h002; 
        10'b0100101100: data <= 9'h002; 
        10'b0100101101: data <= 9'h002; 
        10'b0100101110: data <= 9'h001; 
        10'b0100101111: data <= 9'h000; 
        10'b0100110000: data <= 9'h1ff; 
        10'b0100110001: data <= 9'h000; 
        10'b0100110010: data <= 9'h000; 
        10'b0100110011: data <= 9'h000; 
        10'b0100110100: data <= 9'h000; 
        10'b0100110101: data <= 9'h000; 
        10'b0100110110: data <= 9'h000; 
        10'b0100110111: data <= 9'h001; 
        10'b0100111000: data <= 9'h001; 
        10'b0100111001: data <= 9'h001; 
        10'b0100111010: data <= 9'h000; 
        10'b0100111011: data <= 9'h000; 
        10'b0100111100: data <= 9'h000; 
        10'b0100111101: data <= 9'h001; 
        10'b0100111110: data <= 9'h000; 
        10'b0100111111: data <= 9'h001; 
        10'b0101000000: data <= 9'h001; 
        10'b0101000001: data <= 9'h001; 
        10'b0101000010: data <= 9'h001; 
        10'b0101000011: data <= 9'h003; 
        10'b0101000100: data <= 9'h003; 
        10'b0101000101: data <= 9'h002; 
        10'b0101000110: data <= 9'h002; 
        10'b0101000111: data <= 9'h002; 
        10'b0101001000: data <= 9'h002; 
        10'b0101001001: data <= 9'h001; 
        10'b0101001010: data <= 9'h001; 
        10'b0101001011: data <= 9'h000; 
        10'b0101001100: data <= 9'h1ff; 
        10'b0101001101: data <= 9'h000; 
        10'b0101001110: data <= 9'h000; 
        10'b0101001111: data <= 9'h000; 
        10'b0101010000: data <= 9'h000; 
        10'b0101010001: data <= 9'h000; 
        10'b0101010010: data <= 9'h000; 
        10'b0101010011: data <= 9'h001; 
        10'b0101010100: data <= 9'h001; 
        10'b0101010101: data <= 9'h000; 
        10'b0101010110: data <= 9'h000; 
        10'b0101010111: data <= 9'h001; 
        10'b0101011000: data <= 9'h001; 
        10'b0101011001: data <= 9'h000; 
        10'b0101011010: data <= 9'h1ff; 
        10'b0101011011: data <= 9'h1fe; 
        10'b0101011100: data <= 9'h1fd; 
        10'b0101011101: data <= 9'h1fb; 
        10'b0101011110: data <= 9'h1fc; 
        10'b0101011111: data <= 9'h000; 
        10'b0101100000: data <= 9'h002; 
        10'b0101100001: data <= 9'h002; 
        10'b0101100010: data <= 9'h001; 
        10'b0101100011: data <= 9'h000; 
        10'b0101100100: data <= 9'h000; 
        10'b0101100101: data <= 9'h000; 
        10'b0101100110: data <= 9'h000; 
        10'b0101100111: data <= 9'h000; 
        10'b0101101000: data <= 9'h000; 
        10'b0101101001: data <= 9'h000; 
        10'b0101101010: data <= 9'h000; 
        10'b0101101011: data <= 9'h000; 
        10'b0101101100: data <= 9'h000; 
        10'b0101101101: data <= 9'h000; 
        10'b0101101110: data <= 9'h000; 
        10'b0101101111: data <= 9'h001; 
        10'b0101110000: data <= 9'h000; 
        10'b0101110001: data <= 9'h000; 
        10'b0101110010: data <= 9'h000; 
        10'b0101110011: data <= 9'h000; 
        10'b0101110100: data <= 9'h000; 
        10'b0101110101: data <= 9'h1ff; 
        10'b0101110110: data <= 9'h1fe; 
        10'b0101110111: data <= 9'h1fc; 
        10'b0101111000: data <= 9'h1fa; 
        10'b0101111001: data <= 9'h1f9; 
        10'b0101111010: data <= 9'h1fc; 
        10'b0101111011: data <= 9'h000; 
        10'b0101111100: data <= 9'h001; 
        10'b0101111101: data <= 9'h001; 
        10'b0101111110: data <= 9'h000; 
        10'b0101111111: data <= 9'h000; 
        10'b0110000000: data <= 9'h1ff; 
        10'b0110000001: data <= 9'h1ff; 
        10'b0110000010: data <= 9'h000; 
        10'b0110000011: data <= 9'h000; 
        10'b0110000100: data <= 9'h000; 
        10'b0110000101: data <= 9'h000; 
        10'b0110000110: data <= 9'h000; 
        10'b0110000111: data <= 9'h000; 
        10'b0110001000: data <= 9'h000; 
        10'b0110001001: data <= 9'h000; 
        10'b0110001010: data <= 9'h001; 
        10'b0110001011: data <= 9'h001; 
        10'b0110001100: data <= 9'h000; 
        10'b0110001101: data <= 9'h001; 
        10'b0110001110: data <= 9'h000; 
        10'b0110001111: data <= 9'h000; 
        10'b0110010000: data <= 9'h1ff; 
        10'b0110010001: data <= 9'h1fe; 
        10'b0110010010: data <= 9'h1fd; 
        10'b0110010011: data <= 9'h1fc; 
        10'b0110010100: data <= 9'h1fb; 
        10'b0110010101: data <= 9'h1fb; 
        10'b0110010110: data <= 9'h1fe; 
        10'b0110010111: data <= 9'h000; 
        10'b0110011000: data <= 9'h000; 
        10'b0110011001: data <= 9'h001; 
        10'b0110011010: data <= 9'h002; 
        10'b0110011011: data <= 9'h002; 
        10'b0110011100: data <= 9'h001; 
        10'b0110011101: data <= 9'h001; 
        10'b0110011110: data <= 9'h001; 
        10'b0110011111: data <= 9'h001; 
        10'b0110100000: data <= 9'h000; 
        10'b0110100001: data <= 9'h000; 
        10'b0110100010: data <= 9'h000; 
        10'b0110100011: data <= 9'h000; 
        10'b0110100100: data <= 9'h000; 
        10'b0110100101: data <= 9'h000; 
        10'b0110100110: data <= 9'h000; 
        10'b0110100111: data <= 9'h000; 
        10'b0110101000: data <= 9'h000; 
        10'b0110101001: data <= 9'h1ff; 
        10'b0110101010: data <= 9'h000; 
        10'b0110101011: data <= 9'h000; 
        10'b0110101100: data <= 9'h1fe; 
        10'b0110101101: data <= 9'h1fe; 
        10'b0110101110: data <= 9'h1fd; 
        10'b0110101111: data <= 9'h1fc; 
        10'b0110110000: data <= 9'h1fc; 
        10'b0110110001: data <= 9'h1fd; 
        10'b0110110010: data <= 9'h1fe; 
        10'b0110110011: data <= 9'h000; 
        10'b0110110100: data <= 9'h000; 
        10'b0110110101: data <= 9'h003; 
        10'b0110110110: data <= 9'h003; 
        10'b0110110111: data <= 9'h003; 
        10'b0110111000: data <= 9'h002; 
        10'b0110111001: data <= 9'h002; 
        10'b0110111010: data <= 9'h001; 
        10'b0110111011: data <= 9'h001; 
        10'b0110111100: data <= 9'h000; 
        10'b0110111101: data <= 9'h000; 
        10'b0110111110: data <= 9'h000; 
        10'b0110111111: data <= 9'h000; 
        10'b0111000000: data <= 9'h000; 
        10'b0111000001: data <= 9'h000; 
        10'b0111000010: data <= 9'h000; 
        10'b0111000011: data <= 9'h000; 
        10'b0111000100: data <= 9'h000; 
        10'b0111000101: data <= 9'h000; 
        10'b0111000110: data <= 9'h000; 
        10'b0111000111: data <= 9'h000; 
        10'b0111001000: data <= 9'h1fe; 
        10'b0111001001: data <= 9'h1fe; 
        10'b0111001010: data <= 9'h1fd; 
        10'b0111001011: data <= 9'h1fd; 
        10'b0111001100: data <= 9'h1fe; 
        10'b0111001101: data <= 9'h1ff; 
        10'b0111001110: data <= 9'h1fe; 
        10'b0111001111: data <= 9'h001; 
        10'b0111010000: data <= 9'h001; 
        10'b0111010001: data <= 9'h002; 
        10'b0111010010: data <= 9'h002; 
        10'b0111010011: data <= 9'h002; 
        10'b0111010100: data <= 9'h002; 
        10'b0111010101: data <= 9'h001; 
        10'b0111010110: data <= 9'h000; 
        10'b0111010111: data <= 9'h1ff; 
        10'b0111011000: data <= 9'h000; 
        10'b0111011001: data <= 9'h000; 
        10'b0111011010: data <= 9'h000; 
        10'b0111011011: data <= 9'h000; 
        10'b0111011100: data <= 9'h000; 
        10'b0111011101: data <= 9'h000; 
        10'b0111011110: data <= 9'h000; 
        10'b0111011111: data <= 9'h000; 
        10'b0111100000: data <= 9'h000; 
        10'b0111100001: data <= 9'h000; 
        10'b0111100010: data <= 9'h1ff; 
        10'b0111100011: data <= 9'h1ff; 
        10'b0111100100: data <= 9'h1fe; 
        10'b0111100101: data <= 9'h1ff; 
        10'b0111100110: data <= 9'h1fe; 
        10'b0111100111: data <= 9'h1ff; 
        10'b0111101000: data <= 9'h000; 
        10'b0111101001: data <= 9'h000; 
        10'b0111101010: data <= 9'h000; 
        10'b0111101011: data <= 9'h000; 
        10'b0111101100: data <= 9'h000; 
        10'b0111101101: data <= 9'h001; 
        10'b0111101110: data <= 9'h001; 
        10'b0111101111: data <= 9'h000; 
        10'b0111110000: data <= 9'h000; 
        10'b0111110001: data <= 9'h000; 
        10'b0111110010: data <= 9'h1ff; 
        10'b0111110011: data <= 9'h000; 
        10'b0111110100: data <= 9'h000; 
        10'b0111110101: data <= 9'h000; 
        10'b0111110110: data <= 9'h000; 
        10'b0111110111: data <= 9'h000; 
        10'b0111111000: data <= 9'h000; 
        10'b0111111001: data <= 9'h000; 
        10'b0111111010: data <= 9'h000; 
        10'b0111111011: data <= 9'h000; 
        10'b0111111100: data <= 9'h000; 
        10'b0111111101: data <= 9'h1ff; 
        10'b0111111110: data <= 9'h1fe; 
        10'b0111111111: data <= 9'h1fe; 
        10'b1000000000: data <= 9'h1fe; 
        10'b1000000001: data <= 9'h1fe; 
        10'b1000000010: data <= 9'h1fe; 
        10'b1000000011: data <= 9'h1ff; 
        10'b1000000100: data <= 9'h000; 
        10'b1000000101: data <= 9'h000; 
        10'b1000000110: data <= 9'h001; 
        10'b1000000111: data <= 9'h1ff; 
        10'b1000001000: data <= 9'h1ff; 
        10'b1000001001: data <= 9'h000; 
        10'b1000001010: data <= 9'h1ff; 
        10'b1000001011: data <= 9'h1ff; 
        10'b1000001100: data <= 9'h1ff; 
        10'b1000001101: data <= 9'h1fe; 
        10'b1000001110: data <= 9'h1ff; 
        10'b1000001111: data <= 9'h1ff; 
        10'b1000010000: data <= 9'h1ff; 
        10'b1000010001: data <= 9'h000; 
        10'b1000010010: data <= 9'h000; 
        10'b1000010011: data <= 9'h000; 
        10'b1000010100: data <= 9'h000; 
        10'b1000010101: data <= 9'h000; 
        10'b1000010110: data <= 9'h000; 
        10'b1000010111: data <= 9'h000; 
        10'b1000011000: data <= 9'h000; 
        10'b1000011001: data <= 9'h1ff; 
        10'b1000011010: data <= 9'h1fe; 
        10'b1000011011: data <= 9'h1fe; 
        10'b1000011100: data <= 9'h1fe; 
        10'b1000011101: data <= 9'h1fe; 
        10'b1000011110: data <= 9'h1fe; 
        10'b1000011111: data <= 9'h1ff; 
        10'b1000100000: data <= 9'h1ff; 
        10'b1000100001: data <= 9'h000; 
        10'b1000100010: data <= 9'h001; 
        10'b1000100011: data <= 9'h1ff; 
        10'b1000100100: data <= 9'h1ff; 
        10'b1000100101: data <= 9'h1ff; 
        10'b1000100110: data <= 9'h1fe; 
        10'b1000100111: data <= 9'h1fe; 
        10'b1000101000: data <= 9'h1fe; 
        10'b1000101001: data <= 9'h1fe; 
        10'b1000101010: data <= 9'h1fe; 
        10'b1000101011: data <= 9'h1ff; 
        10'b1000101100: data <= 9'h1ff; 
        10'b1000101101: data <= 9'h000; 
        10'b1000101110: data <= 9'h000; 
        10'b1000101111: data <= 9'h000; 
        10'b1000110000: data <= 9'h000; 
        10'b1000110001: data <= 9'h000; 
        10'b1000110010: data <= 9'h000; 
        10'b1000110011: data <= 9'h000; 
        10'b1000110100: data <= 9'h000; 
        10'b1000110101: data <= 9'h1ff; 
        10'b1000110110: data <= 9'h1fe; 
        10'b1000110111: data <= 9'h1fe; 
        10'b1000111000: data <= 9'h1fe; 
        10'b1000111001: data <= 9'h1fe; 
        10'b1000111010: data <= 9'h1ff; 
        10'b1000111011: data <= 9'h1ff; 
        10'b1000111100: data <= 9'h000; 
        10'b1000111101: data <= 9'h000; 
        10'b1000111110: data <= 9'h001; 
        10'b1000111111: data <= 9'h1ff; 
        10'b1001000000: data <= 9'h1fe; 
        10'b1001000001: data <= 9'h1fe; 
        10'b1001000010: data <= 9'h1fd; 
        10'b1001000011: data <= 9'h1fe; 
        10'b1001000100: data <= 9'h1fd; 
        10'b1001000101: data <= 9'h1fe; 
        10'b1001000110: data <= 9'h1ff; 
        10'b1001000111: data <= 9'h1ff; 
        10'b1001001000: data <= 9'h000; 
        10'b1001001001: data <= 9'h000; 
        10'b1001001010: data <= 9'h000; 
        10'b1001001011: data <= 9'h000; 
        10'b1001001100: data <= 9'h000; 
        10'b1001001101: data <= 9'h000; 
        10'b1001001110: data <= 9'h000; 
        10'b1001001111: data <= 9'h000; 
        10'b1001010000: data <= 9'h000; 
        10'b1001010001: data <= 9'h1ff; 
        10'b1001010010: data <= 9'h1ff; 
        10'b1001010011: data <= 9'h1fe; 
        10'b1001010100: data <= 9'h1ff; 
        10'b1001010101: data <= 9'h1ff; 
        10'b1001010110: data <= 9'h1ff; 
        10'b1001010111: data <= 9'h1ff; 
        10'b1001011000: data <= 9'h000; 
        10'b1001011001: data <= 9'h000; 
        10'b1001011010: data <= 9'h000; 
        10'b1001011011: data <= 9'h1ff; 
        10'b1001011100: data <= 9'h1ff; 
        10'b1001011101: data <= 9'h1fe; 
        10'b1001011110: data <= 9'h1fe; 
        10'b1001011111: data <= 9'h1fe; 
        10'b1001100000: data <= 9'h1fe; 
        10'b1001100001: data <= 9'h1fe; 
        10'b1001100010: data <= 9'h1ff; 
        10'b1001100011: data <= 9'h1ff; 
        10'b1001100100: data <= 9'h000; 
        10'b1001100101: data <= 9'h000; 
        10'b1001100110: data <= 9'h000; 
        10'b1001100111: data <= 9'h000; 
        10'b1001101000: data <= 9'h000; 
        10'b1001101001: data <= 9'h000; 
        10'b1001101010: data <= 9'h000; 
        10'b1001101011: data <= 9'h000; 
        10'b1001101100: data <= 9'h000; 
        10'b1001101101: data <= 9'h000; 
        10'b1001101110: data <= 9'h000; 
        10'b1001101111: data <= 9'h000; 
        10'b1001110000: data <= 9'h000; 
        10'b1001110001: data <= 9'h000; 
        10'b1001110010: data <= 9'h1ff; 
        10'b1001110011: data <= 9'h1ff; 
        10'b1001110100: data <= 9'h1ff; 
        10'b1001110101: data <= 9'h1ff; 
        10'b1001110110: data <= 9'h000; 
        10'b1001110111: data <= 9'h000; 
        10'b1001111000: data <= 9'h1ff; 
        10'b1001111001: data <= 9'h1ff; 
        10'b1001111010: data <= 9'h1fe; 
        10'b1001111011: data <= 9'h1fe; 
        10'b1001111100: data <= 9'h1fe; 
        10'b1001111101: data <= 9'h1fe; 
        10'b1001111110: data <= 9'h1ff; 
        10'b1001111111: data <= 9'h000; 
        10'b1010000000: data <= 9'h000; 
        10'b1010000001: data <= 9'h000; 
        10'b1010000010: data <= 9'h000; 
        10'b1010000011: data <= 9'h000; 
        10'b1010000100: data <= 9'h000; 
        10'b1010000101: data <= 9'h000; 
        10'b1010000110: data <= 9'h000; 
        10'b1010000111: data <= 9'h000; 
        10'b1010001000: data <= 9'h000; 
        10'b1010001001: data <= 9'h000; 
        10'b1010001010: data <= 9'h001; 
        10'b1010001011: data <= 9'h001; 
        10'b1010001100: data <= 9'h001; 
        10'b1010001101: data <= 9'h000; 
        10'b1010001110: data <= 9'h000; 
        10'b1010001111: data <= 9'h1ff; 
        10'b1010010000: data <= 9'h1ff; 
        10'b1010010001: data <= 9'h000; 
        10'b1010010010: data <= 9'h001; 
        10'b1010010011: data <= 9'h000; 
        10'b1010010100: data <= 9'h000; 
        10'b1010010101: data <= 9'h000; 
        10'b1010010110: data <= 9'h1ff; 
        10'b1010010111: data <= 9'h1fe; 
        10'b1010011000: data <= 9'h1fe; 
        10'b1010011001: data <= 9'h1ff; 
        10'b1010011010: data <= 9'h1ff; 
        10'b1010011011: data <= 9'h1ff; 
        10'b1010011100: data <= 9'h000; 
        10'b1010011101: data <= 9'h000; 
        10'b1010011110: data <= 9'h000; 
        10'b1010011111: data <= 9'h000; 
        10'b1010100000: data <= 9'h000; 
        10'b1010100001: data <= 9'h000; 
        10'b1010100010: data <= 9'h000; 
        10'b1010100011: data <= 9'h000; 
        10'b1010100100: data <= 9'h000; 
        10'b1010100101: data <= 9'h001; 
        10'b1010100110: data <= 9'h002; 
        10'b1010100111: data <= 9'h002; 
        10'b1010101000: data <= 9'h002; 
        10'b1010101001: data <= 9'h001; 
        10'b1010101010: data <= 9'h002; 
        10'b1010101011: data <= 9'h001; 
        10'b1010101100: data <= 9'h001; 
        10'b1010101101: data <= 9'h001; 
        10'b1010101110: data <= 9'h001; 
        10'b1010101111: data <= 9'h001; 
        10'b1010110000: data <= 9'h001; 
        10'b1010110001: data <= 9'h001; 
        10'b1010110010: data <= 9'h000; 
        10'b1010110011: data <= 9'h000; 
        10'b1010110100: data <= 9'h1ff; 
        10'b1010110101: data <= 9'h1ff; 
        10'b1010110110: data <= 9'h1ff; 
        10'b1010110111: data <= 9'h1ff; 
        10'b1010111000: data <= 9'h000; 
        10'b1010111001: data <= 9'h000; 
        10'b1010111010: data <= 9'h000; 
        10'b1010111011: data <= 9'h000; 
        10'b1010111100: data <= 9'h000; 
        10'b1010111101: data <= 9'h000; 
        10'b1010111110: data <= 9'h000; 
        10'b1010111111: data <= 9'h000; 
        10'b1011000000: data <= 9'h000; 
        10'b1011000001: data <= 9'h001; 
        10'b1011000010: data <= 9'h001; 
        10'b1011000011: data <= 9'h001; 
        10'b1011000100: data <= 9'h002; 
        10'b1011000101: data <= 9'h002; 
        10'b1011000110: data <= 9'h002; 
        10'b1011000111: data <= 9'h002; 
        10'b1011001000: data <= 9'h002; 
        10'b1011001001: data <= 9'h002; 
        10'b1011001010: data <= 9'h002; 
        10'b1011001011: data <= 9'h002; 
        10'b1011001100: data <= 9'h001; 
        10'b1011001101: data <= 9'h001; 
        10'b1011001110: data <= 9'h001; 
        10'b1011001111: data <= 9'h000; 
        10'b1011010000: data <= 9'h000; 
        10'b1011010001: data <= 9'h000; 
        10'b1011010010: data <= 9'h000; 
        10'b1011010011: data <= 9'h000; 
        10'b1011010100: data <= 9'h000; 
        10'b1011010101: data <= 9'h000; 
        10'b1011010110: data <= 9'h000; 
        10'b1011010111: data <= 9'h000; 
        10'b1011011000: data <= 9'h000; 
        10'b1011011001: data <= 9'h000; 
        10'b1011011010: data <= 9'h000; 
        10'b1011011011: data <= 9'h000; 
        10'b1011011100: data <= 9'h000; 
        10'b1011011101: data <= 9'h000; 
        10'b1011011110: data <= 9'h000; 
        10'b1011011111: data <= 9'h000; 
        10'b1011100000: data <= 9'h000; 
        10'b1011100001: data <= 9'h000; 
        10'b1011100010: data <= 9'h000; 
        10'b1011100011: data <= 9'h001; 
        10'b1011100100: data <= 9'h000; 
        10'b1011100101: data <= 9'h001; 
        10'b1011100110: data <= 9'h001; 
        10'b1011100111: data <= 9'h001; 
        10'b1011101000: data <= 9'h001; 
        10'b1011101001: data <= 9'h001; 
        10'b1011101010: data <= 9'h001; 
        10'b1011101011: data <= 9'h000; 
        10'b1011101100: data <= 9'h000; 
        10'b1011101101: data <= 9'h000; 
        10'b1011101110: data <= 9'h000; 
        10'b1011101111: data <= 9'h000; 
        10'b1011110000: data <= 9'h000; 
        10'b1011110001: data <= 9'h000; 
        10'b1011110010: data <= 9'h000; 
        10'b1011110011: data <= 9'h000; 
        10'b1011110100: data <= 9'h000; 
        10'b1011110101: data <= 9'h000; 
        10'b1011110110: data <= 9'h000; 
        10'b1011110111: data <= 9'h000; 
        10'b1011111000: data <= 9'h000; 
        10'b1011111001: data <= 9'h000; 
        10'b1011111010: data <= 9'h000; 
        10'b1011111011: data <= 9'h000; 
        10'b1011111100: data <= 9'h000; 
        10'b1011111101: data <= 9'h000; 
        10'b1011111110: data <= 9'h000; 
        10'b1011111111: data <= 9'h000; 
        10'b1100000000: data <= 9'h000; 
        10'b1100000001: data <= 9'h000; 
        10'b1100000010: data <= 9'h000; 
        10'b1100000011: data <= 9'h000; 
        10'b1100000100: data <= 9'h001; 
        10'b1100000101: data <= 9'h000; 
        10'b1100000110: data <= 9'h000; 
        10'b1100000111: data <= 9'h000; 
        10'b1100001000: data <= 9'h000; 
        10'b1100001001: data <= 9'h000; 
        10'b1100001010: data <= 9'h000; 
        10'b1100001011: data <= 9'h000; 
        10'b1100001100: data <= 9'h000; 
        10'b1100001101: data <= 9'h000; 
        10'b1100001110: data <= 9'h000; 
        10'b1100001111: data <= 9'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 4) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 10'h000; 
        10'b0000000001: data <= 10'h000; 
        10'b0000000010: data <= 10'h000; 
        10'b0000000011: data <= 10'h000; 
        10'b0000000100: data <= 10'h001; 
        10'b0000000101: data <= 10'h000; 
        10'b0000000110: data <= 10'h000; 
        10'b0000000111: data <= 10'h000; 
        10'b0000001000: data <= 10'h001; 
        10'b0000001001: data <= 10'h001; 
        10'b0000001010: data <= 10'h000; 
        10'b0000001011: data <= 10'h000; 
        10'b0000001100: data <= 10'h000; 
        10'b0000001101: data <= 10'h000; 
        10'b0000001110: data <= 10'h001; 
        10'b0000001111: data <= 10'h000; 
        10'b0000010000: data <= 10'h000; 
        10'b0000010001: data <= 10'h000; 
        10'b0000010010: data <= 10'h000; 
        10'b0000010011: data <= 10'h000; 
        10'b0000010100: data <= 10'h000; 
        10'b0000010101: data <= 10'h001; 
        10'b0000010110: data <= 10'h000; 
        10'b0000010111: data <= 10'h001; 
        10'b0000011000: data <= 10'h000; 
        10'b0000011001: data <= 10'h000; 
        10'b0000011010: data <= 10'h000; 
        10'b0000011011: data <= 10'h000; 
        10'b0000011100: data <= 10'h001; 
        10'b0000011101: data <= 10'h000; 
        10'b0000011110: data <= 10'h000; 
        10'b0000011111: data <= 10'h001; 
        10'b0000100000: data <= 10'h000; 
        10'b0000100001: data <= 10'h000; 
        10'b0000100010: data <= 10'h001; 
        10'b0000100011: data <= 10'h000; 
        10'b0000100100: data <= 10'h000; 
        10'b0000100101: data <= 10'h000; 
        10'b0000100110: data <= 10'h000; 
        10'b0000100111: data <= 10'h000; 
        10'b0000101000: data <= 10'h001; 
        10'b0000101001: data <= 10'h000; 
        10'b0000101010: data <= 10'h001; 
        10'b0000101011: data <= 10'h000; 
        10'b0000101100: data <= 10'h000; 
        10'b0000101101: data <= 10'h001; 
        10'b0000101110: data <= 10'h001; 
        10'b0000101111: data <= 10'h000; 
        10'b0000110000: data <= 10'h000; 
        10'b0000110001: data <= 10'h000; 
        10'b0000110010: data <= 10'h000; 
        10'b0000110011: data <= 10'h001; 
        10'b0000110100: data <= 10'h001; 
        10'b0000110101: data <= 10'h000; 
        10'b0000110110: data <= 10'h000; 
        10'b0000110111: data <= 10'h000; 
        10'b0000111000: data <= 10'h001; 
        10'b0000111001: data <= 10'h001; 
        10'b0000111010: data <= 10'h001; 
        10'b0000111011: data <= 10'h000; 
        10'b0000111100: data <= 10'h001; 
        10'b0000111101: data <= 10'h000; 
        10'b0000111110: data <= 10'h000; 
        10'b0000111111: data <= 10'h000; 
        10'b0001000000: data <= 10'h000; 
        10'b0001000001: data <= 10'h000; 
        10'b0001000010: data <= 10'h000; 
        10'b0001000011: data <= 10'h000; 
        10'b0001000100: data <= 10'h000; 
        10'b0001000101: data <= 10'h000; 
        10'b0001000110: data <= 10'h000; 
        10'b0001000111: data <= 10'h001; 
        10'b0001001000: data <= 10'h000; 
        10'b0001001001: data <= 10'h000; 
        10'b0001001010: data <= 10'h000; 
        10'b0001001011: data <= 10'h001; 
        10'b0001001100: data <= 10'h001; 
        10'b0001001101: data <= 10'h001; 
        10'b0001001110: data <= 10'h000; 
        10'b0001001111: data <= 10'h001; 
        10'b0001010000: data <= 10'h000; 
        10'b0001010001: data <= 10'h000; 
        10'b0001010010: data <= 10'h000; 
        10'b0001010011: data <= 10'h001; 
        10'b0001010100: data <= 10'h000; 
        10'b0001010101: data <= 10'h000; 
        10'b0001010110: data <= 10'h001; 
        10'b0001010111: data <= 10'h000; 
        10'b0001011000: data <= 10'h000; 
        10'b0001011001: data <= 10'h000; 
        10'b0001011010: data <= 10'h000; 
        10'b0001011011: data <= 10'h000; 
        10'b0001011100: data <= 10'h000; 
        10'b0001011101: data <= 10'h000; 
        10'b0001011110: data <= 10'h000; 
        10'b0001011111: data <= 10'h000; 
        10'b0001100000: data <= 10'h000; 
        10'b0001100001: data <= 10'h000; 
        10'b0001100010: data <= 10'h000; 
        10'b0001100011: data <= 10'h000; 
        10'b0001100100: data <= 10'h3ff; 
        10'b0001100101: data <= 10'h3ff; 
        10'b0001100110: data <= 10'h000; 
        10'b0001100111: data <= 10'h000; 
        10'b0001101000: data <= 10'h000; 
        10'b0001101001: data <= 10'h000; 
        10'b0001101010: data <= 10'h000; 
        10'b0001101011: data <= 10'h000; 
        10'b0001101100: data <= 10'h000; 
        10'b0001101101: data <= 10'h001; 
        10'b0001101110: data <= 10'h000; 
        10'b0001101111: data <= 10'h000; 
        10'b0001110000: data <= 10'h001; 
        10'b0001110001: data <= 10'h000; 
        10'b0001110010: data <= 10'h000; 
        10'b0001110011: data <= 10'h000; 
        10'b0001110100: data <= 10'h000; 
        10'b0001110101: data <= 10'h000; 
        10'b0001110110: data <= 10'h000; 
        10'b0001110111: data <= 10'h000; 
        10'b0001111000: data <= 10'h000; 
        10'b0001111001: data <= 10'h000; 
        10'b0001111010: data <= 10'h3ff; 
        10'b0001111011: data <= 10'h3ff; 
        10'b0001111100: data <= 10'h3ff; 
        10'b0001111101: data <= 10'h3ff; 
        10'b0001111110: data <= 10'h3fe; 
        10'b0001111111: data <= 10'h3fd; 
        10'b0010000000: data <= 10'h3fe; 
        10'b0010000001: data <= 10'h3ff; 
        10'b0010000010: data <= 10'h3ff; 
        10'b0010000011: data <= 10'h000; 
        10'b0010000100: data <= 10'h3ff; 
        10'b0010000101: data <= 10'h000; 
        10'b0010000110: data <= 10'h000; 
        10'b0010000111: data <= 10'h000; 
        10'b0010001000: data <= 10'h001; 
        10'b0010001001: data <= 10'h000; 
        10'b0010001010: data <= 10'h001; 
        10'b0010001011: data <= 10'h001; 
        10'b0010001100: data <= 10'h001; 
        10'b0010001101: data <= 10'h000; 
        10'b0010001110: data <= 10'h001; 
        10'b0010001111: data <= 10'h000; 
        10'b0010010000: data <= 10'h000; 
        10'b0010010001: data <= 10'h000; 
        10'b0010010010: data <= 10'h000; 
        10'b0010010011: data <= 10'h000; 
        10'b0010010100: data <= 10'h000; 
        10'b0010010101: data <= 10'h3ff; 
        10'b0010010110: data <= 10'h3fe; 
        10'b0010010111: data <= 10'h3fd; 
        10'b0010011000: data <= 10'h3fc; 
        10'b0010011001: data <= 10'h3fc; 
        10'b0010011010: data <= 10'h3fa; 
        10'b0010011011: data <= 10'h3fa; 
        10'b0010011100: data <= 10'h3fa; 
        10'b0010011101: data <= 10'h3fb; 
        10'b0010011110: data <= 10'h3fc; 
        10'b0010011111: data <= 10'h3fd; 
        10'b0010100000: data <= 10'h3fe; 
        10'b0010100001: data <= 10'h3ff; 
        10'b0010100010: data <= 10'h3ff; 
        10'b0010100011: data <= 10'h000; 
        10'b0010100100: data <= 10'h001; 
        10'b0010100101: data <= 10'h000; 
        10'b0010100110: data <= 10'h000; 
        10'b0010100111: data <= 10'h000; 
        10'b0010101000: data <= 10'h001; 
        10'b0010101001: data <= 10'h001; 
        10'b0010101010: data <= 10'h000; 
        10'b0010101011: data <= 10'h000; 
        10'b0010101100: data <= 10'h001; 
        10'b0010101101: data <= 10'h001; 
        10'b0010101110: data <= 10'h001; 
        10'b0010101111: data <= 10'h002; 
        10'b0010110000: data <= 10'h002; 
        10'b0010110001: data <= 10'h002; 
        10'b0010110010: data <= 10'h002; 
        10'b0010110011: data <= 10'h000; 
        10'b0010110100: data <= 10'h3fe; 
        10'b0010110101: data <= 10'h3fd; 
        10'b0010110110: data <= 10'h3fc; 
        10'b0010110111: data <= 10'h3fe; 
        10'b0010111000: data <= 10'h3ff; 
        10'b0010111001: data <= 10'h3ff; 
        10'b0010111010: data <= 10'h3fe; 
        10'b0010111011: data <= 10'h3fe; 
        10'b0010111100: data <= 10'h3fd; 
        10'b0010111101: data <= 10'h3ff; 
        10'b0010111110: data <= 10'h3fe; 
        10'b0010111111: data <= 10'h3ff; 
        10'b0011000000: data <= 10'h3ff; 
        10'b0011000001: data <= 10'h000; 
        10'b0011000010: data <= 10'h000; 
        10'b0011000011: data <= 10'h000; 
        10'b0011000100: data <= 10'h000; 
        10'b0011000101: data <= 10'h001; 
        10'b0011000110: data <= 10'h001; 
        10'b0011000111: data <= 10'h001; 
        10'b0011001000: data <= 10'h002; 
        10'b0011001001: data <= 10'h002; 
        10'b0011001010: data <= 10'h002; 
        10'b0011001011: data <= 10'h003; 
        10'b0011001100: data <= 10'h005; 
        10'b0011001101: data <= 10'h004; 
        10'b0011001110: data <= 10'h003; 
        10'b0011001111: data <= 10'h003; 
        10'b0011010000: data <= 10'h003; 
        10'b0011010001: data <= 10'h001; 
        10'b0011010010: data <= 10'h000; 
        10'b0011010011: data <= 10'h001; 
        10'b0011010100: data <= 10'h003; 
        10'b0011010101: data <= 10'h003; 
        10'b0011010110: data <= 10'h002; 
        10'b0011010111: data <= 10'h002; 
        10'b0011011000: data <= 10'h000; 
        10'b0011011001: data <= 10'h3ff; 
        10'b0011011010: data <= 10'h000; 
        10'b0011011011: data <= 10'h3ff; 
        10'b0011011100: data <= 10'h3ff; 
        10'b0011011101: data <= 10'h000; 
        10'b0011011110: data <= 10'h000; 
        10'b0011011111: data <= 10'h000; 
        10'b0011100000: data <= 10'h000; 
        10'b0011100001: data <= 10'h001; 
        10'b0011100010: data <= 10'h000; 
        10'b0011100011: data <= 10'h001; 
        10'b0011100100: data <= 10'h002; 
        10'b0011100101: data <= 10'h002; 
        10'b0011100110: data <= 10'h003; 
        10'b0011100111: data <= 10'h005; 
        10'b0011101000: data <= 10'h004; 
        10'b0011101001: data <= 10'h002; 
        10'b0011101010: data <= 10'h003; 
        10'b0011101011: data <= 10'h004; 
        10'b0011101100: data <= 10'h004; 
        10'b0011101101: data <= 10'h002; 
        10'b0011101110: data <= 10'h001; 
        10'b0011101111: data <= 10'h002; 
        10'b0011110000: data <= 10'h003; 
        10'b0011110001: data <= 10'h004; 
        10'b0011110010: data <= 10'h003; 
        10'b0011110011: data <= 10'h003; 
        10'b0011110100: data <= 10'h002; 
        10'b0011110101: data <= 10'h000; 
        10'b0011110110: data <= 10'h001; 
        10'b0011110111: data <= 10'h001; 
        10'b0011111000: data <= 10'h3ff; 
        10'b0011111001: data <= 10'h000; 
        10'b0011111010: data <= 10'h000; 
        10'b0011111011: data <= 10'h001; 
        10'b0011111100: data <= 10'h000; 
        10'b0011111101: data <= 10'h001; 
        10'b0011111110: data <= 10'h001; 
        10'b0011111111: data <= 10'h002; 
        10'b0100000000: data <= 10'h002; 
        10'b0100000001: data <= 10'h003; 
        10'b0100000010: data <= 10'h001; 
        10'b0100000011: data <= 10'h001; 
        10'b0100000100: data <= 10'h001; 
        10'b0100000101: data <= 10'h001; 
        10'b0100000110: data <= 10'h002; 
        10'b0100000111: data <= 10'h003; 
        10'b0100001000: data <= 10'h004; 
        10'b0100001001: data <= 10'h003; 
        10'b0100001010: data <= 10'h004; 
        10'b0100001011: data <= 10'h005; 
        10'b0100001100: data <= 10'h005; 
        10'b0100001101: data <= 10'h006; 
        10'b0100001110: data <= 10'h004; 
        10'b0100001111: data <= 10'h004; 
        10'b0100010000: data <= 10'h003; 
        10'b0100010001: data <= 10'h003; 
        10'b0100010010: data <= 10'h001; 
        10'b0100010011: data <= 10'h000; 
        10'b0100010100: data <= 10'h3ff; 
        10'b0100010101: data <= 10'h000; 
        10'b0100010110: data <= 10'h000; 
        10'b0100010111: data <= 10'h000; 
        10'b0100011000: data <= 10'h000; 
        10'b0100011001: data <= 10'h001; 
        10'b0100011010: data <= 10'h001; 
        10'b0100011011: data <= 10'h002; 
        10'b0100011100: data <= 10'h002; 
        10'b0100011101: data <= 10'h002; 
        10'b0100011110: data <= 10'h000; 
        10'b0100011111: data <= 10'h001; 
        10'b0100100000: data <= 10'h3ff; 
        10'b0100100001: data <= 10'h000; 
        10'b0100100010: data <= 10'h001; 
        10'b0100100011: data <= 10'h003; 
        10'b0100100100: data <= 10'h002; 
        10'b0100100101: data <= 10'h004; 
        10'b0100100110: data <= 10'h005; 
        10'b0100100111: data <= 10'h007; 
        10'b0100101000: data <= 10'h008; 
        10'b0100101001: data <= 10'h006; 
        10'b0100101010: data <= 10'h004; 
        10'b0100101011: data <= 10'h005; 
        10'b0100101100: data <= 10'h004; 
        10'b0100101101: data <= 10'h003; 
        10'b0100101110: data <= 10'h002; 
        10'b0100101111: data <= 10'h3ff; 
        10'b0100110000: data <= 10'h3ff; 
        10'b0100110001: data <= 10'h000; 
        10'b0100110010: data <= 10'h000; 
        10'b0100110011: data <= 10'h000; 
        10'b0100110100: data <= 10'h001; 
        10'b0100110101: data <= 10'h000; 
        10'b0100110110: data <= 10'h001; 
        10'b0100110111: data <= 10'h002; 
        10'b0100111000: data <= 10'h003; 
        10'b0100111001: data <= 10'h001; 
        10'b0100111010: data <= 10'h000; 
        10'b0100111011: data <= 10'h000; 
        10'b0100111100: data <= 10'h000; 
        10'b0100111101: data <= 10'h002; 
        10'b0100111110: data <= 10'h001; 
        10'b0100111111: data <= 10'h001; 
        10'b0101000000: data <= 10'h002; 
        10'b0101000001: data <= 10'h002; 
        10'b0101000010: data <= 10'h002; 
        10'b0101000011: data <= 10'h005; 
        10'b0101000100: data <= 10'h007; 
        10'b0101000101: data <= 10'h004; 
        10'b0101000110: data <= 10'h004; 
        10'b0101000111: data <= 10'h003; 
        10'b0101001000: data <= 10'h003; 
        10'b0101001001: data <= 10'h002; 
        10'b0101001010: data <= 10'h002; 
        10'b0101001011: data <= 10'h3ff; 
        10'b0101001100: data <= 10'h3fe; 
        10'b0101001101: data <= 10'h000; 
        10'b0101001110: data <= 10'h000; 
        10'b0101001111: data <= 10'h001; 
        10'b0101010000: data <= 10'h001; 
        10'b0101010001: data <= 10'h000; 
        10'b0101010010: data <= 10'h000; 
        10'b0101010011: data <= 10'h001; 
        10'b0101010100: data <= 10'h002; 
        10'b0101010101: data <= 10'h000; 
        10'b0101010110: data <= 10'h000; 
        10'b0101010111: data <= 10'h001; 
        10'b0101011000: data <= 10'h001; 
        10'b0101011001: data <= 10'h000; 
        10'b0101011010: data <= 10'h3ff; 
        10'b0101011011: data <= 10'h3fd; 
        10'b0101011100: data <= 10'h3f9; 
        10'b0101011101: data <= 10'h3f6; 
        10'b0101011110: data <= 10'h3f8; 
        10'b0101011111: data <= 10'h000; 
        10'b0101100000: data <= 10'h004; 
        10'b0101100001: data <= 10'h004; 
        10'b0101100010: data <= 10'h002; 
        10'b0101100011: data <= 10'h001; 
        10'b0101100100: data <= 10'h000; 
        10'b0101100101: data <= 10'h3ff; 
        10'b0101100110: data <= 10'h3ff; 
        10'b0101100111: data <= 10'h3ff; 
        10'b0101101000: data <= 10'h3ff; 
        10'b0101101001: data <= 10'h001; 
        10'b0101101010: data <= 10'h000; 
        10'b0101101011: data <= 10'h000; 
        10'b0101101100: data <= 10'h001; 
        10'b0101101101: data <= 10'h000; 
        10'b0101101110: data <= 10'h001; 
        10'b0101101111: data <= 10'h001; 
        10'b0101110000: data <= 10'h000; 
        10'b0101110001: data <= 10'h000; 
        10'b0101110010: data <= 10'h000; 
        10'b0101110011: data <= 10'h000; 
        10'b0101110100: data <= 10'h000; 
        10'b0101110101: data <= 10'h3ff; 
        10'b0101110110: data <= 10'h3fd; 
        10'b0101110111: data <= 10'h3f9; 
        10'b0101111000: data <= 10'h3f4; 
        10'b0101111001: data <= 10'h3f2; 
        10'b0101111010: data <= 10'h3f9; 
        10'b0101111011: data <= 10'h3ff; 
        10'b0101111100: data <= 10'h002; 
        10'b0101111101: data <= 10'h001; 
        10'b0101111110: data <= 10'h000; 
        10'b0101111111: data <= 10'h001; 
        10'b0110000000: data <= 10'h3ff; 
        10'b0110000001: data <= 10'h3fe; 
        10'b0110000010: data <= 10'h000; 
        10'b0110000011: data <= 10'h000; 
        10'b0110000100: data <= 10'h000; 
        10'b0110000101: data <= 10'h000; 
        10'b0110000110: data <= 10'h000; 
        10'b0110000111: data <= 10'h000; 
        10'b0110001000: data <= 10'h000; 
        10'b0110001001: data <= 10'h000; 
        10'b0110001010: data <= 10'h001; 
        10'b0110001011: data <= 10'h001; 
        10'b0110001100: data <= 10'h001; 
        10'b0110001101: data <= 10'h001; 
        10'b0110001110: data <= 10'h000; 
        10'b0110001111: data <= 10'h3ff; 
        10'b0110010000: data <= 10'h3fe; 
        10'b0110010001: data <= 10'h3fc; 
        10'b0110010010: data <= 10'h3fb; 
        10'b0110010011: data <= 10'h3f8; 
        10'b0110010100: data <= 10'h3f5; 
        10'b0110010101: data <= 10'h3f7; 
        10'b0110010110: data <= 10'h3fd; 
        10'b0110010111: data <= 10'h000; 
        10'b0110011000: data <= 10'h001; 
        10'b0110011001: data <= 10'h001; 
        10'b0110011010: data <= 10'h004; 
        10'b0110011011: data <= 10'h004; 
        10'b0110011100: data <= 10'h003; 
        10'b0110011101: data <= 10'h002; 
        10'b0110011110: data <= 10'h002; 
        10'b0110011111: data <= 10'h001; 
        10'b0110100000: data <= 10'h001; 
        10'b0110100001: data <= 10'h000; 
        10'b0110100010: data <= 10'h000; 
        10'b0110100011: data <= 10'h000; 
        10'b0110100100: data <= 10'h000; 
        10'b0110100101: data <= 10'h001; 
        10'b0110100110: data <= 10'h000; 
        10'b0110100111: data <= 10'h001; 
        10'b0110101000: data <= 10'h001; 
        10'b0110101001: data <= 10'h3ff; 
        10'b0110101010: data <= 10'h3ff; 
        10'b0110101011: data <= 10'h3ff; 
        10'b0110101100: data <= 10'h3fc; 
        10'b0110101101: data <= 10'h3fb; 
        10'b0110101110: data <= 10'h3fa; 
        10'b0110101111: data <= 10'h3f9; 
        10'b0110110000: data <= 10'h3f8; 
        10'b0110110001: data <= 10'h3fa; 
        10'b0110110010: data <= 10'h3fd; 
        10'b0110110011: data <= 10'h000; 
        10'b0110110100: data <= 10'h000; 
        10'b0110110101: data <= 10'h006; 
        10'b0110110110: data <= 10'h007; 
        10'b0110110111: data <= 10'h005; 
        10'b0110111000: data <= 10'h005; 
        10'b0110111001: data <= 10'h004; 
        10'b0110111010: data <= 10'h003; 
        10'b0110111011: data <= 10'h001; 
        10'b0110111100: data <= 10'h000; 
        10'b0110111101: data <= 10'h000; 
        10'b0110111110: data <= 10'h000; 
        10'b0110111111: data <= 10'h001; 
        10'b0111000000: data <= 10'h000; 
        10'b0111000001: data <= 10'h001; 
        10'b0111000010: data <= 10'h000; 
        10'b0111000011: data <= 10'h001; 
        10'b0111000100: data <= 10'h001; 
        10'b0111000101: data <= 10'h3ff; 
        10'b0111000110: data <= 10'h3ff; 
        10'b0111000111: data <= 10'h000; 
        10'b0111001000: data <= 10'h3fd; 
        10'b0111001001: data <= 10'h3fc; 
        10'b0111001010: data <= 10'h3fa; 
        10'b0111001011: data <= 10'h3f9; 
        10'b0111001100: data <= 10'h3fc; 
        10'b0111001101: data <= 10'h3fe; 
        10'b0111001110: data <= 10'h3fd; 
        10'b0111001111: data <= 10'h002; 
        10'b0111010000: data <= 10'h002; 
        10'b0111010001: data <= 10'h005; 
        10'b0111010010: data <= 10'h004; 
        10'b0111010011: data <= 10'h004; 
        10'b0111010100: data <= 10'h003; 
        10'b0111010101: data <= 10'h003; 
        10'b0111010110: data <= 10'h001; 
        10'b0111010111: data <= 10'h3ff; 
        10'b0111011000: data <= 10'h3ff; 
        10'b0111011001: data <= 10'h000; 
        10'b0111011010: data <= 10'h000; 
        10'b0111011011: data <= 10'h001; 
        10'b0111011100: data <= 10'h000; 
        10'b0111011101: data <= 10'h000; 
        10'b0111011110: data <= 10'h000; 
        10'b0111011111: data <= 10'h000; 
        10'b0111100000: data <= 10'h000; 
        10'b0111100001: data <= 10'h000; 
        10'b0111100010: data <= 10'h3fe; 
        10'b0111100011: data <= 10'h3fd; 
        10'b0111100100: data <= 10'h3fc; 
        10'b0111100101: data <= 10'h3fd; 
        10'b0111100110: data <= 10'h3fc; 
        10'b0111100111: data <= 10'h3fd; 
        10'b0111101000: data <= 10'h3ff; 
        10'b0111101001: data <= 10'h001; 
        10'b0111101010: data <= 10'h000; 
        10'b0111101011: data <= 10'h001; 
        10'b0111101100: data <= 10'h000; 
        10'b0111101101: data <= 10'h001; 
        10'b0111101110: data <= 10'h001; 
        10'b0111101111: data <= 10'h001; 
        10'b0111110000: data <= 10'h000; 
        10'b0111110001: data <= 10'h3ff; 
        10'b0111110010: data <= 10'h3ff; 
        10'b0111110011: data <= 10'h3ff; 
        10'b0111110100: data <= 10'h3ff; 
        10'b0111110101: data <= 10'h000; 
        10'b0111110110: data <= 10'h000; 
        10'b0111110111: data <= 10'h000; 
        10'b0111111000: data <= 10'h000; 
        10'b0111111001: data <= 10'h000; 
        10'b0111111010: data <= 10'h000; 
        10'b0111111011: data <= 10'h000; 
        10'b0111111100: data <= 10'h3ff; 
        10'b0111111101: data <= 10'h3fe; 
        10'b0111111110: data <= 10'h3fd; 
        10'b0111111111: data <= 10'h3fc; 
        10'b1000000000: data <= 10'h3fc; 
        10'b1000000001: data <= 10'h3fc; 
        10'b1000000010: data <= 10'h3fb; 
        10'b1000000011: data <= 10'h3fe; 
        10'b1000000100: data <= 10'h000; 
        10'b1000000101: data <= 10'h000; 
        10'b1000000110: data <= 10'h001; 
        10'b1000000111: data <= 10'h3ff; 
        10'b1000001000: data <= 10'h3fe; 
        10'b1000001001: data <= 10'h3ff; 
        10'b1000001010: data <= 10'h3fe; 
        10'b1000001011: data <= 10'h3ff; 
        10'b1000001100: data <= 10'h3fe; 
        10'b1000001101: data <= 10'h3fd; 
        10'b1000001110: data <= 10'h3fd; 
        10'b1000001111: data <= 10'h3fe; 
        10'b1000010000: data <= 10'h3ff; 
        10'b1000010001: data <= 10'h000; 
        10'b1000010010: data <= 10'h000; 
        10'b1000010011: data <= 10'h000; 
        10'b1000010100: data <= 10'h001; 
        10'b1000010101: data <= 10'h001; 
        10'b1000010110: data <= 10'h001; 
        10'b1000010111: data <= 10'h000; 
        10'b1000011000: data <= 10'h3ff; 
        10'b1000011001: data <= 10'h3fd; 
        10'b1000011010: data <= 10'h3fc; 
        10'b1000011011: data <= 10'h3fb; 
        10'b1000011100: data <= 10'h3fb; 
        10'b1000011101: data <= 10'h3fb; 
        10'b1000011110: data <= 10'h3fd; 
        10'b1000011111: data <= 10'h3fe; 
        10'b1000100000: data <= 10'h3ff; 
        10'b1000100001: data <= 10'h001; 
        10'b1000100010: data <= 10'h002; 
        10'b1000100011: data <= 10'h3fe; 
        10'b1000100100: data <= 10'h3fe; 
        10'b1000100101: data <= 10'h3fe; 
        10'b1000100110: data <= 10'h3fc; 
        10'b1000100111: data <= 10'h3fc; 
        10'b1000101000: data <= 10'h3fb; 
        10'b1000101001: data <= 10'h3fc; 
        10'b1000101010: data <= 10'h3fd; 
        10'b1000101011: data <= 10'h3fe; 
        10'b1000101100: data <= 10'h3ff; 
        10'b1000101101: data <= 10'h000; 
        10'b1000101110: data <= 10'h001; 
        10'b1000101111: data <= 10'h000; 
        10'b1000110000: data <= 10'h000; 
        10'b1000110001: data <= 10'h000; 
        10'b1000110010: data <= 10'h000; 
        10'b1000110011: data <= 10'h000; 
        10'b1000110100: data <= 10'h3ff; 
        10'b1000110101: data <= 10'h3fe; 
        10'b1000110110: data <= 10'h3fc; 
        10'b1000110111: data <= 10'h3fb; 
        10'b1000111000: data <= 10'h3fc; 
        10'b1000111001: data <= 10'h3fc; 
        10'b1000111010: data <= 10'h3fd; 
        10'b1000111011: data <= 10'h3fd; 
        10'b1000111100: data <= 10'h000; 
        10'b1000111101: data <= 10'h000; 
        10'b1000111110: data <= 10'h001; 
        10'b1000111111: data <= 10'h3fd; 
        10'b1001000000: data <= 10'h3fd; 
        10'b1001000001: data <= 10'h3fc; 
        10'b1001000010: data <= 10'h3fa; 
        10'b1001000011: data <= 10'h3fc; 
        10'b1001000100: data <= 10'h3fb; 
        10'b1001000101: data <= 10'h3fc; 
        10'b1001000110: data <= 10'h3fd; 
        10'b1001000111: data <= 10'h3ff; 
        10'b1001001000: data <= 10'h3ff; 
        10'b1001001001: data <= 10'h001; 
        10'b1001001010: data <= 10'h001; 
        10'b1001001011: data <= 10'h000; 
        10'b1001001100: data <= 10'h001; 
        10'b1001001101: data <= 10'h001; 
        10'b1001001110: data <= 10'h000; 
        10'b1001001111: data <= 10'h3ff; 
        10'b1001010000: data <= 10'h000; 
        10'b1001010001: data <= 10'h3fe; 
        10'b1001010010: data <= 10'h3fe; 
        10'b1001010011: data <= 10'h3fd; 
        10'b1001010100: data <= 10'h3fd; 
        10'b1001010101: data <= 10'h3fe; 
        10'b1001010110: data <= 10'h3fe; 
        10'b1001010111: data <= 10'h3fe; 
        10'b1001011000: data <= 10'h3ff; 
        10'b1001011001: data <= 10'h000; 
        10'b1001011010: data <= 10'h3ff; 
        10'b1001011011: data <= 10'h3fe; 
        10'b1001011100: data <= 10'h3fe; 
        10'b1001011101: data <= 10'h3fc; 
        10'b1001011110: data <= 10'h3fc; 
        10'b1001011111: data <= 10'h3fc; 
        10'b1001100000: data <= 10'h3fc; 
        10'b1001100001: data <= 10'h3fc; 
        10'b1001100010: data <= 10'h3fe; 
        10'b1001100011: data <= 10'h3fe; 
        10'b1001100100: data <= 10'h000; 
        10'b1001100101: data <= 10'h000; 
        10'b1001100110: data <= 10'h001; 
        10'b1001100111: data <= 10'h000; 
        10'b1001101000: data <= 10'h000; 
        10'b1001101001: data <= 10'h000; 
        10'b1001101010: data <= 10'h000; 
        10'b1001101011: data <= 10'h000; 
        10'b1001101100: data <= 10'h000; 
        10'b1001101101: data <= 10'h000; 
        10'b1001101110: data <= 10'h3ff; 
        10'b1001101111: data <= 10'h000; 
        10'b1001110000: data <= 10'h001; 
        10'b1001110001: data <= 10'h3ff; 
        10'b1001110010: data <= 10'h3fe; 
        10'b1001110011: data <= 10'h3fd; 
        10'b1001110100: data <= 10'h3fd; 
        10'b1001110101: data <= 10'h3ff; 
        10'b1001110110: data <= 10'h000; 
        10'b1001110111: data <= 10'h000; 
        10'b1001111000: data <= 10'h3fe; 
        10'b1001111001: data <= 10'h3fe; 
        10'b1001111010: data <= 10'h3fd; 
        10'b1001111011: data <= 10'h3fd; 
        10'b1001111100: data <= 10'h3fc; 
        10'b1001111101: data <= 10'h3fd; 
        10'b1001111110: data <= 10'h3fe; 
        10'b1001111111: data <= 10'h3ff; 
        10'b1010000000: data <= 10'h000; 
        10'b1010000001: data <= 10'h000; 
        10'b1010000010: data <= 10'h000; 
        10'b1010000011: data <= 10'h000; 
        10'b1010000100: data <= 10'h000; 
        10'b1010000101: data <= 10'h001; 
        10'b1010000110: data <= 10'h000; 
        10'b1010000111: data <= 10'h000; 
        10'b1010001000: data <= 10'h001; 
        10'b1010001001: data <= 10'h001; 
        10'b1010001010: data <= 10'h002; 
        10'b1010001011: data <= 10'h003; 
        10'b1010001100: data <= 10'h001; 
        10'b1010001101: data <= 10'h000; 
        10'b1010001110: data <= 10'h3ff; 
        10'b1010001111: data <= 10'h3fe; 
        10'b1010010000: data <= 10'h3fe; 
        10'b1010010001: data <= 10'h000; 
        10'b1010010010: data <= 10'h001; 
        10'b1010010011: data <= 10'h001; 
        10'b1010010100: data <= 10'h000; 
        10'b1010010101: data <= 10'h3ff; 
        10'b1010010110: data <= 10'h3fe; 
        10'b1010010111: data <= 10'h3fd; 
        10'b1010011000: data <= 10'h3fd; 
        10'b1010011001: data <= 10'h3fe; 
        10'b1010011010: data <= 10'h3fe; 
        10'b1010011011: data <= 10'h3ff; 
        10'b1010011100: data <= 10'h3ff; 
        10'b1010011101: data <= 10'h000; 
        10'b1010011110: data <= 10'h000; 
        10'b1010011111: data <= 10'h000; 
        10'b1010100000: data <= 10'h000; 
        10'b1010100001: data <= 10'h000; 
        10'b1010100010: data <= 10'h000; 
        10'b1010100011: data <= 10'h000; 
        10'b1010100100: data <= 10'h001; 
        10'b1010100101: data <= 10'h002; 
        10'b1010100110: data <= 10'h003; 
        10'b1010100111: data <= 10'h004; 
        10'b1010101000: data <= 10'h003; 
        10'b1010101001: data <= 10'h002; 
        10'b1010101010: data <= 10'h004; 
        10'b1010101011: data <= 10'h002; 
        10'b1010101100: data <= 10'h002; 
        10'b1010101101: data <= 10'h003; 
        10'b1010101110: data <= 10'h002; 
        10'b1010101111: data <= 10'h002; 
        10'b1010110000: data <= 10'h001; 
        10'b1010110001: data <= 10'h001; 
        10'b1010110010: data <= 10'h000; 
        10'b1010110011: data <= 10'h3ff; 
        10'b1010110100: data <= 10'h3ff; 
        10'b1010110101: data <= 10'h3ff; 
        10'b1010110110: data <= 10'h3ff; 
        10'b1010110111: data <= 10'h3ff; 
        10'b1010111000: data <= 10'h000; 
        10'b1010111001: data <= 10'h000; 
        10'b1010111010: data <= 10'h000; 
        10'b1010111011: data <= 10'h000; 
        10'b1010111100: data <= 10'h000; 
        10'b1010111101: data <= 10'h000; 
        10'b1010111110: data <= 10'h001; 
        10'b1010111111: data <= 10'h001; 
        10'b1011000000: data <= 10'h000; 
        10'b1011000001: data <= 10'h001; 
        10'b1011000010: data <= 10'h002; 
        10'b1011000011: data <= 10'h003; 
        10'b1011000100: data <= 10'h004; 
        10'b1011000101: data <= 10'h004; 
        10'b1011000110: data <= 10'h005; 
        10'b1011000111: data <= 10'h004; 
        10'b1011001000: data <= 10'h004; 
        10'b1011001001: data <= 10'h003; 
        10'b1011001010: data <= 10'h003; 
        10'b1011001011: data <= 10'h003; 
        10'b1011001100: data <= 10'h003; 
        10'b1011001101: data <= 10'h003; 
        10'b1011001110: data <= 10'h002; 
        10'b1011001111: data <= 10'h001; 
        10'b1011010000: data <= 10'h3ff; 
        10'b1011010001: data <= 10'h000; 
        10'b1011010010: data <= 10'h000; 
        10'b1011010011: data <= 10'h000; 
        10'b1011010100: data <= 10'h000; 
        10'b1011010101: data <= 10'h000; 
        10'b1011010110: data <= 10'h001; 
        10'b1011010111: data <= 10'h001; 
        10'b1011011000: data <= 10'h000; 
        10'b1011011001: data <= 10'h000; 
        10'b1011011010: data <= 10'h001; 
        10'b1011011011: data <= 10'h000; 
        10'b1011011100: data <= 10'h000; 
        10'b1011011101: data <= 10'h001; 
        10'b1011011110: data <= 10'h000; 
        10'b1011011111: data <= 10'h001; 
        10'b1011100000: data <= 10'h001; 
        10'b1011100001: data <= 10'h000; 
        10'b1011100010: data <= 10'h001; 
        10'b1011100011: data <= 10'h001; 
        10'b1011100100: data <= 10'h000; 
        10'b1011100101: data <= 10'h001; 
        10'b1011100110: data <= 10'h002; 
        10'b1011100111: data <= 10'h003; 
        10'b1011101000: data <= 10'h002; 
        10'b1011101001: data <= 10'h003; 
        10'b1011101010: data <= 10'h002; 
        10'b1011101011: data <= 10'h001; 
        10'b1011101100: data <= 10'h000; 
        10'b1011101101: data <= 10'h000; 
        10'b1011101110: data <= 10'h000; 
        10'b1011101111: data <= 10'h000; 
        10'b1011110000: data <= 10'h000; 
        10'b1011110001: data <= 10'h000; 
        10'b1011110010: data <= 10'h000; 
        10'b1011110011: data <= 10'h000; 
        10'b1011110100: data <= 10'h000; 
        10'b1011110101: data <= 10'h000; 
        10'b1011110110: data <= 10'h000; 
        10'b1011110111: data <= 10'h000; 
        10'b1011111000: data <= 10'h001; 
        10'b1011111001: data <= 10'h000; 
        10'b1011111010: data <= 10'h000; 
        10'b1011111011: data <= 10'h000; 
        10'b1011111100: data <= 10'h001; 
        10'b1011111101: data <= 10'h001; 
        10'b1011111110: data <= 10'h000; 
        10'b1011111111: data <= 10'h001; 
        10'b1100000000: data <= 10'h000; 
        10'b1100000001: data <= 10'h001; 
        10'b1100000010: data <= 10'h001; 
        10'b1100000011: data <= 10'h000; 
        10'b1100000100: data <= 10'h001; 
        10'b1100000101: data <= 10'h000; 
        10'b1100000110: data <= 10'h000; 
        10'b1100000111: data <= 10'h001; 
        10'b1100001000: data <= 10'h000; 
        10'b1100001001: data <= 10'h000; 
        10'b1100001010: data <= 10'h001; 
        10'b1100001011: data <= 10'h000; 
        10'b1100001100: data <= 10'h000; 
        10'b1100001101: data <= 10'h000; 
        10'b1100001110: data <= 10'h000; 
        10'b1100001111: data <= 10'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 5) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 11'h000; 
        10'b0000000001: data <= 11'h000; 
        10'b0000000010: data <= 11'h001; 
        10'b0000000011: data <= 11'h000; 
        10'b0000000100: data <= 11'h002; 
        10'b0000000101: data <= 11'h7ff; 
        10'b0000000110: data <= 11'h000; 
        10'b0000000111: data <= 11'h001; 
        10'b0000001000: data <= 11'h001; 
        10'b0000001001: data <= 11'h001; 
        10'b0000001010: data <= 11'h7ff; 
        10'b0000001011: data <= 11'h000; 
        10'b0000001100: data <= 11'h000; 
        10'b0000001101: data <= 11'h000; 
        10'b0000001110: data <= 11'h001; 
        10'b0000001111: data <= 11'h000; 
        10'b0000010000: data <= 11'h000; 
        10'b0000010001: data <= 11'h000; 
        10'b0000010010: data <= 11'h000; 
        10'b0000010011: data <= 11'h000; 
        10'b0000010100: data <= 11'h001; 
        10'b0000010101: data <= 11'h002; 
        10'b0000010110: data <= 11'h000; 
        10'b0000010111: data <= 11'h001; 
        10'b0000011000: data <= 11'h000; 
        10'b0000011001: data <= 11'h001; 
        10'b0000011010: data <= 11'h000; 
        10'b0000011011: data <= 11'h000; 
        10'b0000011100: data <= 11'h001; 
        10'b0000011101: data <= 11'h000; 
        10'b0000011110: data <= 11'h000; 
        10'b0000011111: data <= 11'h001; 
        10'b0000100000: data <= 11'h001; 
        10'b0000100001: data <= 11'h000; 
        10'b0000100010: data <= 11'h001; 
        10'b0000100011: data <= 11'h000; 
        10'b0000100100: data <= 11'h000; 
        10'b0000100101: data <= 11'h000; 
        10'b0000100110: data <= 11'h000; 
        10'b0000100111: data <= 11'h7ff; 
        10'b0000101000: data <= 11'h001; 
        10'b0000101001: data <= 11'h000; 
        10'b0000101010: data <= 11'h001; 
        10'b0000101011: data <= 11'h000; 
        10'b0000101100: data <= 11'h001; 
        10'b0000101101: data <= 11'h001; 
        10'b0000101110: data <= 11'h001; 
        10'b0000101111: data <= 11'h001; 
        10'b0000110000: data <= 11'h000; 
        10'b0000110001: data <= 11'h001; 
        10'b0000110010: data <= 11'h000; 
        10'b0000110011: data <= 11'h002; 
        10'b0000110100: data <= 11'h001; 
        10'b0000110101: data <= 11'h000; 
        10'b0000110110: data <= 11'h000; 
        10'b0000110111: data <= 11'h001; 
        10'b0000111000: data <= 11'h001; 
        10'b0000111001: data <= 11'h001; 
        10'b0000111010: data <= 11'h001; 
        10'b0000111011: data <= 11'h000; 
        10'b0000111100: data <= 11'h001; 
        10'b0000111101: data <= 11'h7ff; 
        10'b0000111110: data <= 11'h000; 
        10'b0000111111: data <= 11'h001; 
        10'b0001000000: data <= 11'h001; 
        10'b0001000001: data <= 11'h000; 
        10'b0001000010: data <= 11'h000; 
        10'b0001000011: data <= 11'h001; 
        10'b0001000100: data <= 11'h000; 
        10'b0001000101: data <= 11'h000; 
        10'b0001000110: data <= 11'h000; 
        10'b0001000111: data <= 11'h001; 
        10'b0001001000: data <= 11'h001; 
        10'b0001001001: data <= 11'h000; 
        10'b0001001010: data <= 11'h000; 
        10'b0001001011: data <= 11'h001; 
        10'b0001001100: data <= 11'h001; 
        10'b0001001101: data <= 11'h001; 
        10'b0001001110: data <= 11'h7ff; 
        10'b0001001111: data <= 11'h001; 
        10'b0001010000: data <= 11'h000; 
        10'b0001010001: data <= 11'h001; 
        10'b0001010010: data <= 11'h001; 
        10'b0001010011: data <= 11'h001; 
        10'b0001010100: data <= 11'h000; 
        10'b0001010101: data <= 11'h000; 
        10'b0001010110: data <= 11'h001; 
        10'b0001010111: data <= 11'h000; 
        10'b0001011000: data <= 11'h000; 
        10'b0001011001: data <= 11'h000; 
        10'b0001011010: data <= 11'h000; 
        10'b0001011011: data <= 11'h001; 
        10'b0001011100: data <= 11'h000; 
        10'b0001011101: data <= 11'h001; 
        10'b0001011110: data <= 11'h7ff; 
        10'b0001011111: data <= 11'h000; 
        10'b0001100000: data <= 11'h001; 
        10'b0001100001: data <= 11'h7ff; 
        10'b0001100010: data <= 11'h001; 
        10'b0001100011: data <= 11'h7ff; 
        10'b0001100100: data <= 11'h7ff; 
        10'b0001100101: data <= 11'h7ff; 
        10'b0001100110: data <= 11'h7ff; 
        10'b0001100111: data <= 11'h7ff; 
        10'b0001101000: data <= 11'h000; 
        10'b0001101001: data <= 11'h7ff; 
        10'b0001101010: data <= 11'h000; 
        10'b0001101011: data <= 11'h000; 
        10'b0001101100: data <= 11'h001; 
        10'b0001101101: data <= 11'h002; 
        10'b0001101110: data <= 11'h7ff; 
        10'b0001101111: data <= 11'h001; 
        10'b0001110000: data <= 11'h001; 
        10'b0001110001: data <= 11'h7ff; 
        10'b0001110010: data <= 11'h001; 
        10'b0001110011: data <= 11'h7ff; 
        10'b0001110100: data <= 11'h000; 
        10'b0001110101: data <= 11'h000; 
        10'b0001110110: data <= 11'h000; 
        10'b0001110111: data <= 11'h7ff; 
        10'b0001111000: data <= 11'h000; 
        10'b0001111001: data <= 11'h000; 
        10'b0001111010: data <= 11'h7ff; 
        10'b0001111011: data <= 11'h7fd; 
        10'b0001111100: data <= 11'h7fd; 
        10'b0001111101: data <= 11'h7fd; 
        10'b0001111110: data <= 11'h7fd; 
        10'b0001111111: data <= 11'h7fb; 
        10'b0010000000: data <= 11'h7fd; 
        10'b0010000001: data <= 11'h7fe; 
        10'b0010000010: data <= 11'h7fe; 
        10'b0010000011: data <= 11'h7ff; 
        10'b0010000100: data <= 11'h7fe; 
        10'b0010000101: data <= 11'h001; 
        10'b0010000110: data <= 11'h000; 
        10'b0010000111: data <= 11'h7ff; 
        10'b0010001000: data <= 11'h001; 
        10'b0010001001: data <= 11'h000; 
        10'b0010001010: data <= 11'h001; 
        10'b0010001011: data <= 11'h001; 
        10'b0010001100: data <= 11'h001; 
        10'b0010001101: data <= 11'h000; 
        10'b0010001110: data <= 11'h001; 
        10'b0010001111: data <= 11'h000; 
        10'b0010010000: data <= 11'h7ff; 
        10'b0010010001: data <= 11'h000; 
        10'b0010010010: data <= 11'h7ff; 
        10'b0010010011: data <= 11'h000; 
        10'b0010010100: data <= 11'h7ff; 
        10'b0010010101: data <= 11'h7fe; 
        10'b0010010110: data <= 11'h7fb; 
        10'b0010010111: data <= 11'h7fa; 
        10'b0010011000: data <= 11'h7f8; 
        10'b0010011001: data <= 11'h7f7; 
        10'b0010011010: data <= 11'h7f5; 
        10'b0010011011: data <= 11'h7f5; 
        10'b0010011100: data <= 11'h7f4; 
        10'b0010011101: data <= 11'h7f6; 
        10'b0010011110: data <= 11'h7f7; 
        10'b0010011111: data <= 11'h7f9; 
        10'b0010100000: data <= 11'h7fb; 
        10'b0010100001: data <= 11'h7fe; 
        10'b0010100010: data <= 11'h7fd; 
        10'b0010100011: data <= 11'h000; 
        10'b0010100100: data <= 11'h001; 
        10'b0010100101: data <= 11'h001; 
        10'b0010100110: data <= 11'h000; 
        10'b0010100111: data <= 11'h000; 
        10'b0010101000: data <= 11'h001; 
        10'b0010101001: data <= 11'h001; 
        10'b0010101010: data <= 11'h000; 
        10'b0010101011: data <= 11'h000; 
        10'b0010101100: data <= 11'h002; 
        10'b0010101101: data <= 11'h002; 
        10'b0010101110: data <= 11'h002; 
        10'b0010101111: data <= 11'h003; 
        10'b0010110000: data <= 11'h005; 
        10'b0010110001: data <= 11'h004; 
        10'b0010110010: data <= 11'h004; 
        10'b0010110011: data <= 11'h001; 
        10'b0010110100: data <= 11'h7fd; 
        10'b0010110101: data <= 11'h7f9; 
        10'b0010110110: data <= 11'h7f9; 
        10'b0010110111: data <= 11'h7fc; 
        10'b0010111000: data <= 11'h7fe; 
        10'b0010111001: data <= 11'h7fd; 
        10'b0010111010: data <= 11'h7fd; 
        10'b0010111011: data <= 11'h7fc; 
        10'b0010111100: data <= 11'h7fa; 
        10'b0010111101: data <= 11'h7fe; 
        10'b0010111110: data <= 11'h7fc; 
        10'b0010111111: data <= 11'h7fd; 
        10'b0011000000: data <= 11'h7fe; 
        10'b0011000001: data <= 11'h7ff; 
        10'b0011000010: data <= 11'h7ff; 
        10'b0011000011: data <= 11'h000; 
        10'b0011000100: data <= 11'h001; 
        10'b0011000101: data <= 11'h001; 
        10'b0011000110: data <= 11'h001; 
        10'b0011000111: data <= 11'h003; 
        10'b0011001000: data <= 11'h003; 
        10'b0011001001: data <= 11'h003; 
        10'b0011001010: data <= 11'h004; 
        10'b0011001011: data <= 11'h007; 
        10'b0011001100: data <= 11'h009; 
        10'b0011001101: data <= 11'h007; 
        10'b0011001110: data <= 11'h005; 
        10'b0011001111: data <= 11'h006; 
        10'b0011010000: data <= 11'h006; 
        10'b0011010001: data <= 11'h001; 
        10'b0011010010: data <= 11'h001; 
        10'b0011010011: data <= 11'h002; 
        10'b0011010100: data <= 11'h006; 
        10'b0011010101: data <= 11'h007; 
        10'b0011010110: data <= 11'h005; 
        10'b0011010111: data <= 11'h004; 
        10'b0011011000: data <= 11'h001; 
        10'b0011011001: data <= 11'h7ff; 
        10'b0011011010: data <= 11'h000; 
        10'b0011011011: data <= 11'h7ff; 
        10'b0011011100: data <= 11'h7ff; 
        10'b0011011101: data <= 11'h000; 
        10'b0011011110: data <= 11'h001; 
        10'b0011011111: data <= 11'h000; 
        10'b0011100000: data <= 11'h7ff; 
        10'b0011100001: data <= 11'h002; 
        10'b0011100010: data <= 11'h001; 
        10'b0011100011: data <= 11'h002; 
        10'b0011100100: data <= 11'h005; 
        10'b0011100101: data <= 11'h004; 
        10'b0011100110: data <= 11'h006; 
        10'b0011100111: data <= 11'h00a; 
        10'b0011101000: data <= 11'h007; 
        10'b0011101001: data <= 11'h005; 
        10'b0011101010: data <= 11'h006; 
        10'b0011101011: data <= 11'h008; 
        10'b0011101100: data <= 11'h008; 
        10'b0011101101: data <= 11'h004; 
        10'b0011101110: data <= 11'h002; 
        10'b0011101111: data <= 11'h003; 
        10'b0011110000: data <= 11'h006; 
        10'b0011110001: data <= 11'h009; 
        10'b0011110010: data <= 11'h006; 
        10'b0011110011: data <= 11'h005; 
        10'b0011110100: data <= 11'h004; 
        10'b0011110101: data <= 11'h000; 
        10'b0011110110: data <= 11'h002; 
        10'b0011110111: data <= 11'h002; 
        10'b0011111000: data <= 11'h7ff; 
        10'b0011111001: data <= 11'h7ff; 
        10'b0011111010: data <= 11'h001; 
        10'b0011111011: data <= 11'h001; 
        10'b0011111100: data <= 11'h001; 
        10'b0011111101: data <= 11'h001; 
        10'b0011111110: data <= 11'h002; 
        10'b0011111111: data <= 11'h003; 
        10'b0100000000: data <= 11'h005; 
        10'b0100000001: data <= 11'h005; 
        10'b0100000010: data <= 11'h002; 
        10'b0100000011: data <= 11'h003; 
        10'b0100000100: data <= 11'h003; 
        10'b0100000101: data <= 11'h002; 
        10'b0100000110: data <= 11'h005; 
        10'b0100000111: data <= 11'h006; 
        10'b0100001000: data <= 11'h007; 
        10'b0100001001: data <= 11'h006; 
        10'b0100001010: data <= 11'h009; 
        10'b0100001011: data <= 11'h00b; 
        10'b0100001100: data <= 11'h00a; 
        10'b0100001101: data <= 11'h00b; 
        10'b0100001110: data <= 11'h007; 
        10'b0100001111: data <= 11'h007; 
        10'b0100010000: data <= 11'h006; 
        10'b0100010001: data <= 11'h005; 
        10'b0100010010: data <= 11'h002; 
        10'b0100010011: data <= 11'h7ff; 
        10'b0100010100: data <= 11'h7fe; 
        10'b0100010101: data <= 11'h7ff; 
        10'b0100010110: data <= 11'h001; 
        10'b0100010111: data <= 11'h000; 
        10'b0100011000: data <= 11'h000; 
        10'b0100011001: data <= 11'h001; 
        10'b0100011010: data <= 11'h001; 
        10'b0100011011: data <= 11'h004; 
        10'b0100011100: data <= 11'h005; 
        10'b0100011101: data <= 11'h004; 
        10'b0100011110: data <= 11'h001; 
        10'b0100011111: data <= 11'h001; 
        10'b0100100000: data <= 11'h7fe; 
        10'b0100100001: data <= 11'h000; 
        10'b0100100010: data <= 11'h003; 
        10'b0100100011: data <= 11'h005; 
        10'b0100100100: data <= 11'h004; 
        10'b0100100101: data <= 11'h008; 
        10'b0100100110: data <= 11'h00b; 
        10'b0100100111: data <= 11'h00d; 
        10'b0100101000: data <= 11'h00f; 
        10'b0100101001: data <= 11'h00b; 
        10'b0100101010: data <= 11'h009; 
        10'b0100101011: data <= 11'h009; 
        10'b0100101100: data <= 11'h008; 
        10'b0100101101: data <= 11'h007; 
        10'b0100101110: data <= 11'h003; 
        10'b0100101111: data <= 11'h7ff; 
        10'b0100110000: data <= 11'h7fe; 
        10'b0100110001: data <= 11'h7ff; 
        10'b0100110010: data <= 11'h000; 
        10'b0100110011: data <= 11'h000; 
        10'b0100110100: data <= 11'h001; 
        10'b0100110101: data <= 11'h001; 
        10'b0100110110: data <= 11'h001; 
        10'b0100110111: data <= 11'h004; 
        10'b0100111000: data <= 11'h005; 
        10'b0100111001: data <= 11'h003; 
        10'b0100111010: data <= 11'h001; 
        10'b0100111011: data <= 11'h001; 
        10'b0100111100: data <= 11'h000; 
        10'b0100111101: data <= 11'h003; 
        10'b0100111110: data <= 11'h002; 
        10'b0100111111: data <= 11'h002; 
        10'b0101000000: data <= 11'h003; 
        10'b0101000001: data <= 11'h003; 
        10'b0101000010: data <= 11'h003; 
        10'b0101000011: data <= 11'h00a; 
        10'b0101000100: data <= 11'h00d; 
        10'b0101000101: data <= 11'h009; 
        10'b0101000110: data <= 11'h009; 
        10'b0101000111: data <= 11'h007; 
        10'b0101001000: data <= 11'h007; 
        10'b0101001001: data <= 11'h004; 
        10'b0101001010: data <= 11'h003; 
        10'b0101001011: data <= 11'h7ff; 
        10'b0101001100: data <= 11'h7fd; 
        10'b0101001101: data <= 11'h000; 
        10'b0101001110: data <= 11'h000; 
        10'b0101001111: data <= 11'h001; 
        10'b0101010000: data <= 11'h001; 
        10'b0101010001: data <= 11'h000; 
        10'b0101010010: data <= 11'h001; 
        10'b0101010011: data <= 11'h003; 
        10'b0101010100: data <= 11'h003; 
        10'b0101010101: data <= 11'h001; 
        10'b0101010110: data <= 11'h001; 
        10'b0101010111: data <= 11'h003; 
        10'b0101011000: data <= 11'h002; 
        10'b0101011001: data <= 11'h000; 
        10'b0101011010: data <= 11'h7fe; 
        10'b0101011011: data <= 11'h7fa; 
        10'b0101011100: data <= 11'h7f2; 
        10'b0101011101: data <= 11'h7eb; 
        10'b0101011110: data <= 11'h7f0; 
        10'b0101011111: data <= 11'h000; 
        10'b0101100000: data <= 11'h009; 
        10'b0101100001: data <= 11'h008; 
        10'b0101100010: data <= 11'h003; 
        10'b0101100011: data <= 11'h001; 
        10'b0101100100: data <= 11'h000; 
        10'b0101100101: data <= 11'h7ff; 
        10'b0101100110: data <= 11'h7ff; 
        10'b0101100111: data <= 11'h7fe; 
        10'b0101101000: data <= 11'h7ff; 
        10'b0101101001: data <= 11'h001; 
        10'b0101101010: data <= 11'h001; 
        10'b0101101011: data <= 11'h000; 
        10'b0101101100: data <= 11'h001; 
        10'b0101101101: data <= 11'h001; 
        10'b0101101110: data <= 11'h001; 
        10'b0101101111: data <= 11'h002; 
        10'b0101110000: data <= 11'h001; 
        10'b0101110001: data <= 11'h000; 
        10'b0101110010: data <= 11'h7ff; 
        10'b0101110011: data <= 11'h001; 
        10'b0101110100: data <= 11'h000; 
        10'b0101110101: data <= 11'h7fe; 
        10'b0101110110: data <= 11'h7f9; 
        10'b0101110111: data <= 11'h7f2; 
        10'b0101111000: data <= 11'h7e7; 
        10'b0101111001: data <= 11'h7e4; 
        10'b0101111010: data <= 11'h7f1; 
        10'b0101111011: data <= 11'h7fe; 
        10'b0101111100: data <= 11'h005; 
        10'b0101111101: data <= 11'h003; 
        10'b0101111110: data <= 11'h001; 
        10'b0101111111: data <= 11'h001; 
        10'b0110000000: data <= 11'h7fd; 
        10'b0110000001: data <= 11'h7fd; 
        10'b0110000010: data <= 11'h7ff; 
        10'b0110000011: data <= 11'h000; 
        10'b0110000100: data <= 11'h7ff; 
        10'b0110000101: data <= 11'h7ff; 
        10'b0110000110: data <= 11'h001; 
        10'b0110000111: data <= 11'h7ff; 
        10'b0110001000: data <= 11'h000; 
        10'b0110001001: data <= 11'h001; 
        10'b0110001010: data <= 11'h002; 
        10'b0110001011: data <= 11'h003; 
        10'b0110001100: data <= 11'h002; 
        10'b0110001101: data <= 11'h002; 
        10'b0110001110: data <= 11'h7ff; 
        10'b0110001111: data <= 11'h7ff; 
        10'b0110010000: data <= 11'h7fd; 
        10'b0110010001: data <= 11'h7f9; 
        10'b0110010010: data <= 11'h7f5; 
        10'b0110010011: data <= 11'h7ef; 
        10'b0110010100: data <= 11'h7eb; 
        10'b0110010101: data <= 11'h7ee; 
        10'b0110010110: data <= 11'h7f9; 
        10'b0110010111: data <= 11'h000; 
        10'b0110011000: data <= 11'h001; 
        10'b0110011001: data <= 11'h003; 
        10'b0110011010: data <= 11'h008; 
        10'b0110011011: data <= 11'h009; 
        10'b0110011100: data <= 11'h005; 
        10'b0110011101: data <= 11'h003; 
        10'b0110011110: data <= 11'h003; 
        10'b0110011111: data <= 11'h003; 
        10'b0110100000: data <= 11'h001; 
        10'b0110100001: data <= 11'h000; 
        10'b0110100010: data <= 11'h000; 
        10'b0110100011: data <= 11'h000; 
        10'b0110100100: data <= 11'h001; 
        10'b0110100101: data <= 11'h001; 
        10'b0110100110: data <= 11'h000; 
        10'b0110100111: data <= 11'h001; 
        10'b0110101000: data <= 11'h001; 
        10'b0110101001: data <= 11'h7fd; 
        10'b0110101010: data <= 11'h7ff; 
        10'b0110101011: data <= 11'h7fe; 
        10'b0110101100: data <= 11'h7f8; 
        10'b0110101101: data <= 11'h7f6; 
        10'b0110101110: data <= 11'h7f3; 
        10'b0110101111: data <= 11'h7f1; 
        10'b0110110000: data <= 11'h7f0; 
        10'b0110110001: data <= 11'h7f4; 
        10'b0110110010: data <= 11'h7f9; 
        10'b0110110011: data <= 11'h000; 
        10'b0110110100: data <= 11'h001; 
        10'b0110110101: data <= 11'h00b; 
        10'b0110110110: data <= 11'h00d; 
        10'b0110110111: data <= 11'h00b; 
        10'b0110111000: data <= 11'h00a; 
        10'b0110111001: data <= 11'h008; 
        10'b0110111010: data <= 11'h005; 
        10'b0110111011: data <= 11'h002; 
        10'b0110111100: data <= 11'h000; 
        10'b0110111101: data <= 11'h7ff; 
        10'b0110111110: data <= 11'h000; 
        10'b0110111111: data <= 11'h001; 
        10'b0111000000: data <= 11'h001; 
        10'b0111000001: data <= 11'h001; 
        10'b0111000010: data <= 11'h000; 
        10'b0111000011: data <= 11'h001; 
        10'b0111000100: data <= 11'h001; 
        10'b0111000101: data <= 11'h7ff; 
        10'b0111000110: data <= 11'h7fe; 
        10'b0111000111: data <= 11'h000; 
        10'b0111001000: data <= 11'h7fa; 
        10'b0111001001: data <= 11'h7f9; 
        10'b0111001010: data <= 11'h7f4; 
        10'b0111001011: data <= 11'h7f2; 
        10'b0111001100: data <= 11'h7f7; 
        10'b0111001101: data <= 11'h7fb; 
        10'b0111001110: data <= 11'h7f9; 
        10'b0111001111: data <= 11'h004; 
        10'b0111010000: data <= 11'h004; 
        10'b0111010001: data <= 11'h009; 
        10'b0111010010: data <= 11'h008; 
        10'b0111010011: data <= 11'h008; 
        10'b0111010100: data <= 11'h007; 
        10'b0111010101: data <= 11'h005; 
        10'b0111010110: data <= 11'h001; 
        10'b0111010111: data <= 11'h7fe; 
        10'b0111011000: data <= 11'h7ff; 
        10'b0111011001: data <= 11'h7ff; 
        10'b0111011010: data <= 11'h001; 
        10'b0111011011: data <= 11'h001; 
        10'b0111011100: data <= 11'h000; 
        10'b0111011101: data <= 11'h000; 
        10'b0111011110: data <= 11'h001; 
        10'b0111011111: data <= 11'h000; 
        10'b0111100000: data <= 11'h000; 
        10'b0111100001: data <= 11'h7ff; 
        10'b0111100010: data <= 11'h7fc; 
        10'b0111100011: data <= 11'h7fa; 
        10'b0111100100: data <= 11'h7f9; 
        10'b0111100101: data <= 11'h7fa; 
        10'b0111100110: data <= 11'h7f8; 
        10'b0111100111: data <= 11'h7fa; 
        10'b0111101000: data <= 11'h7fe; 
        10'b0111101001: data <= 11'h001; 
        10'b0111101010: data <= 11'h001; 
        10'b0111101011: data <= 11'h001; 
        10'b0111101100: data <= 11'h7ff; 
        10'b0111101101: data <= 11'h002; 
        10'b0111101110: data <= 11'h002; 
        10'b0111101111: data <= 11'h001; 
        10'b0111110000: data <= 11'h001; 
        10'b0111110001: data <= 11'h7ff; 
        10'b0111110010: data <= 11'h7fd; 
        10'b0111110011: data <= 11'h7ff; 
        10'b0111110100: data <= 11'h7ff; 
        10'b0111110101: data <= 11'h7ff; 
        10'b0111110110: data <= 11'h000; 
        10'b0111110111: data <= 11'h000; 
        10'b0111111000: data <= 11'h000; 
        10'b0111111001: data <= 11'h000; 
        10'b0111111010: data <= 11'h001; 
        10'b0111111011: data <= 11'h000; 
        10'b0111111100: data <= 11'h7fe; 
        10'b0111111101: data <= 11'h7fc; 
        10'b0111111110: data <= 11'h7f9; 
        10'b0111111111: data <= 11'h7f7; 
        10'b1000000000: data <= 11'h7f8; 
        10'b1000000001: data <= 11'h7f9; 
        10'b1000000010: data <= 11'h7f7; 
        10'b1000000011: data <= 11'h7fd; 
        10'b1000000100: data <= 11'h7ff; 
        10'b1000000101: data <= 11'h000; 
        10'b1000000110: data <= 11'h003; 
        10'b1000000111: data <= 11'h7fd; 
        10'b1000001000: data <= 11'h7fd; 
        10'b1000001001: data <= 11'h7fe; 
        10'b1000001010: data <= 11'h7fc; 
        10'b1000001011: data <= 11'h7fd; 
        10'b1000001100: data <= 11'h7fc; 
        10'b1000001101: data <= 11'h7f9; 
        10'b1000001110: data <= 11'h7fb; 
        10'b1000001111: data <= 11'h7fd; 
        10'b1000010000: data <= 11'h7fd; 
        10'b1000010001: data <= 11'h000; 
        10'b1000010010: data <= 11'h000; 
        10'b1000010011: data <= 11'h000; 
        10'b1000010100: data <= 11'h001; 
        10'b1000010101: data <= 11'h001; 
        10'b1000010110: data <= 11'h001; 
        10'b1000010111: data <= 11'h001; 
        10'b1000011000: data <= 11'h7ff; 
        10'b1000011001: data <= 11'h7fb; 
        10'b1000011010: data <= 11'h7f7; 
        10'b1000011011: data <= 11'h7f7; 
        10'b1000011100: data <= 11'h7f7; 
        10'b1000011101: data <= 11'h7f6; 
        10'b1000011110: data <= 11'h7fa; 
        10'b1000011111: data <= 11'h7fb; 
        10'b1000100000: data <= 11'h7fd; 
        10'b1000100001: data <= 11'h001; 
        10'b1000100010: data <= 11'h004; 
        10'b1000100011: data <= 11'h7fc; 
        10'b1000100100: data <= 11'h7fc; 
        10'b1000100101: data <= 11'h7fb; 
        10'b1000100110: data <= 11'h7f8; 
        10'b1000100111: data <= 11'h7f9; 
        10'b1000101000: data <= 11'h7f7; 
        10'b1000101001: data <= 11'h7f8; 
        10'b1000101010: data <= 11'h7fa; 
        10'b1000101011: data <= 11'h7fc; 
        10'b1000101100: data <= 11'h7fe; 
        10'b1000101101: data <= 11'h7ff; 
        10'b1000101110: data <= 11'h001; 
        10'b1000101111: data <= 11'h7ff; 
        10'b1000110000: data <= 11'h7ff; 
        10'b1000110001: data <= 11'h000; 
        10'b1000110010: data <= 11'h001; 
        10'b1000110011: data <= 11'h000; 
        10'b1000110100: data <= 11'h7ff; 
        10'b1000110101: data <= 11'h7fc; 
        10'b1000110110: data <= 11'h7f7; 
        10'b1000110111: data <= 11'h7f7; 
        10'b1000111000: data <= 11'h7f7; 
        10'b1000111001: data <= 11'h7f8; 
        10'b1000111010: data <= 11'h7fa; 
        10'b1000111011: data <= 11'h7fa; 
        10'b1000111100: data <= 11'h000; 
        10'b1000111101: data <= 11'h001; 
        10'b1000111110: data <= 11'h002; 
        10'b1000111111: data <= 11'h7fb; 
        10'b1001000000: data <= 11'h7f9; 
        10'b1001000001: data <= 11'h7f7; 
        10'b1001000010: data <= 11'h7f4; 
        10'b1001000011: data <= 11'h7f8; 
        10'b1001000100: data <= 11'h7f6; 
        10'b1001000101: data <= 11'h7f8; 
        10'b1001000110: data <= 11'h7fa; 
        10'b1001000111: data <= 11'h7fe; 
        10'b1001001000: data <= 11'h7fe; 
        10'b1001001001: data <= 11'h001; 
        10'b1001001010: data <= 11'h001; 
        10'b1001001011: data <= 11'h001; 
        10'b1001001100: data <= 11'h001; 
        10'b1001001101: data <= 11'h001; 
        10'b1001001110: data <= 11'h000; 
        10'b1001001111: data <= 11'h7fe; 
        10'b1001010000: data <= 11'h7ff; 
        10'b1001010001: data <= 11'h7fc; 
        10'b1001010010: data <= 11'h7fc; 
        10'b1001010011: data <= 11'h7fa; 
        10'b1001010100: data <= 11'h7fa; 
        10'b1001010101: data <= 11'h7fd; 
        10'b1001010110: data <= 11'h7fb; 
        10'b1001010111: data <= 11'h7fc; 
        10'b1001011000: data <= 11'h7fe; 
        10'b1001011001: data <= 11'h000; 
        10'b1001011010: data <= 11'h7ff; 
        10'b1001011011: data <= 11'h7fc; 
        10'b1001011100: data <= 11'h7fc; 
        10'b1001011101: data <= 11'h7f7; 
        10'b1001011110: data <= 11'h7f8; 
        10'b1001011111: data <= 11'h7f8; 
        10'b1001100000: data <= 11'h7f7; 
        10'b1001100001: data <= 11'h7f8; 
        10'b1001100010: data <= 11'h7fc; 
        10'b1001100011: data <= 11'h7fd; 
        10'b1001100100: data <= 11'h000; 
        10'b1001100101: data <= 11'h001; 
        10'b1001100110: data <= 11'h001; 
        10'b1001100111: data <= 11'h000; 
        10'b1001101000: data <= 11'h000; 
        10'b1001101001: data <= 11'h000; 
        10'b1001101010: data <= 11'h000; 
        10'b1001101011: data <= 11'h7ff; 
        10'b1001101100: data <= 11'h000; 
        10'b1001101101: data <= 11'h001; 
        10'b1001101110: data <= 11'h7ff; 
        10'b1001101111: data <= 11'h001; 
        10'b1001110000: data <= 11'h001; 
        10'b1001110001: data <= 11'h7fe; 
        10'b1001110010: data <= 11'h7fd; 
        10'b1001110011: data <= 11'h7fa; 
        10'b1001110100: data <= 11'h7fb; 
        10'b1001110101: data <= 11'h7fe; 
        10'b1001110110: data <= 11'h001; 
        10'b1001110111: data <= 11'h001; 
        10'b1001111000: data <= 11'h7fd; 
        10'b1001111001: data <= 11'h7fc; 
        10'b1001111010: data <= 11'h7f9; 
        10'b1001111011: data <= 11'h7f9; 
        10'b1001111100: data <= 11'h7f8; 
        10'b1001111101: data <= 11'h7f9; 
        10'b1001111110: data <= 11'h7fd; 
        10'b1001111111: data <= 11'h7ff; 
        10'b1010000000: data <= 11'h001; 
        10'b1010000001: data <= 11'h7ff; 
        10'b1010000010: data <= 11'h000; 
        10'b1010000011: data <= 11'h000; 
        10'b1010000100: data <= 11'h001; 
        10'b1010000101: data <= 11'h001; 
        10'b1010000110: data <= 11'h7ff; 
        10'b1010000111: data <= 11'h7ff; 
        10'b1010001000: data <= 11'h001; 
        10'b1010001001: data <= 11'h002; 
        10'b1010001010: data <= 11'h004; 
        10'b1010001011: data <= 11'h005; 
        10'b1010001100: data <= 11'h003; 
        10'b1010001101: data <= 11'h001; 
        10'b1010001110: data <= 11'h7fe; 
        10'b1010001111: data <= 11'h7fc; 
        10'b1010010000: data <= 11'h7fd; 
        10'b1010010001: data <= 11'h000; 
        10'b1010010010: data <= 11'h002; 
        10'b1010010011: data <= 11'h002; 
        10'b1010010100: data <= 11'h7ff; 
        10'b1010010101: data <= 11'h7ff; 
        10'b1010010110: data <= 11'h7fc; 
        10'b1010010111: data <= 11'h7fa; 
        10'b1010011000: data <= 11'h7fa; 
        10'b1010011001: data <= 11'h7fb; 
        10'b1010011010: data <= 11'h7fc; 
        10'b1010011011: data <= 11'h7fd; 
        10'b1010011100: data <= 11'h7ff; 
        10'b1010011101: data <= 11'h000; 
        10'b1010011110: data <= 11'h000; 
        10'b1010011111: data <= 11'h000; 
        10'b1010100000: data <= 11'h000; 
        10'b1010100001: data <= 11'h000; 
        10'b1010100010: data <= 11'h000; 
        10'b1010100011: data <= 11'h001; 
        10'b1010100100: data <= 11'h002; 
        10'b1010100101: data <= 11'h004; 
        10'b1010100110: data <= 11'h007; 
        10'b1010100111: data <= 11'h008; 
        10'b1010101000: data <= 11'h007; 
        10'b1010101001: data <= 11'h003; 
        10'b1010101010: data <= 11'h007; 
        10'b1010101011: data <= 11'h004; 
        10'b1010101100: data <= 11'h004; 
        10'b1010101101: data <= 11'h005; 
        10'b1010101110: data <= 11'h003; 
        10'b1010101111: data <= 11'h005; 
        10'b1010110000: data <= 11'h003; 
        10'b1010110001: data <= 11'h002; 
        10'b1010110010: data <= 11'h000; 
        10'b1010110011: data <= 11'h7fe; 
        10'b1010110100: data <= 11'h7fe; 
        10'b1010110101: data <= 11'h7fd; 
        10'b1010110110: data <= 11'h7fd; 
        10'b1010110111: data <= 11'h7fd; 
        10'b1010111000: data <= 11'h000; 
        10'b1010111001: data <= 11'h000; 
        10'b1010111010: data <= 11'h7ff; 
        10'b1010111011: data <= 11'h001; 
        10'b1010111100: data <= 11'h7ff; 
        10'b1010111101: data <= 11'h001; 
        10'b1010111110: data <= 11'h001; 
        10'b1010111111: data <= 11'h001; 
        10'b1011000000: data <= 11'h001; 
        10'b1011000001: data <= 11'h002; 
        10'b1011000010: data <= 11'h003; 
        10'b1011000011: data <= 11'h005; 
        10'b1011000100: data <= 11'h008; 
        10'b1011000101: data <= 11'h008; 
        10'b1011000110: data <= 11'h009; 
        10'b1011000111: data <= 11'h009; 
        10'b1011001000: data <= 11'h008; 
        10'b1011001001: data <= 11'h006; 
        10'b1011001010: data <= 11'h006; 
        10'b1011001011: data <= 11'h007; 
        10'b1011001100: data <= 11'h005; 
        10'b1011001101: data <= 11'h005; 
        10'b1011001110: data <= 11'h004; 
        10'b1011001111: data <= 11'h001; 
        10'b1011010000: data <= 11'h7fe; 
        10'b1011010001: data <= 11'h000; 
        10'b1011010010: data <= 11'h7ff; 
        10'b1011010011: data <= 11'h7ff; 
        10'b1011010100: data <= 11'h000; 
        10'b1011010101: data <= 11'h000; 
        10'b1011010110: data <= 11'h002; 
        10'b1011010111: data <= 11'h001; 
        10'b1011011000: data <= 11'h7ff; 
        10'b1011011001: data <= 11'h000; 
        10'b1011011010: data <= 11'h001; 
        10'b1011011011: data <= 11'h000; 
        10'b1011011100: data <= 11'h000; 
        10'b1011011101: data <= 11'h001; 
        10'b1011011110: data <= 11'h000; 
        10'b1011011111: data <= 11'h001; 
        10'b1011100000: data <= 11'h001; 
        10'b1011100001: data <= 11'h000; 
        10'b1011100010: data <= 11'h002; 
        10'b1011100011: data <= 11'h003; 
        10'b1011100100: data <= 11'h001; 
        10'b1011100101: data <= 11'h002; 
        10'b1011100110: data <= 11'h005; 
        10'b1011100111: data <= 11'h006; 
        10'b1011101000: data <= 11'h005; 
        10'b1011101001: data <= 11'h006; 
        10'b1011101010: data <= 11'h003; 
        10'b1011101011: data <= 11'h002; 
        10'b1011101100: data <= 11'h000; 
        10'b1011101101: data <= 11'h001; 
        10'b1011101110: data <= 11'h000; 
        10'b1011101111: data <= 11'h000; 
        10'b1011110000: data <= 11'h000; 
        10'b1011110001: data <= 11'h000; 
        10'b1011110010: data <= 11'h000; 
        10'b1011110011: data <= 11'h000; 
        10'b1011110100: data <= 11'h7ff; 
        10'b1011110101: data <= 11'h001; 
        10'b1011110110: data <= 11'h000; 
        10'b1011110111: data <= 11'h001; 
        10'b1011111000: data <= 11'h001; 
        10'b1011111001: data <= 11'h001; 
        10'b1011111010: data <= 11'h000; 
        10'b1011111011: data <= 11'h000; 
        10'b1011111100: data <= 11'h002; 
        10'b1011111101: data <= 11'h001; 
        10'b1011111110: data <= 11'h000; 
        10'b1011111111: data <= 11'h001; 
        10'b1100000000: data <= 11'h000; 
        10'b1100000001: data <= 11'h002; 
        10'b1100000010: data <= 11'h001; 
        10'b1100000011: data <= 11'h001; 
        10'b1100000100: data <= 11'h003; 
        10'b1100000101: data <= 11'h001; 
        10'b1100000110: data <= 11'h001; 
        10'b1100000111: data <= 11'h002; 
        10'b1100001000: data <= 11'h000; 
        10'b1100001001: data <= 11'h000; 
        10'b1100001010: data <= 11'h001; 
        10'b1100001011: data <= 11'h001; 
        10'b1100001100: data <= 11'h000; 
        10'b1100001101: data <= 11'h000; 
        10'b1100001110: data <= 11'h7ff; 
        10'b1100001111: data <= 11'h001; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 6) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 12'h000; 
        10'b0000000001: data <= 12'h000; 
        10'b0000000010: data <= 12'h002; 
        10'b0000000011: data <= 12'h001; 
        10'b0000000100: data <= 12'h003; 
        10'b0000000101: data <= 12'hfff; 
        10'b0000000110: data <= 12'hfff; 
        10'b0000000111: data <= 12'h001; 
        10'b0000001000: data <= 12'h002; 
        10'b0000001001: data <= 12'h002; 
        10'b0000001010: data <= 12'hfff; 
        10'b0000001011: data <= 12'h001; 
        10'b0000001100: data <= 12'h001; 
        10'b0000001101: data <= 12'h000; 
        10'b0000001110: data <= 12'h002; 
        10'b0000001111: data <= 12'h001; 
        10'b0000010000: data <= 12'h000; 
        10'b0000010001: data <= 12'h000; 
        10'b0000010010: data <= 12'h000; 
        10'b0000010011: data <= 12'h001; 
        10'b0000010100: data <= 12'h002; 
        10'b0000010101: data <= 12'h003; 
        10'b0000010110: data <= 12'hfff; 
        10'b0000010111: data <= 12'h002; 
        10'b0000011000: data <= 12'h000; 
        10'b0000011001: data <= 12'h002; 
        10'b0000011010: data <= 12'h000; 
        10'b0000011011: data <= 12'h000; 
        10'b0000011100: data <= 12'h003; 
        10'b0000011101: data <= 12'hfff; 
        10'b0000011110: data <= 12'h001; 
        10'b0000011111: data <= 12'h003; 
        10'b0000100000: data <= 12'h001; 
        10'b0000100001: data <= 12'h000; 
        10'b0000100010: data <= 12'h003; 
        10'b0000100011: data <= 12'h001; 
        10'b0000100100: data <= 12'h000; 
        10'b0000100101: data <= 12'h000; 
        10'b0000100110: data <= 12'h000; 
        10'b0000100111: data <= 12'hfff; 
        10'b0000101000: data <= 12'h002; 
        10'b0000101001: data <= 12'h000; 
        10'b0000101010: data <= 12'h003; 
        10'b0000101011: data <= 12'hfff; 
        10'b0000101100: data <= 12'h001; 
        10'b0000101101: data <= 12'h002; 
        10'b0000101110: data <= 12'h002; 
        10'b0000101111: data <= 12'h002; 
        10'b0000110000: data <= 12'h000; 
        10'b0000110001: data <= 12'h002; 
        10'b0000110010: data <= 12'h000; 
        10'b0000110011: data <= 12'h003; 
        10'b0000110100: data <= 12'h002; 
        10'b0000110101: data <= 12'hfff; 
        10'b0000110110: data <= 12'hfff; 
        10'b0000110111: data <= 12'h001; 
        10'b0000111000: data <= 12'h003; 
        10'b0000111001: data <= 12'h003; 
        10'b0000111010: data <= 12'h002; 
        10'b0000111011: data <= 12'h000; 
        10'b0000111100: data <= 12'h002; 
        10'b0000111101: data <= 12'hfff; 
        10'b0000111110: data <= 12'hfff; 
        10'b0000111111: data <= 12'h002; 
        10'b0001000000: data <= 12'h002; 
        10'b0001000001: data <= 12'hfff; 
        10'b0001000010: data <= 12'h000; 
        10'b0001000011: data <= 12'h001; 
        10'b0001000100: data <= 12'h000; 
        10'b0001000101: data <= 12'hfff; 
        10'b0001000110: data <= 12'h001; 
        10'b0001000111: data <= 12'h002; 
        10'b0001001000: data <= 12'h002; 
        10'b0001001001: data <= 12'h000; 
        10'b0001001010: data <= 12'h001; 
        10'b0001001011: data <= 12'h003; 
        10'b0001001100: data <= 12'h002; 
        10'b0001001101: data <= 12'h003; 
        10'b0001001110: data <= 12'hfff; 
        10'b0001001111: data <= 12'h002; 
        10'b0001010000: data <= 12'h001; 
        10'b0001010001: data <= 12'h002; 
        10'b0001010010: data <= 12'h002; 
        10'b0001010011: data <= 12'h002; 
        10'b0001010100: data <= 12'h000; 
        10'b0001010101: data <= 12'h000; 
        10'b0001010110: data <= 12'h002; 
        10'b0001010111: data <= 12'h000; 
        10'b0001011000: data <= 12'h000; 
        10'b0001011001: data <= 12'h000; 
        10'b0001011010: data <= 12'hfff; 
        10'b0001011011: data <= 12'h002; 
        10'b0001011100: data <= 12'h000; 
        10'b0001011101: data <= 12'h002; 
        10'b0001011110: data <= 12'hfff; 
        10'b0001011111: data <= 12'h000; 
        10'b0001100000: data <= 12'h001; 
        10'b0001100001: data <= 12'hffe; 
        10'b0001100010: data <= 12'h001; 
        10'b0001100011: data <= 12'hfff; 
        10'b0001100100: data <= 12'hffd; 
        10'b0001100101: data <= 12'hffe; 
        10'b0001100110: data <= 12'hffe; 
        10'b0001100111: data <= 12'hfff; 
        10'b0001101000: data <= 12'h000; 
        10'b0001101001: data <= 12'hfff; 
        10'b0001101010: data <= 12'h001; 
        10'b0001101011: data <= 12'h000; 
        10'b0001101100: data <= 12'h001; 
        10'b0001101101: data <= 12'h003; 
        10'b0001101110: data <= 12'hfff; 
        10'b0001101111: data <= 12'h001; 
        10'b0001110000: data <= 12'h003; 
        10'b0001110001: data <= 12'hfff; 
        10'b0001110010: data <= 12'h002; 
        10'b0001110011: data <= 12'hfff; 
        10'b0001110100: data <= 12'h001; 
        10'b0001110101: data <= 12'hfff; 
        10'b0001110110: data <= 12'h000; 
        10'b0001110111: data <= 12'hfff; 
        10'b0001111000: data <= 12'h001; 
        10'b0001111001: data <= 12'h000; 
        10'b0001111010: data <= 12'hffd; 
        10'b0001111011: data <= 12'hffa; 
        10'b0001111100: data <= 12'hffa; 
        10'b0001111101: data <= 12'hffa; 
        10'b0001111110: data <= 12'hff9; 
        10'b0001111111: data <= 12'hff5; 
        10'b0010000000: data <= 12'hffa; 
        10'b0010000001: data <= 12'hffb; 
        10'b0010000010: data <= 12'hffc; 
        10'b0010000011: data <= 12'hfff; 
        10'b0010000100: data <= 12'hffd; 
        10'b0010000101: data <= 12'h001; 
        10'b0010000110: data <= 12'h000; 
        10'b0010000111: data <= 12'hffe; 
        10'b0010001000: data <= 12'h003; 
        10'b0010001001: data <= 12'h000; 
        10'b0010001010: data <= 12'h003; 
        10'b0010001011: data <= 12'h003; 
        10'b0010001100: data <= 12'h003; 
        10'b0010001101: data <= 12'h000; 
        10'b0010001110: data <= 12'h002; 
        10'b0010001111: data <= 12'hfff; 
        10'b0010010000: data <= 12'hffe; 
        10'b0010010001: data <= 12'h000; 
        10'b0010010010: data <= 12'hfff; 
        10'b0010010011: data <= 12'hfff; 
        10'b0010010100: data <= 12'hffe; 
        10'b0010010101: data <= 12'hffc; 
        10'b0010010110: data <= 12'hff6; 
        10'b0010010111: data <= 12'hff4; 
        10'b0010011000: data <= 12'hff1; 
        10'b0010011001: data <= 12'hfee; 
        10'b0010011010: data <= 12'hfea; 
        10'b0010011011: data <= 12'hfea; 
        10'b0010011100: data <= 12'hfe9; 
        10'b0010011101: data <= 12'hfec; 
        10'b0010011110: data <= 12'hfef; 
        10'b0010011111: data <= 12'hff3; 
        10'b0010100000: data <= 12'hff7; 
        10'b0010100001: data <= 12'hffd; 
        10'b0010100010: data <= 12'hffb; 
        10'b0010100011: data <= 12'hfff; 
        10'b0010100100: data <= 12'h002; 
        10'b0010100101: data <= 12'h002; 
        10'b0010100110: data <= 12'h000; 
        10'b0010100111: data <= 12'h000; 
        10'b0010101000: data <= 12'h002; 
        10'b0010101001: data <= 12'h003; 
        10'b0010101010: data <= 12'h000; 
        10'b0010101011: data <= 12'h000; 
        10'b0010101100: data <= 12'h003; 
        10'b0010101101: data <= 12'h004; 
        10'b0010101110: data <= 12'h004; 
        10'b0010101111: data <= 12'h007; 
        10'b0010110000: data <= 12'h00a; 
        10'b0010110001: data <= 12'h008; 
        10'b0010110010: data <= 12'h008; 
        10'b0010110011: data <= 12'h001; 
        10'b0010110100: data <= 12'hff9; 
        10'b0010110101: data <= 12'hff2; 
        10'b0010110110: data <= 12'hff2; 
        10'b0010110111: data <= 12'hff8; 
        10'b0010111000: data <= 12'hffb; 
        10'b0010111001: data <= 12'hffb; 
        10'b0010111010: data <= 12'hff9; 
        10'b0010111011: data <= 12'hff8; 
        10'b0010111100: data <= 12'hff5; 
        10'b0010111101: data <= 12'hffc; 
        10'b0010111110: data <= 12'hff8; 
        10'b0010111111: data <= 12'hffa; 
        10'b0011000000: data <= 12'hffc; 
        10'b0011000001: data <= 12'hfff; 
        10'b0011000010: data <= 12'hfff; 
        10'b0011000011: data <= 12'h000; 
        10'b0011000100: data <= 12'h002; 
        10'b0011000101: data <= 12'h003; 
        10'b0011000110: data <= 12'h002; 
        10'b0011000111: data <= 12'h006; 
        10'b0011001000: data <= 12'h007; 
        10'b0011001001: data <= 12'h006; 
        10'b0011001010: data <= 12'h009; 
        10'b0011001011: data <= 12'h00e; 
        10'b0011001100: data <= 12'h013; 
        10'b0011001101: data <= 12'h00f; 
        10'b0011001110: data <= 12'h00a; 
        10'b0011001111: data <= 12'h00b; 
        10'b0011010000: data <= 12'h00c; 
        10'b0011010001: data <= 12'h002; 
        10'b0011010010: data <= 12'h002; 
        10'b0011010011: data <= 12'h004; 
        10'b0011010100: data <= 12'h00d; 
        10'b0011010101: data <= 12'h00e; 
        10'b0011010110: data <= 12'h009; 
        10'b0011010111: data <= 12'h008; 
        10'b0011011000: data <= 12'h002; 
        10'b0011011001: data <= 12'hffe; 
        10'b0011011010: data <= 12'h001; 
        10'b0011011011: data <= 12'hffe; 
        10'b0011011100: data <= 12'hffe; 
        10'b0011011101: data <= 12'h000; 
        10'b0011011110: data <= 12'h002; 
        10'b0011011111: data <= 12'hfff; 
        10'b0011100000: data <= 12'hfff; 
        10'b0011100001: data <= 12'h003; 
        10'b0011100010: data <= 12'h001; 
        10'b0011100011: data <= 12'h005; 
        10'b0011100100: data <= 12'h00a; 
        10'b0011100101: data <= 12'h009; 
        10'b0011100110: data <= 12'h00c; 
        10'b0011100111: data <= 12'h015; 
        10'b0011101000: data <= 12'h00e; 
        10'b0011101001: data <= 12'h00a; 
        10'b0011101010: data <= 12'h00c; 
        10'b0011101011: data <= 12'h010; 
        10'b0011101100: data <= 12'h010; 
        10'b0011101101: data <= 12'h008; 
        10'b0011101110: data <= 12'h005; 
        10'b0011101111: data <= 12'h006; 
        10'b0011110000: data <= 12'h00b; 
        10'b0011110001: data <= 12'h011; 
        10'b0011110010: data <= 12'h00c; 
        10'b0011110011: data <= 12'h00a; 
        10'b0011110100: data <= 12'h008; 
        10'b0011110101: data <= 12'h000; 
        10'b0011110110: data <= 12'h005; 
        10'b0011110111: data <= 12'h004; 
        10'b0011111000: data <= 12'hffd; 
        10'b0011111001: data <= 12'hfff; 
        10'b0011111010: data <= 12'h002; 
        10'b0011111011: data <= 12'h002; 
        10'b0011111100: data <= 12'h001; 
        10'b0011111101: data <= 12'h002; 
        10'b0011111110: data <= 12'h003; 
        10'b0011111111: data <= 12'h007; 
        10'b0100000000: data <= 12'h009; 
        10'b0100000001: data <= 12'h00b; 
        10'b0100000010: data <= 12'h004; 
        10'b0100000011: data <= 12'h005; 
        10'b0100000100: data <= 12'h006; 
        10'b0100000101: data <= 12'h004; 
        10'b0100000110: data <= 12'h00a; 
        10'b0100000111: data <= 12'h00c; 
        10'b0100001000: data <= 12'h00f; 
        10'b0100001001: data <= 12'h00c; 
        10'b0100001010: data <= 12'h011; 
        10'b0100001011: data <= 12'h016; 
        10'b0100001100: data <= 12'h014; 
        10'b0100001101: data <= 12'h016; 
        10'b0100001110: data <= 12'h00e; 
        10'b0100001111: data <= 12'h00f; 
        10'b0100010000: data <= 12'h00c; 
        10'b0100010001: data <= 12'h00a; 
        10'b0100010010: data <= 12'h005; 
        10'b0100010011: data <= 12'hffe; 
        10'b0100010100: data <= 12'hffd; 
        10'b0100010101: data <= 12'hfff; 
        10'b0100010110: data <= 12'h001; 
        10'b0100010111: data <= 12'hfff; 
        10'b0100011000: data <= 12'h000; 
        10'b0100011001: data <= 12'h003; 
        10'b0100011010: data <= 12'h003; 
        10'b0100011011: data <= 12'h009; 
        10'b0100011100: data <= 12'h00a; 
        10'b0100011101: data <= 12'h008; 
        10'b0100011110: data <= 12'h001; 
        10'b0100011111: data <= 12'h002; 
        10'b0100100000: data <= 12'hffd; 
        10'b0100100001: data <= 12'h000; 
        10'b0100100010: data <= 12'h006; 
        10'b0100100011: data <= 12'h00a; 
        10'b0100100100: data <= 12'h007; 
        10'b0100100101: data <= 12'h011; 
        10'b0100100110: data <= 12'h016; 
        10'b0100100111: data <= 12'h01b; 
        10'b0100101000: data <= 12'h01f; 
        10'b0100101001: data <= 12'h017; 
        10'b0100101010: data <= 12'h012; 
        10'b0100101011: data <= 12'h013; 
        10'b0100101100: data <= 12'h010; 
        10'b0100101101: data <= 12'h00e; 
        10'b0100101110: data <= 12'h006; 
        10'b0100101111: data <= 12'hffe; 
        10'b0100110000: data <= 12'hffc; 
        10'b0100110001: data <= 12'hffe; 
        10'b0100110010: data <= 12'h000; 
        10'b0100110011: data <= 12'hfff; 
        10'b0100110100: data <= 12'h002; 
        10'b0100110101: data <= 12'h002; 
        10'b0100110110: data <= 12'h003; 
        10'b0100110111: data <= 12'h009; 
        10'b0100111000: data <= 12'h00b; 
        10'b0100111001: data <= 12'h005; 
        10'b0100111010: data <= 12'h002; 
        10'b0100111011: data <= 12'h002; 
        10'b0100111100: data <= 12'h000; 
        10'b0100111101: data <= 12'h006; 
        10'b0100111110: data <= 12'h003; 
        10'b0100111111: data <= 12'h004; 
        10'b0101000000: data <= 12'h007; 
        10'b0101000001: data <= 12'h007; 
        10'b0101000010: data <= 12'h007; 
        10'b0101000011: data <= 12'h015; 
        10'b0101000100: data <= 12'h01b; 
        10'b0101000101: data <= 12'h012; 
        10'b0101000110: data <= 12'h012; 
        10'b0101000111: data <= 12'h00e; 
        10'b0101001000: data <= 12'h00d; 
        10'b0101001001: data <= 12'h008; 
        10'b0101001010: data <= 12'h006; 
        10'b0101001011: data <= 12'hffe; 
        10'b0101001100: data <= 12'hffa; 
        10'b0101001101: data <= 12'h000; 
        10'b0101001110: data <= 12'h001; 
        10'b0101001111: data <= 12'h003; 
        10'b0101010000: data <= 12'h002; 
        10'b0101010001: data <= 12'h000; 
        10'b0101010010: data <= 12'h001; 
        10'b0101010011: data <= 12'h005; 
        10'b0101010100: data <= 12'h006; 
        10'b0101010101: data <= 12'h001; 
        10'b0101010110: data <= 12'h001; 
        10'b0101010111: data <= 12'h006; 
        10'b0101011000: data <= 12'h004; 
        10'b0101011001: data <= 12'h000; 
        10'b0101011010: data <= 12'hffb; 
        10'b0101011011: data <= 12'hff3; 
        10'b0101011100: data <= 12'hfe5; 
        10'b0101011101: data <= 12'hfd6; 
        10'b0101011110: data <= 12'hfe1; 
        10'b0101011111: data <= 12'h001; 
        10'b0101100000: data <= 12'h012; 
        10'b0101100001: data <= 12'h010; 
        10'b0101100010: data <= 12'h006; 
        10'b0101100011: data <= 12'h002; 
        10'b0101100100: data <= 12'h000; 
        10'b0101100101: data <= 12'hffe; 
        10'b0101100110: data <= 12'hffe; 
        10'b0101100111: data <= 12'hffc; 
        10'b0101101000: data <= 12'hffd; 
        10'b0101101001: data <= 12'h003; 
        10'b0101101010: data <= 12'h002; 
        10'b0101101011: data <= 12'h000; 
        10'b0101101100: data <= 12'h002; 
        10'b0101101101: data <= 12'h001; 
        10'b0101101110: data <= 12'h002; 
        10'b0101101111: data <= 12'h005; 
        10'b0101110000: data <= 12'h002; 
        10'b0101110001: data <= 12'h001; 
        10'b0101110010: data <= 12'hffe; 
        10'b0101110011: data <= 12'h001; 
        10'b0101110100: data <= 12'hfff; 
        10'b0101110101: data <= 12'hffc; 
        10'b0101110110: data <= 12'hff3; 
        10'b0101110111: data <= 12'hfe4; 
        10'b0101111000: data <= 12'hfce; 
        10'b0101111001: data <= 12'hfc9; 
        10'b0101111010: data <= 12'hfe2; 
        10'b0101111011: data <= 12'hffc; 
        10'b0101111100: data <= 12'h009; 
        10'b0101111101: data <= 12'h006; 
        10'b0101111110: data <= 12'h001; 
        10'b0101111111: data <= 12'h003; 
        10'b0110000000: data <= 12'hffb; 
        10'b0110000001: data <= 12'hff9; 
        10'b0110000010: data <= 12'hffe; 
        10'b0110000011: data <= 12'h001; 
        10'b0110000100: data <= 12'hfff; 
        10'b0110000101: data <= 12'hfff; 
        10'b0110000110: data <= 12'h001; 
        10'b0110000111: data <= 12'hfff; 
        10'b0110001000: data <= 12'hfff; 
        10'b0110001001: data <= 12'h001; 
        10'b0110001010: data <= 12'h004; 
        10'b0110001011: data <= 12'h006; 
        10'b0110001100: data <= 12'h004; 
        10'b0110001101: data <= 12'h004; 
        10'b0110001110: data <= 12'hfff; 
        10'b0110001111: data <= 12'hffd; 
        10'b0110010000: data <= 12'hffa; 
        10'b0110010001: data <= 12'hff1; 
        10'b0110010010: data <= 12'hfea; 
        10'b0110010011: data <= 12'hfde; 
        10'b0110010100: data <= 12'hfd5; 
        10'b0110010101: data <= 12'hfdc; 
        10'b0110010110: data <= 12'hff3; 
        10'b0110010111: data <= 12'h000; 
        10'b0110011000: data <= 12'h003; 
        10'b0110011001: data <= 12'h006; 
        10'b0110011010: data <= 12'h010; 
        10'b0110011011: data <= 12'h012; 
        10'b0110011100: data <= 12'h00b; 
        10'b0110011101: data <= 12'h007; 
        10'b0110011110: data <= 12'h007; 
        10'b0110011111: data <= 12'h006; 
        10'b0110100000: data <= 12'h002; 
        10'b0110100001: data <= 12'h001; 
        10'b0110100010: data <= 12'hfff; 
        10'b0110100011: data <= 12'hfff; 
        10'b0110100100: data <= 12'h001; 
        10'b0110100101: data <= 12'h002; 
        10'b0110100110: data <= 12'h001; 
        10'b0110100111: data <= 12'h002; 
        10'b0110101000: data <= 12'h002; 
        10'b0110101001: data <= 12'hffa; 
        10'b0110101010: data <= 12'hffd; 
        10'b0110101011: data <= 12'hffc; 
        10'b0110101100: data <= 12'hff0; 
        10'b0110101101: data <= 12'hfed; 
        10'b0110101110: data <= 12'hfe6; 
        10'b0110101111: data <= 12'hfe3; 
        10'b0110110000: data <= 12'hfe0; 
        10'b0110110001: data <= 12'hfe9; 
        10'b0110110010: data <= 12'hff2; 
        10'b0110110011: data <= 12'h000; 
        10'b0110110100: data <= 12'h001; 
        10'b0110110101: data <= 12'h016; 
        10'b0110110110: data <= 12'h01a; 
        10'b0110110111: data <= 12'h016; 
        10'b0110111000: data <= 12'h013; 
        10'b0110111001: data <= 12'h010; 
        10'b0110111010: data <= 12'h00b; 
        10'b0110111011: data <= 12'h005; 
        10'b0110111100: data <= 12'h000; 
        10'b0110111101: data <= 12'hfff; 
        10'b0110111110: data <= 12'h000; 
        10'b0110111111: data <= 12'h002; 
        10'b0111000000: data <= 12'h001; 
        10'b0111000001: data <= 12'h003; 
        10'b0111000010: data <= 12'h000; 
        10'b0111000011: data <= 12'h003; 
        10'b0111000100: data <= 12'h002; 
        10'b0111000101: data <= 12'hffd; 
        10'b0111000110: data <= 12'hffc; 
        10'b0111000111: data <= 12'hfff; 
        10'b0111001000: data <= 12'hff3; 
        10'b0111001001: data <= 12'hff2; 
        10'b0111001010: data <= 12'hfe9; 
        10'b0111001011: data <= 12'hfe4; 
        10'b0111001100: data <= 12'hfef; 
        10'b0111001101: data <= 12'hff6; 
        10'b0111001110: data <= 12'hff2; 
        10'b0111001111: data <= 12'h007; 
        10'b0111010000: data <= 12'h009; 
        10'b0111010001: data <= 12'h013; 
        10'b0111010010: data <= 12'h010; 
        10'b0111010011: data <= 12'h011; 
        10'b0111010100: data <= 12'h00d; 
        10'b0111010101: data <= 12'h00a; 
        10'b0111010110: data <= 12'h002; 
        10'b0111010111: data <= 12'hffc; 
        10'b0111011000: data <= 12'hffd; 
        10'b0111011001: data <= 12'hfff; 
        10'b0111011010: data <= 12'h002; 
        10'b0111011011: data <= 12'h003; 
        10'b0111011100: data <= 12'h000; 
        10'b0111011101: data <= 12'h000; 
        10'b0111011110: data <= 12'h002; 
        10'b0111011111: data <= 12'h000; 
        10'b0111100000: data <= 12'h001; 
        10'b0111100001: data <= 12'hffe; 
        10'b0111100010: data <= 12'hff7; 
        10'b0111100011: data <= 12'hff5; 
        10'b0111100100: data <= 12'hff2; 
        10'b0111100101: data <= 12'hff4; 
        10'b0111100110: data <= 12'hff0; 
        10'b0111100111: data <= 12'hff4; 
        10'b0111101000: data <= 12'hffc; 
        10'b0111101001: data <= 12'h003; 
        10'b0111101010: data <= 12'h002; 
        10'b0111101011: data <= 12'h003; 
        10'b0111101100: data <= 12'hffe; 
        10'b0111101101: data <= 12'h005; 
        10'b0111101110: data <= 12'h004; 
        10'b0111101111: data <= 12'h003; 
        10'b0111110000: data <= 12'h002; 
        10'b0111110001: data <= 12'hffe; 
        10'b0111110010: data <= 12'hffb; 
        10'b0111110011: data <= 12'hffe; 
        10'b0111110100: data <= 12'hffe; 
        10'b0111110101: data <= 12'hffe; 
        10'b0111110110: data <= 12'hfff; 
        10'b0111110111: data <= 12'hfff; 
        10'b0111111000: data <= 12'hfff; 
        10'b0111111001: data <= 12'h000; 
        10'b0111111010: data <= 12'h002; 
        10'b0111111011: data <= 12'h001; 
        10'b0111111100: data <= 12'hffd; 
        10'b0111111101: data <= 12'hff8; 
        10'b0111111110: data <= 12'hff2; 
        10'b0111111111: data <= 12'hfef; 
        10'b1000000000: data <= 12'hff0; 
        10'b1000000001: data <= 12'hff1; 
        10'b1000000010: data <= 12'hfed; 
        10'b1000000011: data <= 12'hff9; 
        10'b1000000100: data <= 12'hffe; 
        10'b1000000101: data <= 12'h000; 
        10'b1000000110: data <= 12'h005; 
        10'b1000000111: data <= 12'hffa; 
        10'b1000001000: data <= 12'hff9; 
        10'b1000001001: data <= 12'hffc; 
        10'b1000001010: data <= 12'hff7; 
        10'b1000001011: data <= 12'hffb; 
        10'b1000001100: data <= 12'hff7; 
        10'b1000001101: data <= 12'hff2; 
        10'b1000001110: data <= 12'hff6; 
        10'b1000001111: data <= 12'hffa; 
        10'b1000010000: data <= 12'hffb; 
        10'b1000010001: data <= 12'h001; 
        10'b1000010010: data <= 12'hfff; 
        10'b1000010011: data <= 12'h000; 
        10'b1000010100: data <= 12'h003; 
        10'b1000010101: data <= 12'h003; 
        10'b1000010110: data <= 12'h003; 
        10'b1000010111: data <= 12'h001; 
        10'b1000011000: data <= 12'hffe; 
        10'b1000011001: data <= 12'hff5; 
        10'b1000011010: data <= 12'hfef; 
        10'b1000011011: data <= 12'hfee; 
        10'b1000011100: data <= 12'hfed; 
        10'b1000011101: data <= 12'hfed; 
        10'b1000011110: data <= 12'hff3; 
        10'b1000011111: data <= 12'hff7; 
        10'b1000100000: data <= 12'hffa; 
        10'b1000100001: data <= 12'h002; 
        10'b1000100010: data <= 12'h008; 
        10'b1000100011: data <= 12'hff8; 
        10'b1000100100: data <= 12'hff8; 
        10'b1000100101: data <= 12'hff6; 
        10'b1000100110: data <= 12'hff1; 
        10'b1000100111: data <= 12'hff1; 
        10'b1000101000: data <= 12'hfee; 
        10'b1000101001: data <= 12'hfef; 
        10'b1000101010: data <= 12'hff3; 
        10'b1000101011: data <= 12'hff7; 
        10'b1000101100: data <= 12'hffc; 
        10'b1000101101: data <= 12'hffe; 
        10'b1000101110: data <= 12'h003; 
        10'b1000101111: data <= 12'hfff; 
        10'b1000110000: data <= 12'hfff; 
        10'b1000110001: data <= 12'hfff; 
        10'b1000110010: data <= 12'h001; 
        10'b1000110011: data <= 12'h000; 
        10'b1000110100: data <= 12'hffd; 
        10'b1000110101: data <= 12'hff8; 
        10'b1000110110: data <= 12'hfef; 
        10'b1000110111: data <= 12'hfee; 
        10'b1000111000: data <= 12'hfef; 
        10'b1000111001: data <= 12'hfef; 
        10'b1000111010: data <= 12'hff4; 
        10'b1000111011: data <= 12'hff4; 
        10'b1000111100: data <= 12'h001; 
        10'b1000111101: data <= 12'h001; 
        10'b1000111110: data <= 12'h004; 
        10'b1000111111: data <= 12'hff5; 
        10'b1001000000: data <= 12'hff3; 
        10'b1001000001: data <= 12'hfef; 
        10'b1001000010: data <= 12'hfe8; 
        10'b1001000011: data <= 12'hff1; 
        10'b1001000100: data <= 12'hfeb; 
        10'b1001000101: data <= 12'hff0; 
        10'b1001000110: data <= 12'hff4; 
        10'b1001000111: data <= 12'hffb; 
        10'b1001001000: data <= 12'hffd; 
        10'b1001001001: data <= 12'h002; 
        10'b1001001010: data <= 12'h002; 
        10'b1001001011: data <= 12'h002; 
        10'b1001001100: data <= 12'h002; 
        10'b1001001101: data <= 12'h002; 
        10'b1001001110: data <= 12'h001; 
        10'b1001001111: data <= 12'hffd; 
        10'b1001010000: data <= 12'hffe; 
        10'b1001010001: data <= 12'hff9; 
        10'b1001010010: data <= 12'hff7; 
        10'b1001010011: data <= 12'hff4; 
        10'b1001010100: data <= 12'hff5; 
        10'b1001010101: data <= 12'hff9; 
        10'b1001010110: data <= 12'hff6; 
        10'b1001010111: data <= 12'hff8; 
        10'b1001011000: data <= 12'hffd; 
        10'b1001011001: data <= 12'h000; 
        10'b1001011010: data <= 12'hffe; 
        10'b1001011011: data <= 12'hff9; 
        10'b1001011100: data <= 12'hff8; 
        10'b1001011101: data <= 12'hfef; 
        10'b1001011110: data <= 12'hfef; 
        10'b1001011111: data <= 12'hfef; 
        10'b1001100000: data <= 12'hfee; 
        10'b1001100001: data <= 12'hff1; 
        10'b1001100010: data <= 12'hff7; 
        10'b1001100011: data <= 12'hff9; 
        10'b1001100100: data <= 12'h000; 
        10'b1001100101: data <= 12'h001; 
        10'b1001100110: data <= 12'h002; 
        10'b1001100111: data <= 12'h000; 
        10'b1001101000: data <= 12'h001; 
        10'b1001101001: data <= 12'h000; 
        10'b1001101010: data <= 12'h001; 
        10'b1001101011: data <= 12'hffe; 
        10'b1001101100: data <= 12'hfff; 
        10'b1001101101: data <= 12'h001; 
        10'b1001101110: data <= 12'hffd; 
        10'b1001101111: data <= 12'h001; 
        10'b1001110000: data <= 12'h002; 
        10'b1001110001: data <= 12'hffd; 
        10'b1001110010: data <= 12'hff9; 
        10'b1001110011: data <= 12'hff5; 
        10'b1001110100: data <= 12'hff6; 
        10'b1001110101: data <= 12'hffc; 
        10'b1001110110: data <= 12'h001; 
        10'b1001110111: data <= 12'h001; 
        10'b1001111000: data <= 12'hffa; 
        10'b1001111001: data <= 12'hff8; 
        10'b1001111010: data <= 12'hff2; 
        10'b1001111011: data <= 12'hff2; 
        10'b1001111100: data <= 12'hff1; 
        10'b1001111101: data <= 12'hff3; 
        10'b1001111110: data <= 12'hff9; 
        10'b1001111111: data <= 12'hffe; 
        10'b1010000000: data <= 12'h001; 
        10'b1010000001: data <= 12'hfff; 
        10'b1010000010: data <= 12'h001; 
        10'b1010000011: data <= 12'h000; 
        10'b1010000100: data <= 12'h001; 
        10'b1010000101: data <= 12'h002; 
        10'b1010000110: data <= 12'hffe; 
        10'b1010000111: data <= 12'hfff; 
        10'b1010001000: data <= 12'h003; 
        10'b1010001001: data <= 12'h004; 
        10'b1010001010: data <= 12'h008; 
        10'b1010001011: data <= 12'h00b; 
        10'b1010001100: data <= 12'h005; 
        10'b1010001101: data <= 12'h001; 
        10'b1010001110: data <= 12'hffd; 
        10'b1010001111: data <= 12'hff9; 
        10'b1010010000: data <= 12'hffa; 
        10'b1010010001: data <= 12'h000; 
        10'b1010010010: data <= 12'h004; 
        10'b1010010011: data <= 12'h004; 
        10'b1010010100: data <= 12'hffe; 
        10'b1010010101: data <= 12'hffe; 
        10'b1010010110: data <= 12'hff7; 
        10'b1010010111: data <= 12'hff4; 
        10'b1010011000: data <= 12'hff4; 
        10'b1010011001: data <= 12'hff6; 
        10'b1010011010: data <= 12'hff8; 
        10'b1010011011: data <= 12'hffb; 
        10'b1010011100: data <= 12'hffe; 
        10'b1010011101: data <= 12'h000; 
        10'b1010011110: data <= 12'h000; 
        10'b1010011111: data <= 12'hfff; 
        10'b1010100000: data <= 12'h000; 
        10'b1010100001: data <= 12'h000; 
        10'b1010100010: data <= 12'h001; 
        10'b1010100011: data <= 12'h002; 
        10'b1010100100: data <= 12'h004; 
        10'b1010100101: data <= 12'h009; 
        10'b1010100110: data <= 12'h00e; 
        10'b1010100111: data <= 12'h00f; 
        10'b1010101000: data <= 12'h00d; 
        10'b1010101001: data <= 12'h007; 
        10'b1010101010: data <= 12'h00e; 
        10'b1010101011: data <= 12'h009; 
        10'b1010101100: data <= 12'h007; 
        10'b1010101101: data <= 12'h00a; 
        10'b1010101110: data <= 12'h006; 
        10'b1010101111: data <= 12'h009; 
        10'b1010110000: data <= 12'h005; 
        10'b1010110001: data <= 12'h004; 
        10'b1010110010: data <= 12'h000; 
        10'b1010110011: data <= 12'hffc; 
        10'b1010110100: data <= 12'hffc; 
        10'b1010110101: data <= 12'hffb; 
        10'b1010110110: data <= 12'hffa; 
        10'b1010110111: data <= 12'hffb; 
        10'b1010111000: data <= 12'h001; 
        10'b1010111001: data <= 12'h000; 
        10'b1010111010: data <= 12'hfff; 
        10'b1010111011: data <= 12'h002; 
        10'b1010111100: data <= 12'hfff; 
        10'b1010111101: data <= 12'h001; 
        10'b1010111110: data <= 12'h002; 
        10'b1010111111: data <= 12'h002; 
        10'b1011000000: data <= 12'h001; 
        10'b1011000001: data <= 12'h004; 
        10'b1011000010: data <= 12'h007; 
        10'b1011000011: data <= 12'h00a; 
        10'b1011000100: data <= 12'h010; 
        10'b1011000101: data <= 12'h00f; 
        10'b1011000110: data <= 12'h012; 
        10'b1011000111: data <= 12'h011; 
        10'b1011001000: data <= 12'h00f; 
        10'b1011001001: data <= 12'h00c; 
        10'b1011001010: data <= 12'h00c; 
        10'b1011001011: data <= 12'h00d; 
        10'b1011001100: data <= 12'h00b; 
        10'b1011001101: data <= 12'h00a; 
        10'b1011001110: data <= 12'h008; 
        10'b1011001111: data <= 12'h003; 
        10'b1011010000: data <= 12'hffd; 
        10'b1011010001: data <= 12'h000; 
        10'b1011010010: data <= 12'hffe; 
        10'b1011010011: data <= 12'hfff; 
        10'b1011010100: data <= 12'h000; 
        10'b1011010101: data <= 12'h001; 
        10'b1011010110: data <= 12'h003; 
        10'b1011010111: data <= 12'h002; 
        10'b1011011000: data <= 12'hfff; 
        10'b1011011001: data <= 12'h001; 
        10'b1011011010: data <= 12'h003; 
        10'b1011011011: data <= 12'h000; 
        10'b1011011100: data <= 12'hfff; 
        10'b1011011101: data <= 12'h003; 
        10'b1011011110: data <= 12'h000; 
        10'b1011011111: data <= 12'h003; 
        10'b1011100000: data <= 12'h002; 
        10'b1011100001: data <= 12'h000; 
        10'b1011100010: data <= 12'h003; 
        10'b1011100011: data <= 12'h005; 
        10'b1011100100: data <= 12'h001; 
        10'b1011100101: data <= 12'h004; 
        10'b1011100110: data <= 12'h009; 
        10'b1011100111: data <= 12'h00c; 
        10'b1011101000: data <= 12'h009; 
        10'b1011101001: data <= 12'h00c; 
        10'b1011101010: data <= 12'h007; 
        10'b1011101011: data <= 12'h003; 
        10'b1011101100: data <= 12'h000; 
        10'b1011101101: data <= 12'h001; 
        10'b1011101110: data <= 12'h000; 
        10'b1011101111: data <= 12'h001; 
        10'b1011110000: data <= 12'h000; 
        10'b1011110001: data <= 12'hfff; 
        10'b1011110010: data <= 12'h000; 
        10'b1011110011: data <= 12'h000; 
        10'b1011110100: data <= 12'hfff; 
        10'b1011110101: data <= 12'h001; 
        10'b1011110110: data <= 12'h001; 
        10'b1011110111: data <= 12'h001; 
        10'b1011111000: data <= 12'h002; 
        10'b1011111001: data <= 12'h001; 
        10'b1011111010: data <= 12'h001; 
        10'b1011111011: data <= 12'h000; 
        10'b1011111100: data <= 12'h003; 
        10'b1011111101: data <= 12'h002; 
        10'b1011111110: data <= 12'h001; 
        10'b1011111111: data <= 12'h002; 
        10'b1100000000: data <= 12'h001; 
        10'b1100000001: data <= 12'h004; 
        10'b1100000010: data <= 12'h002; 
        10'b1100000011: data <= 12'h002; 
        10'b1100000100: data <= 12'h005; 
        10'b1100000101: data <= 12'h002; 
        10'b1100000110: data <= 12'h002; 
        10'b1100000111: data <= 12'h004; 
        10'b1100001000: data <= 12'h000; 
        10'b1100001001: data <= 12'hfff; 
        10'b1100001010: data <= 12'h003; 
        10'b1100001011: data <= 12'h002; 
        10'b1100001100: data <= 12'h001; 
        10'b1100001101: data <= 12'hfff; 
        10'b1100001110: data <= 12'hfff; 
        10'b1100001111: data <= 12'h002; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 7) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 13'h0000; 
        10'b0000000001: data <= 13'h0001; 
        10'b0000000010: data <= 13'h0004; 
        10'b0000000011: data <= 13'h0001; 
        10'b0000000100: data <= 13'h0006; 
        10'b0000000101: data <= 13'h1ffd; 
        10'b0000000110: data <= 13'h1ffe; 
        10'b0000000111: data <= 13'h0002; 
        10'b0000001000: data <= 13'h0005; 
        10'b0000001001: data <= 13'h0005; 
        10'b0000001010: data <= 13'h1ffd; 
        10'b0000001011: data <= 13'h0001; 
        10'b0000001100: data <= 13'h0001; 
        10'b0000001101: data <= 13'h1fff; 
        10'b0000001110: data <= 13'h0005; 
        10'b0000001111: data <= 13'h0001; 
        10'b0000010000: data <= 13'h0000; 
        10'b0000010001: data <= 13'h0000; 
        10'b0000010010: data <= 13'h0001; 
        10'b0000010011: data <= 13'h0002; 
        10'b0000010100: data <= 13'h0003; 
        10'b0000010101: data <= 13'h0006; 
        10'b0000010110: data <= 13'h1ffe; 
        10'b0000010111: data <= 13'h0004; 
        10'b0000011000: data <= 13'h1fff; 
        10'b0000011001: data <= 13'h0003; 
        10'b0000011010: data <= 13'h0000; 
        10'b0000011011: data <= 13'h0000; 
        10'b0000011100: data <= 13'h0006; 
        10'b0000011101: data <= 13'h1fff; 
        10'b0000011110: data <= 13'h0001; 
        10'b0000011111: data <= 13'h0006; 
        10'b0000100000: data <= 13'h0002; 
        10'b0000100001: data <= 13'h0000; 
        10'b0000100010: data <= 13'h0006; 
        10'b0000100011: data <= 13'h0002; 
        10'b0000100100: data <= 13'h0001; 
        10'b0000100101: data <= 13'h1fff; 
        10'b0000100110: data <= 13'h1fff; 
        10'b0000100111: data <= 13'h1ffd; 
        10'b0000101000: data <= 13'h0005; 
        10'b0000101001: data <= 13'h0000; 
        10'b0000101010: data <= 13'h0006; 
        10'b0000101011: data <= 13'h1ffe; 
        10'b0000101100: data <= 13'h0002; 
        10'b0000101101: data <= 13'h0004; 
        10'b0000101110: data <= 13'h0005; 
        10'b0000101111: data <= 13'h0004; 
        10'b0000110000: data <= 13'h0000; 
        10'b0000110001: data <= 13'h0004; 
        10'b0000110010: data <= 13'h0000; 
        10'b0000110011: data <= 13'h0006; 
        10'b0000110100: data <= 13'h0005; 
        10'b0000110101: data <= 13'h1ffe; 
        10'b0000110110: data <= 13'h1ffe; 
        10'b0000110111: data <= 13'h0002; 
        10'b0000111000: data <= 13'h0005; 
        10'b0000111001: data <= 13'h0005; 
        10'b0000111010: data <= 13'h0004; 
        10'b0000111011: data <= 13'h1fff; 
        10'b0000111100: data <= 13'h0005; 
        10'b0000111101: data <= 13'h1ffe; 
        10'b0000111110: data <= 13'h1ffe; 
        10'b0000111111: data <= 13'h0004; 
        10'b0001000000: data <= 13'h0003; 
        10'b0001000001: data <= 13'h1ffe; 
        10'b0001000010: data <= 13'h0000; 
        10'b0001000011: data <= 13'h0002; 
        10'b0001000100: data <= 13'h1fff; 
        10'b0001000101: data <= 13'h1fff; 
        10'b0001000110: data <= 13'h0001; 
        10'b0001000111: data <= 13'h0005; 
        10'b0001001000: data <= 13'h0004; 
        10'b0001001001: data <= 13'h0001; 
        10'b0001001010: data <= 13'h0002; 
        10'b0001001011: data <= 13'h0006; 
        10'b0001001100: data <= 13'h0005; 
        10'b0001001101: data <= 13'h0005; 
        10'b0001001110: data <= 13'h1ffd; 
        10'b0001001111: data <= 13'h0004; 
        10'b0001010000: data <= 13'h0002; 
        10'b0001010001: data <= 13'h0004; 
        10'b0001010010: data <= 13'h0003; 
        10'b0001010011: data <= 13'h0005; 
        10'b0001010100: data <= 13'h0000; 
        10'b0001010101: data <= 13'h0000; 
        10'b0001010110: data <= 13'h0005; 
        10'b0001010111: data <= 13'h1fff; 
        10'b0001011000: data <= 13'h0001; 
        10'b0001011001: data <= 13'h0000; 
        10'b0001011010: data <= 13'h1ffe; 
        10'b0001011011: data <= 13'h0003; 
        10'b0001011100: data <= 13'h0000; 
        10'b0001011101: data <= 13'h0003; 
        10'b0001011110: data <= 13'h1ffd; 
        10'b0001011111: data <= 13'h0001; 
        10'b0001100000: data <= 13'h0003; 
        10'b0001100001: data <= 13'h1ffc; 
        10'b0001100010: data <= 13'h0003; 
        10'b0001100011: data <= 13'h1ffe; 
        10'b0001100100: data <= 13'h1ffb; 
        10'b0001100101: data <= 13'h1ffc; 
        10'b0001100110: data <= 13'h1ffc; 
        10'b0001100111: data <= 13'h1ffe; 
        10'b0001101000: data <= 13'h1fff; 
        10'b0001101001: data <= 13'h1ffe; 
        10'b0001101010: data <= 13'h0002; 
        10'b0001101011: data <= 13'h0000; 
        10'b0001101100: data <= 13'h0002; 
        10'b0001101101: data <= 13'h0006; 
        10'b0001101110: data <= 13'h1ffe; 
        10'b0001101111: data <= 13'h0003; 
        10'b0001110000: data <= 13'h0006; 
        10'b0001110001: data <= 13'h1ffe; 
        10'b0001110010: data <= 13'h0003; 
        10'b0001110011: data <= 13'h1ffd; 
        10'b0001110100: data <= 13'h0001; 
        10'b0001110101: data <= 13'h1fff; 
        10'b0001110110: data <= 13'h0000; 
        10'b0001110111: data <= 13'h1ffe; 
        10'b0001111000: data <= 13'h0002; 
        10'b0001111001: data <= 13'h1fff; 
        10'b0001111010: data <= 13'h1ffa; 
        10'b0001111011: data <= 13'h1ff5; 
        10'b0001111100: data <= 13'h1ff4; 
        10'b0001111101: data <= 13'h1ff5; 
        10'b0001111110: data <= 13'h1ff3; 
        10'b0001111111: data <= 13'h1fea; 
        10'b0010000000: data <= 13'h1ff3; 
        10'b0010000001: data <= 13'h1ff6; 
        10'b0010000010: data <= 13'h1ff8; 
        10'b0010000011: data <= 13'h1ffe; 
        10'b0010000100: data <= 13'h1ffa; 
        10'b0010000101: data <= 13'h0003; 
        10'b0010000110: data <= 13'h0000; 
        10'b0010000111: data <= 13'h1ffd; 
        10'b0010001000: data <= 13'h0006; 
        10'b0010001001: data <= 13'h0000; 
        10'b0010001010: data <= 13'h0005; 
        10'b0010001011: data <= 13'h0005; 
        10'b0010001100: data <= 13'h0005; 
        10'b0010001101: data <= 13'h0000; 
        10'b0010001110: data <= 13'h0005; 
        10'b0010001111: data <= 13'h1fff; 
        10'b0010010000: data <= 13'h1ffc; 
        10'b0010010001: data <= 13'h1fff; 
        10'b0010010010: data <= 13'h1ffd; 
        10'b0010010011: data <= 13'h1fff; 
        10'b0010010100: data <= 13'h1ffd; 
        10'b0010010101: data <= 13'h1ff8; 
        10'b0010010110: data <= 13'h1fec; 
        10'b0010010111: data <= 13'h1fe8; 
        10'b0010011000: data <= 13'h1fe2; 
        10'b0010011001: data <= 13'h1fdc; 
        10'b0010011010: data <= 13'h1fd4; 
        10'b0010011011: data <= 13'h1fd4; 
        10'b0010011100: data <= 13'h1fd2; 
        10'b0010011101: data <= 13'h1fd7; 
        10'b0010011110: data <= 13'h1fdd; 
        10'b0010011111: data <= 13'h1fe6; 
        10'b0010100000: data <= 13'h1fed; 
        10'b0010100001: data <= 13'h1ff9; 
        10'b0010100010: data <= 13'h1ff6; 
        10'b0010100011: data <= 13'h1fff; 
        10'b0010100100: data <= 13'h0005; 
        10'b0010100101: data <= 13'h0004; 
        10'b0010100110: data <= 13'h1fff; 
        10'b0010100111: data <= 13'h0000; 
        10'b0010101000: data <= 13'h0004; 
        10'b0010101001: data <= 13'h0006; 
        10'b0010101010: data <= 13'h0000; 
        10'b0010101011: data <= 13'h0001; 
        10'b0010101100: data <= 13'h0006; 
        10'b0010101101: data <= 13'h0007; 
        10'b0010101110: data <= 13'h0009; 
        10'b0010101111: data <= 13'h000d; 
        10'b0010110000: data <= 13'h0013; 
        10'b0010110001: data <= 13'h000f; 
        10'b0010110010: data <= 13'h0010; 
        10'b0010110011: data <= 13'h0003; 
        10'b0010110100: data <= 13'h1ff3; 
        10'b0010110101: data <= 13'h1fe4; 
        10'b0010110110: data <= 13'h1fe3; 
        10'b0010110111: data <= 13'h1ff1; 
        10'b0010111000: data <= 13'h1ff7; 
        10'b0010111001: data <= 13'h1ff5; 
        10'b0010111010: data <= 13'h1ff3; 
        10'b0010111011: data <= 13'h1ff1; 
        10'b0010111100: data <= 13'h1fe9; 
        10'b0010111101: data <= 13'h1ff7; 
        10'b0010111110: data <= 13'h1ff0; 
        10'b0010111111: data <= 13'h1ff4; 
        10'b0011000000: data <= 13'h1ff8; 
        10'b0011000001: data <= 13'h1ffd; 
        10'b0011000010: data <= 13'h1ffd; 
        10'b0011000011: data <= 13'h0001; 
        10'b0011000100: data <= 13'h0004; 
        10'b0011000101: data <= 13'h0006; 
        10'b0011000110: data <= 13'h0005; 
        10'b0011000111: data <= 13'h000b; 
        10'b0011001000: data <= 13'h000e; 
        10'b0011001001: data <= 13'h000c; 
        10'b0011001010: data <= 13'h0012; 
        10'b0011001011: data <= 13'h001b; 
        10'b0011001100: data <= 13'h0025; 
        10'b0011001101: data <= 13'h001d; 
        10'b0011001110: data <= 13'h0014; 
        10'b0011001111: data <= 13'h0016; 
        10'b0011010000: data <= 13'h0018; 
        10'b0011010001: data <= 13'h0005; 
        10'b0011010010: data <= 13'h0003; 
        10'b0011010011: data <= 13'h0009; 
        10'b0011010100: data <= 13'h0019; 
        10'b0011010101: data <= 13'h001c; 
        10'b0011010110: data <= 13'h0013; 
        10'b0011010111: data <= 13'h000f; 
        10'b0011011000: data <= 13'h0004; 
        10'b0011011001: data <= 13'h1ffc; 
        10'b0011011010: data <= 13'h0002; 
        10'b0011011011: data <= 13'h1ffb; 
        10'b0011011100: data <= 13'h1ffc; 
        10'b0011011101: data <= 13'h0000; 
        10'b0011011110: data <= 13'h0003; 
        10'b0011011111: data <= 13'h1fff; 
        10'b0011100000: data <= 13'h1ffd; 
        10'b0011100001: data <= 13'h0006; 
        10'b0011100010: data <= 13'h0002; 
        10'b0011100011: data <= 13'h000a; 
        10'b0011100100: data <= 13'h0013; 
        10'b0011100101: data <= 13'h0011; 
        10'b0011100110: data <= 13'h0017; 
        10'b0011100111: data <= 13'h002a; 
        10'b0011101000: data <= 13'h001c; 
        10'b0011101001: data <= 13'h0013; 
        10'b0011101010: data <= 13'h0019; 
        10'b0011101011: data <= 13'h0021; 
        10'b0011101100: data <= 13'h001f; 
        10'b0011101101: data <= 13'h0010; 
        10'b0011101110: data <= 13'h0009; 
        10'b0011101111: data <= 13'h000d; 
        10'b0011110000: data <= 13'h0016; 
        10'b0011110001: data <= 13'h0022; 
        10'b0011110010: data <= 13'h0017; 
        10'b0011110011: data <= 13'h0014; 
        10'b0011110100: data <= 13'h0010; 
        10'b0011110101: data <= 13'h0000; 
        10'b0011110110: data <= 13'h000a; 
        10'b0011110111: data <= 13'h0008; 
        10'b0011111000: data <= 13'h1ffa; 
        10'b0011111001: data <= 13'h1ffd; 
        10'b0011111010: data <= 13'h0003; 
        10'b0011111011: data <= 13'h0005; 
        10'b0011111100: data <= 13'h0003; 
        10'b0011111101: data <= 13'h0005; 
        10'b0011111110: data <= 13'h0006; 
        10'b0011111111: data <= 13'h000e; 
        10'b0100000000: data <= 13'h0013; 
        10'b0100000001: data <= 13'h0015; 
        10'b0100000010: data <= 13'h0008; 
        10'b0100000011: data <= 13'h000a; 
        10'b0100000100: data <= 13'h000c; 
        10'b0100000101: data <= 13'h0008; 
        10'b0100000110: data <= 13'h0013; 
        10'b0100000111: data <= 13'h0018; 
        10'b0100001000: data <= 13'h001e; 
        10'b0100001001: data <= 13'h0018; 
        10'b0100001010: data <= 13'h0023; 
        10'b0100001011: data <= 13'h002b; 
        10'b0100001100: data <= 13'h0028; 
        10'b0100001101: data <= 13'h002c; 
        10'b0100001110: data <= 13'h001d; 
        10'b0100001111: data <= 13'h001d; 
        10'b0100010000: data <= 13'h0019; 
        10'b0100010001: data <= 13'h0015; 
        10'b0100010010: data <= 13'h000a; 
        10'b0100010011: data <= 13'h1ffc; 
        10'b0100010100: data <= 13'h1ffa; 
        10'b0100010101: data <= 13'h1ffd; 
        10'b0100010110: data <= 13'h0003; 
        10'b0100010111: data <= 13'h1fff; 
        10'b0100011000: data <= 13'h0001; 
        10'b0100011001: data <= 13'h0005; 
        10'b0100011010: data <= 13'h0006; 
        10'b0100011011: data <= 13'h0011; 
        10'b0100011100: data <= 13'h0014; 
        10'b0100011101: data <= 13'h0010; 
        10'b0100011110: data <= 13'h0003; 
        10'b0100011111: data <= 13'h0005; 
        10'b0100100000: data <= 13'h1ff9; 
        10'b0100100001: data <= 13'h0000; 
        10'b0100100010: data <= 13'h000c; 
        10'b0100100011: data <= 13'h0015; 
        10'b0100100100: data <= 13'h000f; 
        10'b0100100101: data <= 13'h0022; 
        10'b0100100110: data <= 13'h002c; 
        10'b0100100111: data <= 13'h0036; 
        10'b0100101000: data <= 13'h003d; 
        10'b0100101001: data <= 13'h002d; 
        10'b0100101010: data <= 13'h0024; 
        10'b0100101011: data <= 13'h0025; 
        10'b0100101100: data <= 13'h0021; 
        10'b0100101101: data <= 13'h001c; 
        10'b0100101110: data <= 13'h000c; 
        10'b0100101111: data <= 13'h1ffb; 
        10'b0100110000: data <= 13'h1ff8; 
        10'b0100110001: data <= 13'h1ffd; 
        10'b0100110010: data <= 13'h0001; 
        10'b0100110011: data <= 13'h1fff; 
        10'b0100110100: data <= 13'h0005; 
        10'b0100110101: data <= 13'h0003; 
        10'b0100110110: data <= 13'h0006; 
        10'b0100110111: data <= 13'h0011; 
        10'b0100111000: data <= 13'h0015; 
        10'b0100111001: data <= 13'h000a; 
        10'b0100111010: data <= 13'h0004; 
        10'b0100111011: data <= 13'h0003; 
        10'b0100111100: data <= 13'h0001; 
        10'b0100111101: data <= 13'h000d; 
        10'b0100111110: data <= 13'h0007; 
        10'b0100111111: data <= 13'h0008; 
        10'b0101000000: data <= 13'h000e; 
        10'b0101000001: data <= 13'h000d; 
        10'b0101000010: data <= 13'h000e; 
        10'b0101000011: data <= 13'h0029; 
        10'b0101000100: data <= 13'h0035; 
        10'b0101000101: data <= 13'h0024; 
        10'b0101000110: data <= 13'h0024; 
        10'b0101000111: data <= 13'h001c; 
        10'b0101001000: data <= 13'h001b; 
        10'b0101001001: data <= 13'h0011; 
        10'b0101001010: data <= 13'h000c; 
        10'b0101001011: data <= 13'h1ffc; 
        10'b0101001100: data <= 13'h1ff4; 
        10'b0101001101: data <= 13'h0000; 
        10'b0101001110: data <= 13'h0001; 
        10'b0101001111: data <= 13'h0005; 
        10'b0101010000: data <= 13'h0004; 
        10'b0101010001: data <= 13'h0000; 
        10'b0101010010: data <= 13'h0003; 
        10'b0101010011: data <= 13'h000b; 
        10'b0101010100: data <= 13'h000c; 
        10'b0101010101: data <= 13'h0002; 
        10'b0101010110: data <= 13'h0003; 
        10'b0101010111: data <= 13'h000c; 
        10'b0101011000: data <= 13'h0008; 
        10'b0101011001: data <= 13'h0000; 
        10'b0101011010: data <= 13'h1ff6; 
        10'b0101011011: data <= 13'h1fe6; 
        10'b0101011100: data <= 13'h1fca; 
        10'b0101011101: data <= 13'h1fac; 
        10'b0101011110: data <= 13'h1fc1; 
        10'b0101011111: data <= 13'h0001; 
        10'b0101100000: data <= 13'h0023; 
        10'b0101100001: data <= 13'h0020; 
        10'b0101100010: data <= 13'h000d; 
        10'b0101100011: data <= 13'h0005; 
        10'b0101100100: data <= 13'h0001; 
        10'b0101100101: data <= 13'h1ffb; 
        10'b0101100110: data <= 13'h1ffc; 
        10'b0101100111: data <= 13'h1ff8; 
        10'b0101101000: data <= 13'h1ffb; 
        10'b0101101001: data <= 13'h0005; 
        10'b0101101010: data <= 13'h0004; 
        10'b0101101011: data <= 13'h0000; 
        10'b0101101100: data <= 13'h0004; 
        10'b0101101101: data <= 13'h0003; 
        10'b0101101110: data <= 13'h0005; 
        10'b0101101111: data <= 13'h000a; 
        10'b0101110000: data <= 13'h0004; 
        10'b0101110001: data <= 13'h0002; 
        10'b0101110010: data <= 13'h1ffd; 
        10'b0101110011: data <= 13'h0002; 
        10'b0101110100: data <= 13'h1ffe; 
        10'b0101110101: data <= 13'h1ff8; 
        10'b0101110110: data <= 13'h1fe5; 
        10'b0101110111: data <= 13'h1fc7; 
        10'b0101111000: data <= 13'h1f9d; 
        10'b0101111001: data <= 13'h1f91; 
        10'b0101111010: data <= 13'h1fc5; 
        10'b0101111011: data <= 13'h1ff8; 
        10'b0101111100: data <= 13'h0012; 
        10'b0101111101: data <= 13'h000c; 
        10'b0101111110: data <= 13'h0003; 
        10'b0101111111: data <= 13'h0005; 
        10'b0110000000: data <= 13'h1ff5; 
        10'b0110000001: data <= 13'h1ff2; 
        10'b0110000010: data <= 13'h1ffd; 
        10'b0110000011: data <= 13'h0001; 
        10'b0110000100: data <= 13'h1ffd; 
        10'b0110000101: data <= 13'h1ffe; 
        10'b0110000110: data <= 13'h0003; 
        10'b0110000111: data <= 13'h1ffd; 
        10'b0110001000: data <= 13'h1fff; 
        10'b0110001001: data <= 13'h0002; 
        10'b0110001010: data <= 13'h0009; 
        10'b0110001011: data <= 13'h000b; 
        10'b0110001100: data <= 13'h0007; 
        10'b0110001101: data <= 13'h0008; 
        10'b0110001110: data <= 13'h1ffd; 
        10'b0110001111: data <= 13'h1ffa; 
        10'b0110010000: data <= 13'h1ff3; 
        10'b0110010001: data <= 13'h1fe3; 
        10'b0110010010: data <= 13'h1fd5; 
        10'b0110010011: data <= 13'h1fbd; 
        10'b0110010100: data <= 13'h1faa; 
        10'b0110010101: data <= 13'h1fb8; 
        10'b0110010110: data <= 13'h1fe5; 
        10'b0110010111: data <= 13'h0001; 
        10'b0110011000: data <= 13'h0006; 
        10'b0110011001: data <= 13'h000b; 
        10'b0110011010: data <= 13'h0021; 
        10'b0110011011: data <= 13'h0023; 
        10'b0110011100: data <= 13'h0015; 
        10'b0110011101: data <= 13'h000e; 
        10'b0110011110: data <= 13'h000e; 
        10'b0110011111: data <= 13'h000c; 
        10'b0110100000: data <= 13'h0004; 
        10'b0110100001: data <= 13'h0001; 
        10'b0110100010: data <= 13'h1ffe; 
        10'b0110100011: data <= 13'h1ffe; 
        10'b0110100100: data <= 13'h0003; 
        10'b0110100101: data <= 13'h0004; 
        10'b0110100110: data <= 13'h0002; 
        10'b0110100111: data <= 13'h0004; 
        10'b0110101000: data <= 13'h0004; 
        10'b0110101001: data <= 13'h1ff4; 
        10'b0110101010: data <= 13'h1ffb; 
        10'b0110101011: data <= 13'h1ff9; 
        10'b0110101100: data <= 13'h1fe0; 
        10'b0110101101: data <= 13'h1fda; 
        10'b0110101110: data <= 13'h1fcd; 
        10'b0110101111: data <= 13'h1fc6; 
        10'b0110110000: data <= 13'h1fc0; 
        10'b0110110001: data <= 13'h1fd1; 
        10'b0110110010: data <= 13'h1fe5; 
        10'b0110110011: data <= 13'h0001; 
        10'b0110110100: data <= 13'h0003; 
        10'b0110110101: data <= 13'h002d; 
        10'b0110110110: data <= 13'h0034; 
        10'b0110110111: data <= 13'h002b; 
        10'b0110111000: data <= 13'h0026; 
        10'b0110111001: data <= 13'h0021; 
        10'b0110111010: data <= 13'h0015; 
        10'b0110111011: data <= 13'h000a; 
        10'b0110111100: data <= 13'h0000; 
        10'b0110111101: data <= 13'h1ffd; 
        10'b0110111110: data <= 13'h0001; 
        10'b0110111111: data <= 13'h0005; 
        10'b0111000000: data <= 13'h0003; 
        10'b0111000001: data <= 13'h0006; 
        10'b0111000010: data <= 13'h0000; 
        10'b0111000011: data <= 13'h0006; 
        10'b0111000100: data <= 13'h0005; 
        10'b0111000101: data <= 13'h1ffb; 
        10'b0111000110: data <= 13'h1ff8; 
        10'b0111000111: data <= 13'h1fff; 
        10'b0111001000: data <= 13'h1fe7; 
        10'b0111001001: data <= 13'h1fe3; 
        10'b0111001010: data <= 13'h1fd2; 
        10'b0111001011: data <= 13'h1fc9; 
        10'b0111001100: data <= 13'h1fde; 
        10'b0111001101: data <= 13'h1fed; 
        10'b0111001110: data <= 13'h1fe4; 
        10'b0111001111: data <= 13'h000e; 
        10'b0111010000: data <= 13'h0011; 
        10'b0111010001: data <= 13'h0026; 
        10'b0111010010: data <= 13'h0020; 
        10'b0111010011: data <= 13'h0022; 
        10'b0111010100: data <= 13'h001b; 
        10'b0111010101: data <= 13'h0015; 
        10'b0111010110: data <= 13'h0004; 
        10'b0111010111: data <= 13'h1ff8; 
        10'b0111011000: data <= 13'h1ffb; 
        10'b0111011001: data <= 13'h1ffd; 
        10'b0111011010: data <= 13'h0003; 
        10'b0111011011: data <= 13'h0006; 
        10'b0111011100: data <= 13'h0000; 
        10'b0111011101: data <= 13'h0001; 
        10'b0111011110: data <= 13'h0003; 
        10'b0111011111: data <= 13'h0000; 
        10'b0111100000: data <= 13'h0001; 
        10'b0111100001: data <= 13'h1ffd; 
        10'b0111100010: data <= 13'h1fef; 
        10'b0111100011: data <= 13'h1fe9; 
        10'b0111100100: data <= 13'h1fe4; 
        10'b0111100101: data <= 13'h1fe9; 
        10'b0111100110: data <= 13'h1fe1; 
        10'b0111100111: data <= 13'h1fe9; 
        10'b0111101000: data <= 13'h1ff9; 
        10'b0111101001: data <= 13'h0006; 
        10'b0111101010: data <= 13'h0003; 
        10'b0111101011: data <= 13'h0006; 
        10'b0111101100: data <= 13'h1ffd; 
        10'b0111101101: data <= 13'h0009; 
        10'b0111101110: data <= 13'h0008; 
        10'b0111101111: data <= 13'h0006; 
        10'b0111110000: data <= 13'h0003; 
        10'b0111110001: data <= 13'h1ffb; 
        10'b0111110010: data <= 13'h1ff6; 
        10'b0111110011: data <= 13'h1ffb; 
        10'b0111110100: data <= 13'h1ffc; 
        10'b0111110101: data <= 13'h1ffd; 
        10'b0111110110: data <= 13'h1ffe; 
        10'b0111110111: data <= 13'h1ffe; 
        10'b0111111000: data <= 13'h1ffe; 
        10'b0111111001: data <= 13'h1fff; 
        10'b0111111010: data <= 13'h0004; 
        10'b0111111011: data <= 13'h0001; 
        10'b0111111100: data <= 13'h1ff9; 
        10'b0111111101: data <= 13'h1fef; 
        10'b0111111110: data <= 13'h1fe5; 
        10'b0111111111: data <= 13'h1fde; 
        10'b1000000000: data <= 13'h1fe0; 
        10'b1000000001: data <= 13'h1fe2; 
        10'b1000000010: data <= 13'h1fda; 
        10'b1000000011: data <= 13'h1ff3; 
        10'b1000000100: data <= 13'h1ffc; 
        10'b1000000101: data <= 13'h0000; 
        10'b1000000110: data <= 13'h000b; 
        10'b1000000111: data <= 13'h1ff5; 
        10'b1000001000: data <= 13'h1ff2; 
        10'b1000001001: data <= 13'h1ff8; 
        10'b1000001010: data <= 13'h1fef; 
        10'b1000001011: data <= 13'h1ff5; 
        10'b1000001100: data <= 13'h1fee; 
        10'b1000001101: data <= 13'h1fe4; 
        10'b1000001110: data <= 13'h1fec; 
        10'b1000001111: data <= 13'h1ff3; 
        10'b1000010000: data <= 13'h1ff6; 
        10'b1000010001: data <= 13'h0001; 
        10'b1000010010: data <= 13'h1fff; 
        10'b1000010011: data <= 13'h0000; 
        10'b1000010100: data <= 13'h0005; 
        10'b1000010101: data <= 13'h0006; 
        10'b1000010110: data <= 13'h0005; 
        10'b1000010111: data <= 13'h0003; 
        10'b1000011000: data <= 13'h1ffb; 
        10'b1000011001: data <= 13'h1feb; 
        10'b1000011010: data <= 13'h1fde; 
        10'b1000011011: data <= 13'h1fdb; 
        10'b1000011100: data <= 13'h1fda; 
        10'b1000011101: data <= 13'h1fda; 
        10'b1000011110: data <= 13'h1fe6; 
        10'b1000011111: data <= 13'h1fed; 
        10'b1000100000: data <= 13'h1ff5; 
        10'b1000100001: data <= 13'h0005; 
        10'b1000100010: data <= 13'h000f; 
        10'b1000100011: data <= 13'h1ff0; 
        10'b1000100100: data <= 13'h1ff1; 
        10'b1000100101: data <= 13'h1fed; 
        10'b1000100110: data <= 13'h1fe1; 
        10'b1000100111: data <= 13'h1fe3; 
        10'b1000101000: data <= 13'h1fdc; 
        10'b1000101001: data <= 13'h1fdf; 
        10'b1000101010: data <= 13'h1fe7; 
        10'b1000101011: data <= 13'h1fef; 
        10'b1000101100: data <= 13'h1ff7; 
        10'b1000101101: data <= 13'h1ffd; 
        10'b1000101110: data <= 13'h0006; 
        10'b1000101111: data <= 13'h1ffd; 
        10'b1000110000: data <= 13'h1ffd; 
        10'b1000110001: data <= 13'h1fff; 
        10'b1000110010: data <= 13'h0002; 
        10'b1000110011: data <= 13'h1fff; 
        10'b1000110100: data <= 13'h1ffb; 
        10'b1000110101: data <= 13'h1fef; 
        10'b1000110110: data <= 13'h1fdd; 
        10'b1000110111: data <= 13'h1fdc; 
        10'b1000111000: data <= 13'h1fde; 
        10'b1000111001: data <= 13'h1fdf; 
        10'b1000111010: data <= 13'h1fe9; 
        10'b1000111011: data <= 13'h1fe8; 
        10'b1000111100: data <= 13'h0002; 
        10'b1000111101: data <= 13'h0002; 
        10'b1000111110: data <= 13'h0008; 
        10'b1000111111: data <= 13'h1feb; 
        10'b1001000000: data <= 13'h1fe6; 
        10'b1001000001: data <= 13'h1fdd; 
        10'b1001000010: data <= 13'h1fd0; 
        10'b1001000011: data <= 13'h1fe2; 
        10'b1001000100: data <= 13'h1fd6; 
        10'b1001000101: data <= 13'h1fe0; 
        10'b1001000110: data <= 13'h1fe9; 
        10'b1001000111: data <= 13'h1ff6; 
        10'b1001001000: data <= 13'h1ff9; 
        10'b1001001001: data <= 13'h0005; 
        10'b1001001010: data <= 13'h0005; 
        10'b1001001011: data <= 13'h0003; 
        10'b1001001100: data <= 13'h0004; 
        10'b1001001101: data <= 13'h0005; 
        10'b1001001110: data <= 13'h0001; 
        10'b1001001111: data <= 13'h1ffa; 
        10'b1001010000: data <= 13'h1ffd; 
        10'b1001010001: data <= 13'h1ff1; 
        10'b1001010010: data <= 13'h1fef; 
        10'b1001010011: data <= 13'h1fe7; 
        10'b1001010100: data <= 13'h1fe9; 
        10'b1001010101: data <= 13'h1ff3; 
        10'b1001010110: data <= 13'h1fed; 
        10'b1001010111: data <= 13'h1ff0; 
        10'b1001011000: data <= 13'h1ff9; 
        10'b1001011001: data <= 13'h0001; 
        10'b1001011010: data <= 13'h1ffc; 
        10'b1001011011: data <= 13'h1ff2; 
        10'b1001011100: data <= 13'h1ff0; 
        10'b1001011101: data <= 13'h1fde; 
        10'b1001011110: data <= 13'h1fde; 
        10'b1001011111: data <= 13'h1fde; 
        10'b1001100000: data <= 13'h1fdc; 
        10'b1001100001: data <= 13'h1fe2; 
        10'b1001100010: data <= 13'h1fee; 
        10'b1001100011: data <= 13'h1ff3; 
        10'b1001100100: data <= 13'h1fff; 
        10'b1001100101: data <= 13'h0002; 
        10'b1001100110: data <= 13'h0004; 
        10'b1001100111: data <= 13'h1fff; 
        10'b1001101000: data <= 13'h0002; 
        10'b1001101001: data <= 13'h0000; 
        10'b1001101010: data <= 13'h0001; 
        10'b1001101011: data <= 13'h1ffc; 
        10'b1001101100: data <= 13'h1ffe; 
        10'b1001101101: data <= 13'h0002; 
        10'b1001101110: data <= 13'h1ffb; 
        10'b1001101111: data <= 13'h0003; 
        10'b1001110000: data <= 13'h0004; 
        10'b1001110001: data <= 13'h1ff9; 
        10'b1001110010: data <= 13'h1ff3; 
        10'b1001110011: data <= 13'h1fea; 
        10'b1001110100: data <= 13'h1feb; 
        10'b1001110101: data <= 13'h1ff8; 
        10'b1001110110: data <= 13'h0002; 
        10'b1001110111: data <= 13'h0002; 
        10'b1001111000: data <= 13'h1ff3; 
        10'b1001111001: data <= 13'h1ff0; 
        10'b1001111010: data <= 13'h1fe5; 
        10'b1001111011: data <= 13'h1fe5; 
        10'b1001111100: data <= 13'h1fe1; 
        10'b1001111101: data <= 13'h1fe5; 
        10'b1001111110: data <= 13'h1ff2; 
        10'b1001111111: data <= 13'h1ffb; 
        10'b1010000000: data <= 13'h0003; 
        10'b1010000001: data <= 13'h1ffd; 
        10'b1010000010: data <= 13'h0001; 
        10'b1010000011: data <= 13'h0000; 
        10'b1010000100: data <= 13'h0002; 
        10'b1010000101: data <= 13'h0004; 
        10'b1010000110: data <= 13'h1ffd; 
        10'b1010000111: data <= 13'h1ffd; 
        10'b1010001000: data <= 13'h0006; 
        10'b1010001001: data <= 13'h0008; 
        10'b1010001010: data <= 13'h0010; 
        10'b1010001011: data <= 13'h0016; 
        10'b1010001100: data <= 13'h000a; 
        10'b1010001101: data <= 13'h0002; 
        10'b1010001110: data <= 13'h1ffa; 
        10'b1010001111: data <= 13'h1ff1; 
        10'b1010010000: data <= 13'h1ff4; 
        10'b1010010001: data <= 13'h0001; 
        10'b1010010010: data <= 13'h0009; 
        10'b1010010011: data <= 13'h0008; 
        10'b1010010100: data <= 13'h1ffd; 
        10'b1010010101: data <= 13'h1ffb; 
        10'b1010010110: data <= 13'h1fef; 
        10'b1010010111: data <= 13'h1fe8; 
        10'b1010011000: data <= 13'h1fe7; 
        10'b1010011001: data <= 13'h1fed; 
        10'b1010011010: data <= 13'h1ff0; 
        10'b1010011011: data <= 13'h1ff6; 
        10'b1010011100: data <= 13'h1ffb; 
        10'b1010011101: data <= 13'h0000; 
        10'b1010011110: data <= 13'h0000; 
        10'b1010011111: data <= 13'h1ffe; 
        10'b1010100000: data <= 13'h0000; 
        10'b1010100001: data <= 13'h1fff; 
        10'b1010100010: data <= 13'h0002; 
        10'b1010100011: data <= 13'h0004; 
        10'b1010100100: data <= 13'h0008; 
        10'b1010100101: data <= 13'h0012; 
        10'b1010100110: data <= 13'h001b; 
        10'b1010100111: data <= 13'h001f; 
        10'b1010101000: data <= 13'h001a; 
        10'b1010101001: data <= 13'h000d; 
        10'b1010101010: data <= 13'h001d; 
        10'b1010101011: data <= 13'h0011; 
        10'b1010101100: data <= 13'h000f; 
        10'b1010101101: data <= 13'h0015; 
        10'b1010101110: data <= 13'h000d; 
        10'b1010101111: data <= 13'h0013; 
        10'b1010110000: data <= 13'h000b; 
        10'b1010110001: data <= 13'h0009; 
        10'b1010110010: data <= 13'h1fff; 
        10'b1010110011: data <= 13'h1ff8; 
        10'b1010110100: data <= 13'h1ff7; 
        10'b1010110101: data <= 13'h1ff6; 
        10'b1010110110: data <= 13'h1ff4; 
        10'b1010110111: data <= 13'h1ff5; 
        10'b1010111000: data <= 13'h0002; 
        10'b1010111001: data <= 13'h1fff; 
        10'b1010111010: data <= 13'h1ffd; 
        10'b1010111011: data <= 13'h0003; 
        10'b1010111100: data <= 13'h1ffd; 
        10'b1010111101: data <= 13'h0003; 
        10'b1010111110: data <= 13'h0005; 
        10'b1010111111: data <= 13'h0004; 
        10'b1011000000: data <= 13'h0003; 
        10'b1011000001: data <= 13'h0009; 
        10'b1011000010: data <= 13'h000d; 
        10'b1011000011: data <= 13'h0015; 
        10'b1011000100: data <= 13'h0020; 
        10'b1011000101: data <= 13'h001f; 
        10'b1011000110: data <= 13'h0025; 
        10'b1011000111: data <= 13'h0022; 
        10'b1011001000: data <= 13'h001e; 
        10'b1011001001: data <= 13'h0018; 
        10'b1011001010: data <= 13'h0019; 
        10'b1011001011: data <= 13'h001a; 
        10'b1011001100: data <= 13'h0016; 
        10'b1011001101: data <= 13'h0014; 
        10'b1011001110: data <= 13'h0010; 
        10'b1011001111: data <= 13'h0006; 
        10'b1011010000: data <= 13'h1ff9; 
        10'b1011010001: data <= 13'h0001; 
        10'b1011010010: data <= 13'h1ffd; 
        10'b1011010011: data <= 13'h1ffd; 
        10'b1011010100: data <= 13'h1fff; 
        10'b1011010101: data <= 13'h0002; 
        10'b1011010110: data <= 13'h0006; 
        10'b1011010111: data <= 13'h0004; 
        10'b1011011000: data <= 13'h1ffe; 
        10'b1011011001: data <= 13'h0001; 
        10'b1011011010: data <= 13'h0006; 
        10'b1011011011: data <= 13'h1fff; 
        10'b1011011100: data <= 13'h1ffe; 
        10'b1011011101: data <= 13'h0005; 
        10'b1011011110: data <= 13'h0000; 
        10'b1011011111: data <= 13'h0005; 
        10'b1011100000: data <= 13'h0005; 
        10'b1011100001: data <= 13'h0001; 
        10'b1011100010: data <= 13'h0007; 
        10'b1011100011: data <= 13'h000a; 
        10'b1011100100: data <= 13'h0003; 
        10'b1011100101: data <= 13'h0009; 
        10'b1011100110: data <= 13'h0013; 
        10'b1011100111: data <= 13'h0017; 
        10'b1011101000: data <= 13'h0012; 
        10'b1011101001: data <= 13'h0017; 
        10'b1011101010: data <= 13'h000d; 
        10'b1011101011: data <= 13'h0006; 
        10'b1011101100: data <= 13'h0000; 
        10'b1011101101: data <= 13'h0002; 
        10'b1011101110: data <= 13'h1fff; 
        10'b1011101111: data <= 13'h0001; 
        10'b1011110000: data <= 13'h0000; 
        10'b1011110001: data <= 13'h1ffe; 
        10'b1011110010: data <= 13'h0000; 
        10'b1011110011: data <= 13'h1fff; 
        10'b1011110100: data <= 13'h1ffd; 
        10'b1011110101: data <= 13'h0002; 
        10'b1011110110: data <= 13'h0002; 
        10'b1011110111: data <= 13'h0003; 
        10'b1011111000: data <= 13'h0004; 
        10'b1011111001: data <= 13'h0002; 
        10'b1011111010: data <= 13'h0001; 
        10'b1011111011: data <= 13'h0000; 
        10'b1011111100: data <= 13'h0007; 
        10'b1011111101: data <= 13'h0004; 
        10'b1011111110: data <= 13'h0001; 
        10'b1011111111: data <= 13'h0004; 
        10'b1100000000: data <= 13'h0002; 
        10'b1100000001: data <= 13'h0008; 
        10'b1100000010: data <= 13'h0005; 
        10'b1100000011: data <= 13'h0003; 
        10'b1100000100: data <= 13'h000b; 
        10'b1100000101: data <= 13'h0004; 
        10'b1100000110: data <= 13'h0003; 
        10'b1100000111: data <= 13'h0007; 
        10'b1100001000: data <= 13'h0001; 
        10'b1100001001: data <= 13'h1fff; 
        10'b1100001010: data <= 13'h0006; 
        10'b1100001011: data <= 13'h0003; 
        10'b1100001100: data <= 13'h0002; 
        10'b1100001101: data <= 13'h1fff; 
        10'b1100001110: data <= 13'h1ffe; 
        10'b1100001111: data <= 13'h0004; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 8) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 14'h0001; 
        10'b0000000001: data <= 14'h0001; 
        10'b0000000010: data <= 14'h0008; 
        10'b0000000011: data <= 14'h0003; 
        10'b0000000100: data <= 14'h000c; 
        10'b0000000101: data <= 14'h3ffb; 
        10'b0000000110: data <= 14'h3ffc; 
        10'b0000000111: data <= 14'h0004; 
        10'b0000001000: data <= 14'h000a; 
        10'b0000001001: data <= 14'h0009; 
        10'b0000001010: data <= 14'h3ffb; 
        10'b0000001011: data <= 14'h0002; 
        10'b0000001100: data <= 14'h0003; 
        10'b0000001101: data <= 14'h3fff; 
        10'b0000001110: data <= 14'h000a; 
        10'b0000001111: data <= 14'h0003; 
        10'b0000010000: data <= 14'h0000; 
        10'b0000010001: data <= 14'h0000; 
        10'b0000010010: data <= 14'h0001; 
        10'b0000010011: data <= 14'h0003; 
        10'b0000010100: data <= 14'h0006; 
        10'b0000010101: data <= 14'h000c; 
        10'b0000010110: data <= 14'h3ffd; 
        10'b0000010111: data <= 14'h0009; 
        10'b0000011000: data <= 14'h3fff; 
        10'b0000011001: data <= 14'h0006; 
        10'b0000011010: data <= 14'h3fff; 
        10'b0000011011: data <= 14'h0000; 
        10'b0000011100: data <= 14'h000b; 
        10'b0000011101: data <= 14'h3ffe; 
        10'b0000011110: data <= 14'h0003; 
        10'b0000011111: data <= 14'h000b; 
        10'b0000100000: data <= 14'h0004; 
        10'b0000100001: data <= 14'h0000; 
        10'b0000100010: data <= 14'h000b; 
        10'b0000100011: data <= 14'h0004; 
        10'b0000100100: data <= 14'h0001; 
        10'b0000100101: data <= 14'h3ffe; 
        10'b0000100110: data <= 14'h3fff; 
        10'b0000100111: data <= 14'h3ffa; 
        10'b0000101000: data <= 14'h000a; 
        10'b0000101001: data <= 14'h3fff; 
        10'b0000101010: data <= 14'h000c; 
        10'b0000101011: data <= 14'h3ffd; 
        10'b0000101100: data <= 14'h0005; 
        10'b0000101101: data <= 14'h0009; 
        10'b0000101110: data <= 14'h000a; 
        10'b0000101111: data <= 14'h0008; 
        10'b0000110000: data <= 14'h0000; 
        10'b0000110001: data <= 14'h0008; 
        10'b0000110010: data <= 14'h0000; 
        10'b0000110011: data <= 14'h000c; 
        10'b0000110100: data <= 14'h0009; 
        10'b0000110101: data <= 14'h3ffd; 
        10'b0000110110: data <= 14'h3ffd; 
        10'b0000110111: data <= 14'h0005; 
        10'b0000111000: data <= 14'h000b; 
        10'b0000111001: data <= 14'h000b; 
        10'b0000111010: data <= 14'h0008; 
        10'b0000111011: data <= 14'h3ffe; 
        10'b0000111100: data <= 14'h000a; 
        10'b0000111101: data <= 14'h3ffb; 
        10'b0000111110: data <= 14'h3ffc; 
        10'b0000111111: data <= 14'h0008; 
        10'b0001000000: data <= 14'h0006; 
        10'b0001000001: data <= 14'h3ffc; 
        10'b0001000010: data <= 14'h3fff; 
        10'b0001000011: data <= 14'h0005; 
        10'b0001000100: data <= 14'h3fff; 
        10'b0001000101: data <= 14'h3ffe; 
        10'b0001000110: data <= 14'h0003; 
        10'b0001000111: data <= 14'h000a; 
        10'b0001001000: data <= 14'h0008; 
        10'b0001001001: data <= 14'h0001; 
        10'b0001001010: data <= 14'h0004; 
        10'b0001001011: data <= 14'h000b; 
        10'b0001001100: data <= 14'h0009; 
        10'b0001001101: data <= 14'h000b; 
        10'b0001001110: data <= 14'h3ffb; 
        10'b0001001111: data <= 14'h0008; 
        10'b0001010000: data <= 14'h0003; 
        10'b0001010001: data <= 14'h0007; 
        10'b0001010010: data <= 14'h0006; 
        10'b0001010011: data <= 14'h000a; 
        10'b0001010100: data <= 14'h3fff; 
        10'b0001010101: data <= 14'h0001; 
        10'b0001010110: data <= 14'h000a; 
        10'b0001010111: data <= 14'h3ffe; 
        10'b0001011000: data <= 14'h0001; 
        10'b0001011001: data <= 14'h3fff; 
        10'b0001011010: data <= 14'h3ffc; 
        10'b0001011011: data <= 14'h0006; 
        10'b0001011100: data <= 14'h0000; 
        10'b0001011101: data <= 14'h0006; 
        10'b0001011110: data <= 14'h3ffb; 
        10'b0001011111: data <= 14'h0001; 
        10'b0001100000: data <= 14'h0005; 
        10'b0001100001: data <= 14'h3ff9; 
        10'b0001100010: data <= 14'h0006; 
        10'b0001100011: data <= 14'h3ffb; 
        10'b0001100100: data <= 14'h3ff6; 
        10'b0001100101: data <= 14'h3ff7; 
        10'b0001100110: data <= 14'h3ff9; 
        10'b0001100111: data <= 14'h3ffb; 
        10'b0001101000: data <= 14'h3fff; 
        10'b0001101001: data <= 14'h3ffb; 
        10'b0001101010: data <= 14'h0004; 
        10'b0001101011: data <= 14'h3fff; 
        10'b0001101100: data <= 14'h0005; 
        10'b0001101101: data <= 14'h000c; 
        10'b0001101110: data <= 14'h3ffc; 
        10'b0001101111: data <= 14'h0005; 
        10'b0001110000: data <= 14'h000c; 
        10'b0001110001: data <= 14'h3ffc; 
        10'b0001110010: data <= 14'h0007; 
        10'b0001110011: data <= 14'h3ffb; 
        10'b0001110100: data <= 14'h0003; 
        10'b0001110101: data <= 14'h3ffe; 
        10'b0001110110: data <= 14'h0001; 
        10'b0001110111: data <= 14'h3ffb; 
        10'b0001111000: data <= 14'h0004; 
        10'b0001111001: data <= 14'h3ffe; 
        10'b0001111010: data <= 14'h3ff4; 
        10'b0001111011: data <= 14'h3fea; 
        10'b0001111100: data <= 14'h3fe9; 
        10'b0001111101: data <= 14'h3fea; 
        10'b0001111110: data <= 14'h3fe5; 
        10'b0001111111: data <= 14'h3fd4; 
        10'b0010000000: data <= 14'h3fe6; 
        10'b0010000001: data <= 14'h3fec; 
        10'b0010000010: data <= 14'h3fef; 
        10'b0010000011: data <= 14'h3ffb; 
        10'b0010000100: data <= 14'h3ff3; 
        10'b0010000101: data <= 14'h0006; 
        10'b0010000110: data <= 14'h0001; 
        10'b0010000111: data <= 14'h3ffa; 
        10'b0010001000: data <= 14'h000b; 
        10'b0010001001: data <= 14'h0000; 
        10'b0010001010: data <= 14'h000b; 
        10'b0010001011: data <= 14'h000b; 
        10'b0010001100: data <= 14'h000a; 
        10'b0010001101: data <= 14'h0000; 
        10'b0010001110: data <= 14'h000a; 
        10'b0010001111: data <= 14'h3ffd; 
        10'b0010010000: data <= 14'h3ff8; 
        10'b0010010001: data <= 14'h3fff; 
        10'b0010010010: data <= 14'h3ffa; 
        10'b0010010011: data <= 14'h3ffe; 
        10'b0010010100: data <= 14'h3ff9; 
        10'b0010010101: data <= 14'h3ff0; 
        10'b0010010110: data <= 14'h3fd9; 
        10'b0010010111: data <= 14'h3fd0; 
        10'b0010011000: data <= 14'h3fc3; 
        10'b0010011001: data <= 14'h3fb9; 
        10'b0010011010: data <= 14'h3fa7; 
        10'b0010011011: data <= 14'h3fa8; 
        10'b0010011100: data <= 14'h3fa4; 
        10'b0010011101: data <= 14'h3fae; 
        10'b0010011110: data <= 14'h3fbb; 
        10'b0010011111: data <= 14'h3fcb; 
        10'b0010100000: data <= 14'h3fdb; 
        10'b0010100001: data <= 14'h3ff3; 
        10'b0010100010: data <= 14'h3feb; 
        10'b0010100011: data <= 14'h3ffd; 
        10'b0010100100: data <= 14'h0009; 
        10'b0010100101: data <= 14'h0007; 
        10'b0010100110: data <= 14'h3ffe; 
        10'b0010100111: data <= 14'h0000; 
        10'b0010101000: data <= 14'h0008; 
        10'b0010101001: data <= 14'h000b; 
        10'b0010101010: data <= 14'h0001; 
        10'b0010101011: data <= 14'h0002; 
        10'b0010101100: data <= 14'h000c; 
        10'b0010101101: data <= 14'h000f; 
        10'b0010101110: data <= 14'h0011; 
        10'b0010101111: data <= 14'h001a; 
        10'b0010110000: data <= 14'h0027; 
        10'b0010110001: data <= 14'h001f; 
        10'b0010110010: data <= 14'h0021; 
        10'b0010110011: data <= 14'h0006; 
        10'b0010110100: data <= 14'h3fe6; 
        10'b0010110101: data <= 14'h3fc9; 
        10'b0010110110: data <= 14'h3fc6; 
        10'b0010110111: data <= 14'h3fe2; 
        10'b0010111000: data <= 14'h3fee; 
        10'b0010111001: data <= 14'h3fea; 
        10'b0010111010: data <= 14'h3fe6; 
        10'b0010111011: data <= 14'h3fe2; 
        10'b0010111100: data <= 14'h3fd2; 
        10'b0010111101: data <= 14'h3fef; 
        10'b0010111110: data <= 14'h3fe0; 
        10'b0010111111: data <= 14'h3fe9; 
        10'b0011000000: data <= 14'h3ff0; 
        10'b0011000001: data <= 14'h3ffb; 
        10'b0011000010: data <= 14'h3ffb; 
        10'b0011000011: data <= 14'h0001; 
        10'b0011000100: data <= 14'h0008; 
        10'b0011000101: data <= 14'h000c; 
        10'b0011000110: data <= 14'h000a; 
        10'b0011000111: data <= 14'h0017; 
        10'b0011001000: data <= 14'h001b; 
        10'b0011001001: data <= 14'h0019; 
        10'b0011001010: data <= 14'h0024; 
        10'b0011001011: data <= 14'h0036; 
        10'b0011001100: data <= 14'h004a; 
        10'b0011001101: data <= 14'h003b; 
        10'b0011001110: data <= 14'h0029; 
        10'b0011001111: data <= 14'h002d; 
        10'b0011010000: data <= 14'h0030; 
        10'b0011010001: data <= 14'h0009; 
        10'b0011010010: data <= 14'h0007; 
        10'b0011010011: data <= 14'h0011; 
        10'b0011010100: data <= 14'h0032; 
        10'b0011010101: data <= 14'h0038; 
        10'b0011010110: data <= 14'h0026; 
        10'b0011010111: data <= 14'h001e; 
        10'b0011011000: data <= 14'h0007; 
        10'b0011011001: data <= 14'h3ff8; 
        10'b0011011010: data <= 14'h0004; 
        10'b0011011011: data <= 14'h3ff7; 
        10'b0011011100: data <= 14'h3ff8; 
        10'b0011011101: data <= 14'h0000; 
        10'b0011011110: data <= 14'h0006; 
        10'b0011011111: data <= 14'h3ffe; 
        10'b0011100000: data <= 14'h3ffa; 
        10'b0011100001: data <= 14'h000c; 
        10'b0011100010: data <= 14'h0005; 
        10'b0011100011: data <= 14'h0013; 
        10'b0011100100: data <= 14'h0026; 
        10'b0011100101: data <= 14'h0023; 
        10'b0011100110: data <= 14'h002e; 
        10'b0011100111: data <= 14'h0053; 
        10'b0011101000: data <= 14'h0038; 
        10'b0011101001: data <= 14'h0027; 
        10'b0011101010: data <= 14'h0031; 
        10'b0011101011: data <= 14'h0042; 
        10'b0011101100: data <= 14'h003f; 
        10'b0011101101: data <= 14'h0020; 
        10'b0011101110: data <= 14'h0012; 
        10'b0011101111: data <= 14'h001a; 
        10'b0011110000: data <= 14'h002c; 
        10'b0011110001: data <= 14'h0044; 
        10'b0011110010: data <= 14'h002f; 
        10'b0011110011: data <= 14'h0028; 
        10'b0011110100: data <= 14'h0020; 
        10'b0011110101: data <= 14'h0001; 
        10'b0011110110: data <= 14'h0013; 
        10'b0011110111: data <= 14'h0010; 
        10'b0011111000: data <= 14'h3ff4; 
        10'b0011111001: data <= 14'h3ffa; 
        10'b0011111010: data <= 14'h0006; 
        10'b0011111011: data <= 14'h000a; 
        10'b0011111100: data <= 14'h0005; 
        10'b0011111101: data <= 14'h000a; 
        10'b0011111110: data <= 14'h000d; 
        10'b0011111111: data <= 14'h001b; 
        10'b0100000000: data <= 14'h0026; 
        10'b0100000001: data <= 14'h002b; 
        10'b0100000010: data <= 14'h0010; 
        10'b0100000011: data <= 14'h0015; 
        10'b0100000100: data <= 14'h0018; 
        10'b0100000101: data <= 14'h0010; 
        10'b0100000110: data <= 14'h0026; 
        10'b0100000111: data <= 14'h002f; 
        10'b0100001000: data <= 14'h003c; 
        10'b0100001001: data <= 14'h0031; 
        10'b0100001010: data <= 14'h0046; 
        10'b0100001011: data <= 14'h0056; 
        10'b0100001100: data <= 14'h004f; 
        10'b0100001101: data <= 14'h0058; 
        10'b0100001110: data <= 14'h003a; 
        10'b0100001111: data <= 14'h003b; 
        10'b0100010000: data <= 14'h0031; 
        10'b0100010001: data <= 14'h0029; 
        10'b0100010010: data <= 14'h0014; 
        10'b0100010011: data <= 14'h3ff9; 
        10'b0100010100: data <= 14'h3ff4; 
        10'b0100010101: data <= 14'h3ffa; 
        10'b0100010110: data <= 14'h0005; 
        10'b0100010111: data <= 14'h3ffd; 
        10'b0100011000: data <= 14'h0002; 
        10'b0100011001: data <= 14'h000b; 
        10'b0100011010: data <= 14'h000c; 
        10'b0100011011: data <= 14'h0022; 
        10'b0100011100: data <= 14'h0027; 
        10'b0100011101: data <= 14'h0020; 
        10'b0100011110: data <= 14'h0006; 
        10'b0100011111: data <= 14'h000a; 
        10'b0100100000: data <= 14'h3ff3; 
        10'b0100100001: data <= 14'h0000; 
        10'b0100100010: data <= 14'h0018; 
        10'b0100100011: data <= 14'h002a; 
        10'b0100100100: data <= 14'h001d; 
        10'b0100100101: data <= 14'h0044; 
        10'b0100100110: data <= 14'h0057; 
        10'b0100100111: data <= 14'h006b; 
        10'b0100101000: data <= 14'h007a; 
        10'b0100101001: data <= 14'h005b; 
        10'b0100101010: data <= 14'h0047; 
        10'b0100101011: data <= 14'h004a; 
        10'b0100101100: data <= 14'h0041; 
        10'b0100101101: data <= 14'h0037; 
        10'b0100101110: data <= 14'h0018; 
        10'b0100101111: data <= 14'h3ff6; 
        10'b0100110000: data <= 14'h3fef; 
        10'b0100110001: data <= 14'h3ff9; 
        10'b0100110010: data <= 14'h0001; 
        10'b0100110011: data <= 14'h3ffd; 
        10'b0100110100: data <= 14'h0009; 
        10'b0100110101: data <= 14'h0007; 
        10'b0100110110: data <= 14'h000c; 
        10'b0100110111: data <= 14'h0023; 
        10'b0100111000: data <= 14'h002a; 
        10'b0100111001: data <= 14'h0015; 
        10'b0100111010: data <= 14'h0008; 
        10'b0100111011: data <= 14'h0007; 
        10'b0100111100: data <= 14'h0002; 
        10'b0100111101: data <= 14'h0019; 
        10'b0100111110: data <= 14'h000d; 
        10'b0100111111: data <= 14'h0010; 
        10'b0101000000: data <= 14'h001b; 
        10'b0101000001: data <= 14'h001b; 
        10'b0101000010: data <= 14'h001c; 
        10'b0101000011: data <= 14'h0052; 
        10'b0101000100: data <= 14'h006b; 
        10'b0101000101: data <= 14'h0047; 
        10'b0101000110: data <= 14'h0048; 
        10'b0101000111: data <= 14'h0037; 
        10'b0101001000: data <= 14'h0036; 
        10'b0101001001: data <= 14'h0022; 
        10'b0101001010: data <= 14'h0018; 
        10'b0101001011: data <= 14'h3ff8; 
        10'b0101001100: data <= 14'h3fe7; 
        10'b0101001101: data <= 14'h3fff; 
        10'b0101001110: data <= 14'h0002; 
        10'b0101001111: data <= 14'h000b; 
        10'b0101010000: data <= 14'h0008; 
        10'b0101010001: data <= 14'h3fff; 
        10'b0101010010: data <= 14'h0006; 
        10'b0101010011: data <= 14'h0016; 
        10'b0101010100: data <= 14'h0019; 
        10'b0101010101: data <= 14'h0004; 
        10'b0101010110: data <= 14'h0006; 
        10'b0101010111: data <= 14'h0017; 
        10'b0101011000: data <= 14'h0010; 
        10'b0101011001: data <= 14'h3fff; 
        10'b0101011010: data <= 14'h3fed; 
        10'b0101011011: data <= 14'h3fcd; 
        10'b0101011100: data <= 14'h3f94; 
        10'b0101011101: data <= 14'h3f59; 
        10'b0101011110: data <= 14'h3f83; 
        10'b0101011111: data <= 14'h0003; 
        10'b0101100000: data <= 14'h0047; 
        10'b0101100001: data <= 14'h0040; 
        10'b0101100010: data <= 14'h0019; 
        10'b0101100011: data <= 14'h0009; 
        10'b0101100100: data <= 14'h0002; 
        10'b0101100101: data <= 14'h3ff7; 
        10'b0101100110: data <= 14'h3ff8; 
        10'b0101100111: data <= 14'h3ff1; 
        10'b0101101000: data <= 14'h3ff5; 
        10'b0101101001: data <= 14'h000a; 
        10'b0101101010: data <= 14'h0007; 
        10'b0101101011: data <= 14'h0000; 
        10'b0101101100: data <= 14'h0009; 
        10'b0101101101: data <= 14'h0005; 
        10'b0101101110: data <= 14'h000a; 
        10'b0101101111: data <= 14'h0014; 
        10'b0101110000: data <= 14'h0007; 
        10'b0101110001: data <= 14'h0003; 
        10'b0101110010: data <= 14'h3ff9; 
        10'b0101110011: data <= 14'h0004; 
        10'b0101110100: data <= 14'h3ffd; 
        10'b0101110101: data <= 14'h3ff0; 
        10'b0101110110: data <= 14'h3fca; 
        10'b0101110111: data <= 14'h3f8f; 
        10'b0101111000: data <= 14'h3f39; 
        10'b0101111001: data <= 14'h3f22; 
        10'b0101111010: data <= 14'h3f89; 
        10'b0101111011: data <= 14'h3ff0; 
        10'b0101111100: data <= 14'h0024; 
        10'b0101111101: data <= 14'h0017; 
        10'b0101111110: data <= 14'h0005; 
        10'b0101111111: data <= 14'h000b; 
        10'b0110000000: data <= 14'h3fea; 
        10'b0110000001: data <= 14'h3fe4; 
        10'b0110000010: data <= 14'h3ff9; 
        10'b0110000011: data <= 14'h0002; 
        10'b0110000100: data <= 14'h3ffb; 
        10'b0110000101: data <= 14'h3ffc; 
        10'b0110000110: data <= 14'h0006; 
        10'b0110000111: data <= 14'h3ffb; 
        10'b0110001000: data <= 14'h3ffe; 
        10'b0110001001: data <= 14'h0005; 
        10'b0110001010: data <= 14'h0012; 
        10'b0110001011: data <= 14'h0016; 
        10'b0110001100: data <= 14'h000e; 
        10'b0110001101: data <= 14'h0010; 
        10'b0110001110: data <= 14'h3ffb; 
        10'b0110001111: data <= 14'h3ff5; 
        10'b0110010000: data <= 14'h3fe7; 
        10'b0110010001: data <= 14'h3fc5; 
        10'b0110010010: data <= 14'h3fa9; 
        10'b0110010011: data <= 14'h3f7a; 
        10'b0110010100: data <= 14'h3f54; 
        10'b0110010101: data <= 14'h3f6f; 
        10'b0110010110: data <= 14'h3fcb; 
        10'b0110010111: data <= 14'h0001; 
        10'b0110011000: data <= 14'h000b; 
        10'b0110011001: data <= 14'h0017; 
        10'b0110011010: data <= 14'h0042; 
        10'b0110011011: data <= 14'h0047; 
        10'b0110011100: data <= 14'h002a; 
        10'b0110011101: data <= 14'h001b; 
        10'b0110011110: data <= 14'h001b; 
        10'b0110011111: data <= 14'h0018; 
        10'b0110100000: data <= 14'h0008; 
        10'b0110100001: data <= 14'h0002; 
        10'b0110100010: data <= 14'h3ffc; 
        10'b0110100011: data <= 14'h3ffd; 
        10'b0110100100: data <= 14'h0006; 
        10'b0110100101: data <= 14'h0008; 
        10'b0110100110: data <= 14'h0003; 
        10'b0110100111: data <= 14'h0008; 
        10'b0110101000: data <= 14'h0008; 
        10'b0110101001: data <= 14'h3fe8; 
        10'b0110101010: data <= 14'h3ff5; 
        10'b0110101011: data <= 14'h3ff1; 
        10'b0110101100: data <= 14'h3fc1; 
        10'b0110101101: data <= 14'h3fb3; 
        10'b0110101110: data <= 14'h3f9a; 
        10'b0110101111: data <= 14'h3f8b; 
        10'b0110110000: data <= 14'h3f81; 
        10'b0110110001: data <= 14'h3fa2; 
        10'b0110110010: data <= 14'h3fc9; 
        10'b0110110011: data <= 14'h0002; 
        10'b0110110100: data <= 14'h0006; 
        10'b0110110101: data <= 14'h0059; 
        10'b0110110110: data <= 14'h0069; 
        10'b0110110111: data <= 14'h0056; 
        10'b0110111000: data <= 14'h004d; 
        10'b0110111001: data <= 14'h0042; 
        10'b0110111010: data <= 14'h002b; 
        10'b0110111011: data <= 14'h0013; 
        10'b0110111100: data <= 14'h3fff; 
        10'b0110111101: data <= 14'h3ffb; 
        10'b0110111110: data <= 14'h0001; 
        10'b0110111111: data <= 14'h0009; 
        10'b0111000000: data <= 14'h0006; 
        10'b0111000001: data <= 14'h000b; 
        10'b0111000010: data <= 14'h3fff; 
        10'b0111000011: data <= 14'h000c; 
        10'b0111000100: data <= 14'h0009; 
        10'b0111000101: data <= 14'h3ff5; 
        10'b0111000110: data <= 14'h3ff1; 
        10'b0111000111: data <= 14'h3ffe; 
        10'b0111001000: data <= 14'h3fcd; 
        10'b0111001001: data <= 14'h3fc7; 
        10'b0111001010: data <= 14'h3fa3; 
        10'b0111001011: data <= 14'h3f92; 
        10'b0111001100: data <= 14'h3fbb; 
        10'b0111001101: data <= 14'h3fd9; 
        10'b0111001110: data <= 14'h3fc8; 
        10'b0111001111: data <= 14'h001d; 
        10'b0111010000: data <= 14'h0023; 
        10'b0111010001: data <= 14'h004c; 
        10'b0111010010: data <= 14'h0041; 
        10'b0111010011: data <= 14'h0044; 
        10'b0111010100: data <= 14'h0036; 
        10'b0111010101: data <= 14'h0029; 
        10'b0111010110: data <= 14'h0008; 
        10'b0111010111: data <= 14'h3fef; 
        10'b0111011000: data <= 14'h3ff6; 
        10'b0111011001: data <= 14'h3ffa; 
        10'b0111011010: data <= 14'h0006; 
        10'b0111011011: data <= 14'h000b; 
        10'b0111011100: data <= 14'h0000; 
        10'b0111011101: data <= 14'h0001; 
        10'b0111011110: data <= 14'h0007; 
        10'b0111011111: data <= 14'h0000; 
        10'b0111100000: data <= 14'h0002; 
        10'b0111100001: data <= 14'h3ff9; 
        10'b0111100010: data <= 14'h3fde; 
        10'b0111100011: data <= 14'h3fd3; 
        10'b0111100100: data <= 14'h3fc7; 
        10'b0111100101: data <= 14'h3fd1; 
        10'b0111100110: data <= 14'h3fc2; 
        10'b0111100111: data <= 14'h3fd2; 
        10'b0111101000: data <= 14'h3ff1; 
        10'b0111101001: data <= 14'h000b; 
        10'b0111101010: data <= 14'h0007; 
        10'b0111101011: data <= 14'h000b; 
        10'b0111101100: data <= 14'h3ff9; 
        10'b0111101101: data <= 14'h0012; 
        10'b0111101110: data <= 14'h0010; 
        10'b0111101111: data <= 14'h000c; 
        10'b0111110000: data <= 14'h0006; 
        10'b0111110001: data <= 14'h3ff7; 
        10'b0111110010: data <= 14'h3feb; 
        10'b0111110011: data <= 14'h3ff7; 
        10'b0111110100: data <= 14'h3ff8; 
        10'b0111110101: data <= 14'h3ffa; 
        10'b0111110110: data <= 14'h3ffd; 
        10'b0111110111: data <= 14'h3ffd; 
        10'b0111111000: data <= 14'h3ffd; 
        10'b0111111001: data <= 14'h3fff; 
        10'b0111111010: data <= 14'h0008; 
        10'b0111111011: data <= 14'h0002; 
        10'b0111111100: data <= 14'h3ff2; 
        10'b0111111101: data <= 14'h3fdf; 
        10'b0111111110: data <= 14'h3fc9; 
        10'b0111111111: data <= 14'h3fbc; 
        10'b1000000000: data <= 14'h3fc1; 
        10'b1000000001: data <= 14'h3fc5; 
        10'b1000000010: data <= 14'h3fb4; 
        10'b1000000011: data <= 14'h3fe6; 
        10'b1000000100: data <= 14'h3ff8; 
        10'b1000000101: data <= 14'h0001; 
        10'b1000000110: data <= 14'h0015; 
        10'b1000000111: data <= 14'h3fe9; 
        10'b1000001000: data <= 14'h3fe4; 
        10'b1000001001: data <= 14'h3ff1; 
        10'b1000001010: data <= 14'h3fdd; 
        10'b1000001011: data <= 14'h3feb; 
        10'b1000001100: data <= 14'h3fdc; 
        10'b1000001101: data <= 14'h3fc9; 
        10'b1000001110: data <= 14'h3fd8; 
        10'b1000001111: data <= 14'h3fe7; 
        10'b1000010000: data <= 14'h3fec; 
        10'b1000010001: data <= 14'h0002; 
        10'b1000010010: data <= 14'h3ffe; 
        10'b1000010011: data <= 14'h0000; 
        10'b1000010100: data <= 14'h000b; 
        10'b1000010101: data <= 14'h000c; 
        10'b1000010110: data <= 14'h000b; 
        10'b1000010111: data <= 14'h0005; 
        10'b1000011000: data <= 14'h3ff7; 
        10'b1000011001: data <= 14'h3fd5; 
        10'b1000011010: data <= 14'h3fbb; 
        10'b1000011011: data <= 14'h3fb6; 
        10'b1000011100: data <= 14'h3fb4; 
        10'b1000011101: data <= 14'h3fb4; 
        10'b1000011110: data <= 14'h3fcc; 
        10'b1000011111: data <= 14'h3fdb; 
        10'b1000100000: data <= 14'h3fea; 
        10'b1000100001: data <= 14'h000a; 
        10'b1000100010: data <= 14'h001e; 
        10'b1000100011: data <= 14'h3fe0; 
        10'b1000100100: data <= 14'h3fe1; 
        10'b1000100101: data <= 14'h3fd9; 
        10'b1000100110: data <= 14'h3fc2; 
        10'b1000100111: data <= 14'h3fc5; 
        10'b1000101000: data <= 14'h3fb8; 
        10'b1000101001: data <= 14'h3fbd; 
        10'b1000101010: data <= 14'h3fcd; 
        10'b1000101011: data <= 14'h3fdd; 
        10'b1000101100: data <= 14'h3fee; 
        10'b1000101101: data <= 14'h3ff9; 
        10'b1000101110: data <= 14'h000b; 
        10'b1000101111: data <= 14'h3ffb; 
        10'b1000110000: data <= 14'h3ffa; 
        10'b1000110001: data <= 14'h3ffd; 
        10'b1000110010: data <= 14'h0005; 
        10'b1000110011: data <= 14'h3ffe; 
        10'b1000110100: data <= 14'h3ff5; 
        10'b1000110101: data <= 14'h3fdf; 
        10'b1000110110: data <= 14'h3fbb; 
        10'b1000110111: data <= 14'h3fb8; 
        10'b1000111000: data <= 14'h3fbc; 
        10'b1000111001: data <= 14'h3fbd; 
        10'b1000111010: data <= 14'h3fd2; 
        10'b1000111011: data <= 14'h3fd0; 
        10'b1000111100: data <= 14'h0003; 
        10'b1000111101: data <= 14'h0005; 
        10'b1000111110: data <= 14'h0010; 
        10'b1000111111: data <= 14'h3fd6; 
        10'b1001000000: data <= 14'h3fcb; 
        10'b1001000001: data <= 14'h3fbb; 
        10'b1001000010: data <= 14'h3fa1; 
        10'b1001000011: data <= 14'h3fc3; 
        10'b1001000100: data <= 14'h3fac; 
        10'b1001000101: data <= 14'h3fc0; 
        10'b1001000110: data <= 14'h3fd2; 
        10'b1001000111: data <= 14'h3fec; 
        10'b1001001000: data <= 14'h3ff3; 
        10'b1001001001: data <= 14'h000a; 
        10'b1001001010: data <= 14'h0009; 
        10'b1001001011: data <= 14'h0006; 
        10'b1001001100: data <= 14'h0009; 
        10'b1001001101: data <= 14'h0009; 
        10'b1001001110: data <= 14'h0002; 
        10'b1001001111: data <= 14'h3ff4; 
        10'b1001010000: data <= 14'h3ffa; 
        10'b1001010001: data <= 14'h3fe2; 
        10'b1001010010: data <= 14'h3fdd; 
        10'b1001010011: data <= 14'h3fce; 
        10'b1001010100: data <= 14'h3fd3; 
        10'b1001010101: data <= 14'h3fe5; 
        10'b1001010110: data <= 14'h3fda; 
        10'b1001010111: data <= 14'h3fe1; 
        10'b1001011000: data <= 14'h3ff2; 
        10'b1001011001: data <= 14'h0002; 
        10'b1001011010: data <= 14'h3ff8; 
        10'b1001011011: data <= 14'h3fe3; 
        10'b1001011100: data <= 14'h3fdf; 
        10'b1001011101: data <= 14'h3fbc; 
        10'b1001011110: data <= 14'h3fbc; 
        10'b1001011111: data <= 14'h3fbc; 
        10'b1001100000: data <= 14'h3fb8; 
        10'b1001100001: data <= 14'h3fc3; 
        10'b1001100010: data <= 14'h3fdc; 
        10'b1001100011: data <= 14'h3fe5; 
        10'b1001100100: data <= 14'h3fff; 
        10'b1001100101: data <= 14'h0004; 
        10'b1001100110: data <= 14'h0009; 
        10'b1001100111: data <= 14'h3ffe; 
        10'b1001101000: data <= 14'h0003; 
        10'b1001101001: data <= 14'h0001; 
        10'b1001101010: data <= 14'h0002; 
        10'b1001101011: data <= 14'h3ff8; 
        10'b1001101100: data <= 14'h3ffd; 
        10'b1001101101: data <= 14'h0004; 
        10'b1001101110: data <= 14'h3ff5; 
        10'b1001101111: data <= 14'h0005; 
        10'b1001110000: data <= 14'h0009; 
        10'b1001110001: data <= 14'h3ff2; 
        10'b1001110010: data <= 14'h3fe6; 
        10'b1001110011: data <= 14'h3fd4; 
        10'b1001110100: data <= 14'h3fd6; 
        10'b1001110101: data <= 14'h3fef; 
        10'b1001110110: data <= 14'h0005; 
        10'b1001110111: data <= 14'h0005; 
        10'b1001111000: data <= 14'h3fe6; 
        10'b1001111001: data <= 14'h3fe0; 
        10'b1001111010: data <= 14'h3fc9; 
        10'b1001111011: data <= 14'h3fca; 
        10'b1001111100: data <= 14'h3fc3; 
        10'b1001111101: data <= 14'h3fca; 
        10'b1001111110: data <= 14'h3fe5; 
        10'b1001111111: data <= 14'h3ff7; 
        10'b1010000000: data <= 14'h0006; 
        10'b1010000001: data <= 14'h3ffa; 
        10'b1010000010: data <= 14'h0003; 
        10'b1010000011: data <= 14'h0000; 
        10'b1010000100: data <= 14'h0004; 
        10'b1010000101: data <= 14'h0008; 
        10'b1010000110: data <= 14'h3ff9; 
        10'b1010000111: data <= 14'h3ffa; 
        10'b1010001000: data <= 14'h000b; 
        10'b1010001001: data <= 14'h000f; 
        10'b1010001010: data <= 14'h0021; 
        10'b1010001011: data <= 14'h002c; 
        10'b1010001100: data <= 14'h0015; 
        10'b1010001101: data <= 14'h0004; 
        10'b1010001110: data <= 14'h3ff3; 
        10'b1010001111: data <= 14'h3fe2; 
        10'b1010010000: data <= 14'h3fe8; 
        10'b1010010001: data <= 14'h0002; 
        10'b1010010010: data <= 14'h0011; 
        10'b1010010011: data <= 14'h0010; 
        10'b1010010100: data <= 14'h3ff9; 
        10'b1010010101: data <= 14'h3ff6; 
        10'b1010010110: data <= 14'h3fdd; 
        10'b1010010111: data <= 14'h3fcf; 
        10'b1010011000: data <= 14'h3fce; 
        10'b1010011001: data <= 14'h3fd9; 
        10'b1010011010: data <= 14'h3fe0; 
        10'b1010011011: data <= 14'h3feb; 
        10'b1010011100: data <= 14'h3ff7; 
        10'b1010011101: data <= 14'h0001; 
        10'b1010011110: data <= 14'h0001; 
        10'b1010011111: data <= 14'h3ffd; 
        10'b1010100000: data <= 14'h0000; 
        10'b1010100001: data <= 14'h3fff; 
        10'b1010100010: data <= 14'h0003; 
        10'b1010100011: data <= 14'h0007; 
        10'b1010100100: data <= 14'h0010; 
        10'b1010100101: data <= 14'h0024; 
        10'b1010100110: data <= 14'h0036; 
        10'b1010100111: data <= 14'h003d; 
        10'b1010101000: data <= 14'h0034; 
        10'b1010101001: data <= 14'h001b; 
        10'b1010101010: data <= 14'h003a; 
        10'b1010101011: data <= 14'h0022; 
        10'b1010101100: data <= 14'h001e; 
        10'b1010101101: data <= 14'h002a; 
        10'b1010101110: data <= 14'h001a; 
        10'b1010101111: data <= 14'h0025; 
        10'b1010110000: data <= 14'h0016; 
        10'b1010110001: data <= 14'h0011; 
        10'b1010110010: data <= 14'h3fff; 
        10'b1010110011: data <= 14'h3ff0; 
        10'b1010110100: data <= 14'h3fef; 
        10'b1010110101: data <= 14'h3feb; 
        10'b1010110110: data <= 14'h3fe9; 
        10'b1010110111: data <= 14'h3feb; 
        10'b1010111000: data <= 14'h0003; 
        10'b1010111001: data <= 14'h3ffe; 
        10'b1010111010: data <= 14'h3ffa; 
        10'b1010111011: data <= 14'h0006; 
        10'b1010111100: data <= 14'h3ffa; 
        10'b1010111101: data <= 14'h0005; 
        10'b1010111110: data <= 14'h0009; 
        10'b1010111111: data <= 14'h0009; 
        10'b1011000000: data <= 14'h0005; 
        10'b1011000001: data <= 14'h0012; 
        10'b1011000010: data <= 14'h001b; 
        10'b1011000011: data <= 14'h0029; 
        10'b1011000100: data <= 14'h003f; 
        10'b1011000101: data <= 14'h003e; 
        10'b1011000110: data <= 14'h0049; 
        10'b1011000111: data <= 14'h0044; 
        10'b1011001000: data <= 14'h003d; 
        10'b1011001001: data <= 14'h0030; 
        10'b1011001010: data <= 14'h0031; 
        10'b1011001011: data <= 14'h0034; 
        10'b1011001100: data <= 14'h002c; 
        10'b1011001101: data <= 14'h0029; 
        10'b1011001110: data <= 14'h0021; 
        10'b1011001111: data <= 14'h000b; 
        10'b1011010000: data <= 14'h3ff2; 
        10'b1011010001: data <= 14'h0002; 
        10'b1011010010: data <= 14'h3ff9; 
        10'b1011010011: data <= 14'h3ffb; 
        10'b1011010100: data <= 14'h3ffe; 
        10'b1011010101: data <= 14'h0003; 
        10'b1011010110: data <= 14'h000c; 
        10'b1011010111: data <= 14'h0008; 
        10'b1011011000: data <= 14'h3ffc; 
        10'b1011011001: data <= 14'h0002; 
        10'b1011011010: data <= 14'h000c; 
        10'b1011011011: data <= 14'h3ffe; 
        10'b1011011100: data <= 14'h3ffc; 
        10'b1011011101: data <= 14'h000b; 
        10'b1011011110: data <= 14'h0001; 
        10'b1011011111: data <= 14'h000a; 
        10'b1011100000: data <= 14'h000a; 
        10'b1011100001: data <= 14'h0001; 
        10'b1011100010: data <= 14'h000e; 
        10'b1011100011: data <= 14'h0014; 
        10'b1011100100: data <= 14'h0006; 
        10'b1011100101: data <= 14'h0011; 
        10'b1011100110: data <= 14'h0025; 
        10'b1011100111: data <= 14'h002e; 
        10'b1011101000: data <= 14'h0024; 
        10'b1011101001: data <= 14'h002f; 
        10'b1011101010: data <= 14'h001b; 
        10'b1011101011: data <= 14'h000d; 
        10'b1011101100: data <= 14'h0000; 
        10'b1011101101: data <= 14'h0005; 
        10'b1011101110: data <= 14'h3fff; 
        10'b1011101111: data <= 14'h0003; 
        10'b1011110000: data <= 14'h0001; 
        10'b1011110001: data <= 14'h3ffd; 
        10'b1011110010: data <= 14'h3fff; 
        10'b1011110011: data <= 14'h3ffe; 
        10'b1011110100: data <= 14'h3ffa; 
        10'b1011110101: data <= 14'h0005; 
        10'b1011110110: data <= 14'h0003; 
        10'b1011110111: data <= 14'h0006; 
        10'b1011111000: data <= 14'h0008; 
        10'b1011111001: data <= 14'h0005; 
        10'b1011111010: data <= 14'h0002; 
        10'b1011111011: data <= 14'h0001; 
        10'b1011111100: data <= 14'h000d; 
        10'b1011111101: data <= 14'h0008; 
        10'b1011111110: data <= 14'h0002; 
        10'b1011111111: data <= 14'h0008; 
        10'b1100000000: data <= 14'h0004; 
        10'b1100000001: data <= 14'h000f; 
        10'b1100000010: data <= 14'h0009; 
        10'b1100000011: data <= 14'h0007; 
        10'b1100000100: data <= 14'h0015; 
        10'b1100000101: data <= 14'h0007; 
        10'b1100000110: data <= 14'h0006; 
        10'b1100000111: data <= 14'h000f; 
        10'b1100001000: data <= 14'h0002; 
        10'b1100001001: data <= 14'h3ffe; 
        10'b1100001010: data <= 14'h000c; 
        10'b1100001011: data <= 14'h0007; 
        10'b1100001100: data <= 14'h0003; 
        10'b1100001101: data <= 14'h3ffe; 
        10'b1100001110: data <= 14'h3ffb; 
        10'b1100001111: data <= 14'h0008; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 9) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 15'h0002; 
        10'b0000000001: data <= 15'h0002; 
        10'b0000000010: data <= 15'h000f; 
        10'b0000000011: data <= 15'h0006; 
        10'b0000000100: data <= 15'h0019; 
        10'b0000000101: data <= 15'h7ff5; 
        10'b0000000110: data <= 15'h7ff9; 
        10'b0000000111: data <= 15'h0008; 
        10'b0000001000: data <= 15'h0013; 
        10'b0000001001: data <= 15'h0013; 
        10'b0000001010: data <= 15'h7ff5; 
        10'b0000001011: data <= 15'h0005; 
        10'b0000001100: data <= 15'h0005; 
        10'b0000001101: data <= 15'h7ffd; 
        10'b0000001110: data <= 15'h0014; 
        10'b0000001111: data <= 15'h0005; 
        10'b0000010000: data <= 15'h0000; 
        10'b0000010001: data <= 15'h7fff; 
        10'b0000010010: data <= 15'h0002; 
        10'b0000010011: data <= 15'h0007; 
        10'b0000010100: data <= 15'h000d; 
        10'b0000010101: data <= 15'h0018; 
        10'b0000010110: data <= 15'h7ffa; 
        10'b0000010111: data <= 15'h0012; 
        10'b0000011000: data <= 15'h7ffe; 
        10'b0000011001: data <= 15'h000d; 
        10'b0000011010: data <= 15'h7fff; 
        10'b0000011011: data <= 15'h0000; 
        10'b0000011100: data <= 15'h0017; 
        10'b0000011101: data <= 15'h7ffb; 
        10'b0000011110: data <= 15'h0005; 
        10'b0000011111: data <= 15'h0016; 
        10'b0000100000: data <= 15'h0009; 
        10'b0000100001: data <= 15'h0001; 
        10'b0000100010: data <= 15'h0016; 
        10'b0000100011: data <= 15'h0007; 
        10'b0000100100: data <= 15'h0002; 
        10'b0000100101: data <= 15'h7ffc; 
        10'b0000100110: data <= 15'h7ffd; 
        10'b0000100111: data <= 15'h7ff4; 
        10'b0000101000: data <= 15'h0013; 
        10'b0000101001: data <= 15'h7fff; 
        10'b0000101010: data <= 15'h0017; 
        10'b0000101011: data <= 15'h7ffa; 
        10'b0000101100: data <= 15'h000a; 
        10'b0000101101: data <= 15'h0011; 
        10'b0000101110: data <= 15'h0013; 
        10'b0000101111: data <= 15'h0010; 
        10'b0000110000: data <= 15'h0001; 
        10'b0000110001: data <= 15'h000f; 
        10'b0000110010: data <= 15'h0000; 
        10'b0000110011: data <= 15'h0018; 
        10'b0000110100: data <= 15'h0013; 
        10'b0000110101: data <= 15'h7ff9; 
        10'b0000110110: data <= 15'h7ff9; 
        10'b0000110111: data <= 15'h000a; 
        10'b0000111000: data <= 15'h0016; 
        10'b0000111001: data <= 15'h0015; 
        10'b0000111010: data <= 15'h0011; 
        10'b0000111011: data <= 15'h7ffd; 
        10'b0000111100: data <= 15'h0013; 
        10'b0000111101: data <= 15'h7ff7; 
        10'b0000111110: data <= 15'h7ff8; 
        10'b0000111111: data <= 15'h000f; 
        10'b0001000000: data <= 15'h000d; 
        10'b0001000001: data <= 15'h7ff8; 
        10'b0001000010: data <= 15'h7ffe; 
        10'b0001000011: data <= 15'h0009; 
        10'b0001000100: data <= 15'h7ffd; 
        10'b0001000101: data <= 15'h7ffb; 
        10'b0001000110: data <= 15'h0006; 
        10'b0001000111: data <= 15'h0014; 
        10'b0001001000: data <= 15'h0010; 
        10'b0001001001: data <= 15'h0003; 
        10'b0001001010: data <= 15'h0008; 
        10'b0001001011: data <= 15'h0016; 
        10'b0001001100: data <= 15'h0013; 
        10'b0001001101: data <= 15'h0016; 
        10'b0001001110: data <= 15'h7ff5; 
        10'b0001001111: data <= 15'h0011; 
        10'b0001010000: data <= 15'h0006; 
        10'b0001010001: data <= 15'h000f; 
        10'b0001010010: data <= 15'h000d; 
        10'b0001010011: data <= 15'h0013; 
        10'b0001010100: data <= 15'h7ffe; 
        10'b0001010101: data <= 15'h0001; 
        10'b0001010110: data <= 15'h0014; 
        10'b0001010111: data <= 15'h7ffd; 
        10'b0001011000: data <= 15'h0002; 
        10'b0001011001: data <= 15'h7fff; 
        10'b0001011010: data <= 15'h7ff9; 
        10'b0001011011: data <= 15'h000d; 
        10'b0001011100: data <= 15'h0000; 
        10'b0001011101: data <= 15'h000d; 
        10'b0001011110: data <= 15'h7ff5; 
        10'b0001011111: data <= 15'h0003; 
        10'b0001100000: data <= 15'h000a; 
        10'b0001100001: data <= 15'h7ff2; 
        10'b0001100010: data <= 15'h000c; 
        10'b0001100011: data <= 15'h7ff6; 
        10'b0001100100: data <= 15'h7feb; 
        10'b0001100101: data <= 15'h7fef; 
        10'b0001100110: data <= 15'h7ff1; 
        10'b0001100111: data <= 15'h7ff6; 
        10'b0001101000: data <= 15'h7ffe; 
        10'b0001101001: data <= 15'h7ff7; 
        10'b0001101010: data <= 15'h0008; 
        10'b0001101011: data <= 15'h7fff; 
        10'b0001101100: data <= 15'h000a; 
        10'b0001101101: data <= 15'h0018; 
        10'b0001101110: data <= 15'h7ff8; 
        10'b0001101111: data <= 15'h000a; 
        10'b0001110000: data <= 15'h0018; 
        10'b0001110001: data <= 15'h7ff7; 
        10'b0001110010: data <= 15'h000d; 
        10'b0001110011: data <= 15'h7ff6; 
        10'b0001110100: data <= 15'h0006; 
        10'b0001110101: data <= 15'h7ffb; 
        10'b0001110110: data <= 15'h0001; 
        10'b0001110111: data <= 15'h7ff6; 
        10'b0001111000: data <= 15'h0007; 
        10'b0001111001: data <= 15'h7ffd; 
        10'b0001111010: data <= 15'h7fe9; 
        10'b0001111011: data <= 15'h7fd3; 
        10'b0001111100: data <= 15'h7fd1; 
        10'b0001111101: data <= 15'h7fd3; 
        10'b0001111110: data <= 15'h7fcb; 
        10'b0001111111: data <= 15'h7fa8; 
        10'b0010000000: data <= 15'h7fcc; 
        10'b0010000001: data <= 15'h7fd9; 
        10'b0010000010: data <= 15'h7fde; 
        10'b0010000011: data <= 15'h7ff7; 
        10'b0010000100: data <= 15'h7fe7; 
        10'b0010000101: data <= 15'h000c; 
        10'b0010000110: data <= 15'h0002; 
        10'b0010000111: data <= 15'h7ff4; 
        10'b0010001000: data <= 15'h0016; 
        10'b0010001001: data <= 15'h7fff; 
        10'b0010001010: data <= 15'h0016; 
        10'b0010001011: data <= 15'h0015; 
        10'b0010001100: data <= 15'h0014; 
        10'b0010001101: data <= 15'h0001; 
        10'b0010001110: data <= 15'h0013; 
        10'b0010001111: data <= 15'h7ffb; 
        10'b0010010000: data <= 15'h7ff1; 
        10'b0010010001: data <= 15'h7ffd; 
        10'b0010010010: data <= 15'h7ff4; 
        10'b0010010011: data <= 15'h7ffc; 
        10'b0010010100: data <= 15'h7ff2; 
        10'b0010010101: data <= 15'h7fe0; 
        10'b0010010110: data <= 15'h7fb1; 
        10'b0010010111: data <= 15'h7f9f; 
        10'b0010011000: data <= 15'h7f86; 
        10'b0010011001: data <= 15'h7f72; 
        10'b0010011010: data <= 15'h7f4e; 
        10'b0010011011: data <= 15'h7f50; 
        10'b0010011100: data <= 15'h7f47; 
        10'b0010011101: data <= 15'h7f5d; 
        10'b0010011110: data <= 15'h7f76; 
        10'b0010011111: data <= 15'h7f97; 
        10'b0010100000: data <= 15'h7fb5; 
        10'b0010100001: data <= 15'h7fe5; 
        10'b0010100010: data <= 15'h7fd7; 
        10'b0010100011: data <= 15'h7ffb; 
        10'b0010100100: data <= 15'h0012; 
        10'b0010100101: data <= 15'h000e; 
        10'b0010100110: data <= 15'h7ffc; 
        10'b0010100111: data <= 15'h0001; 
        10'b0010101000: data <= 15'h0011; 
        10'b0010101001: data <= 15'h0017; 
        10'b0010101010: data <= 15'h0002; 
        10'b0010101011: data <= 15'h0004; 
        10'b0010101100: data <= 15'h0019; 
        10'b0010101101: data <= 15'h001e; 
        10'b0010101110: data <= 15'h0023; 
        10'b0010101111: data <= 15'h0034; 
        10'b0010110000: data <= 15'h004d; 
        10'b0010110001: data <= 15'h003e; 
        10'b0010110010: data <= 15'h0042; 
        10'b0010110011: data <= 15'h000c; 
        10'b0010110100: data <= 15'h7fcb; 
        10'b0010110101: data <= 15'h7f91; 
        10'b0010110110: data <= 15'h7f8c; 
        10'b0010110111: data <= 15'h7fc4; 
        10'b0010111000: data <= 15'h7fdc; 
        10'b0010111001: data <= 15'h7fd5; 
        10'b0010111010: data <= 15'h7fcb; 
        10'b0010111011: data <= 15'h7fc3; 
        10'b0010111100: data <= 15'h7fa4; 
        10'b0010111101: data <= 15'h7fdd; 
        10'b0010111110: data <= 15'h7fc0; 
        10'b0010111111: data <= 15'h7fd1; 
        10'b0011000000: data <= 15'h7fe1; 
        10'b0011000001: data <= 15'h7ff5; 
        10'b0011000010: data <= 15'h7ff5; 
        10'b0011000011: data <= 15'h0003; 
        10'b0011000100: data <= 15'h000f; 
        10'b0011000101: data <= 15'h0017; 
        10'b0011000110: data <= 15'h0013; 
        10'b0011000111: data <= 15'h002d; 
        10'b0011001000: data <= 15'h0037; 
        10'b0011001001: data <= 15'h0031; 
        10'b0011001010: data <= 15'h0047; 
        10'b0011001011: data <= 15'h006d; 
        10'b0011001100: data <= 15'h0095; 
        10'b0011001101: data <= 15'h0076; 
        10'b0011001110: data <= 15'h0051; 
        10'b0011001111: data <= 15'h005a; 
        10'b0011010000: data <= 15'h005f; 
        10'b0011010001: data <= 15'h0012; 
        10'b0011010010: data <= 15'h000e; 
        10'b0011010011: data <= 15'h0022; 
        10'b0011010100: data <= 15'h0065; 
        10'b0011010101: data <= 15'h0070; 
        10'b0011010110: data <= 15'h004c; 
        10'b0011010111: data <= 15'h003d; 
        10'b0011011000: data <= 15'h000f; 
        10'b0011011001: data <= 15'h7fef; 
        10'b0011011010: data <= 15'h0008; 
        10'b0011011011: data <= 15'h7fee; 
        10'b0011011100: data <= 15'h7fef; 
        10'b0011011101: data <= 15'h7fff; 
        10'b0011011110: data <= 15'h000c; 
        10'b0011011111: data <= 15'h7ffb; 
        10'b0011100000: data <= 15'h7ff4; 
        10'b0011100001: data <= 15'h0018; 
        10'b0011100010: data <= 15'h0009; 
        10'b0011100011: data <= 15'h0026; 
        10'b0011100100: data <= 15'h004d; 
        10'b0011100101: data <= 15'h0045; 
        10'b0011100110: data <= 15'h005d; 
        10'b0011100111: data <= 15'h00a7; 
        10'b0011101000: data <= 15'h0070; 
        10'b0011101001: data <= 15'h004d; 
        10'b0011101010: data <= 15'h0062; 
        10'b0011101011: data <= 15'h0084; 
        10'b0011101100: data <= 15'h007d; 
        10'b0011101101: data <= 15'h003f; 
        10'b0011101110: data <= 15'h0025; 
        10'b0011101111: data <= 15'h0033; 
        10'b0011110000: data <= 15'h0059; 
        10'b0011110001: data <= 15'h0089; 
        10'b0011110010: data <= 15'h005e; 
        10'b0011110011: data <= 15'h0050; 
        10'b0011110100: data <= 15'h0040; 
        10'b0011110101: data <= 15'h0001; 
        10'b0011110110: data <= 15'h0027; 
        10'b0011110111: data <= 15'h0021; 
        10'b0011111000: data <= 15'h7fe9; 
        10'b0011111001: data <= 15'h7ff5; 
        10'b0011111010: data <= 15'h000d; 
        10'b0011111011: data <= 15'h0014; 
        10'b0011111100: data <= 15'h000a; 
        10'b0011111101: data <= 15'h0013; 
        10'b0011111110: data <= 15'h001a; 
        10'b0011111111: data <= 15'h0037; 
        10'b0100000000: data <= 15'h004b; 
        10'b0100000001: data <= 15'h0056; 
        10'b0100000010: data <= 15'h001f; 
        10'b0100000011: data <= 15'h002a; 
        10'b0100000100: data <= 15'h002f; 
        10'b0100000101: data <= 15'h001f; 
        10'b0100000110: data <= 15'h004d; 
        10'b0100000111: data <= 15'h005e; 
        10'b0100001000: data <= 15'h0078; 
        10'b0100001001: data <= 15'h0062; 
        10'b0100001010: data <= 15'h008c; 
        10'b0100001011: data <= 15'h00ac; 
        10'b0100001100: data <= 15'h009f; 
        10'b0100001101: data <= 15'h00b1; 
        10'b0100001110: data <= 15'h0074; 
        10'b0100001111: data <= 15'h0076; 
        10'b0100010000: data <= 15'h0063; 
        10'b0100010001: data <= 15'h0053; 
        10'b0100010010: data <= 15'h0027; 
        10'b0100010011: data <= 15'h7ff2; 
        10'b0100010100: data <= 15'h7fe8; 
        10'b0100010101: data <= 15'h7ff4; 
        10'b0100010110: data <= 15'h000a; 
        10'b0100010111: data <= 15'h7ffb; 
        10'b0100011000: data <= 15'h0004; 
        10'b0100011001: data <= 15'h0015; 
        10'b0100011010: data <= 15'h0017; 
        10'b0100011011: data <= 15'h0044; 
        10'b0100011100: data <= 15'h004e; 
        10'b0100011101: data <= 15'h0041; 
        10'b0100011110: data <= 15'h000c; 
        10'b0100011111: data <= 15'h0014; 
        10'b0100100000: data <= 15'h7fe6; 
        10'b0100100001: data <= 15'h7fff; 
        10'b0100100010: data <= 15'h0030; 
        10'b0100100011: data <= 15'h0054; 
        10'b0100100100: data <= 15'h003a; 
        10'b0100100101: data <= 15'h0088; 
        10'b0100100110: data <= 15'h00af; 
        10'b0100100111: data <= 15'h00d7; 
        10'b0100101000: data <= 15'h00f4; 
        10'b0100101001: data <= 15'h00b5; 
        10'b0100101010: data <= 15'h008f; 
        10'b0100101011: data <= 15'h0094; 
        10'b0100101100: data <= 15'h0082; 
        10'b0100101101: data <= 15'h006f; 
        10'b0100101110: data <= 15'h0031; 
        10'b0100101111: data <= 15'h7fec; 
        10'b0100110000: data <= 15'h7fdf; 
        10'b0100110001: data <= 15'h7ff3; 
        10'b0100110010: data <= 15'h0003; 
        10'b0100110011: data <= 15'h7ffb; 
        10'b0100110100: data <= 15'h0013; 
        10'b0100110101: data <= 15'h000d; 
        10'b0100110110: data <= 15'h0018; 
        10'b0100110111: data <= 15'h0046; 
        10'b0100111000: data <= 15'h0054; 
        10'b0100111001: data <= 15'h002a; 
        10'b0100111010: data <= 15'h000f; 
        10'b0100111011: data <= 15'h000e; 
        10'b0100111100: data <= 15'h0004; 
        10'b0100111101: data <= 15'h0032; 
        10'b0100111110: data <= 15'h001a; 
        10'b0100111111: data <= 15'h0021; 
        10'b0101000000: data <= 15'h0036; 
        10'b0101000001: data <= 15'h0036; 
        10'b0101000010: data <= 15'h0038; 
        10'b0101000011: data <= 15'h00a4; 
        10'b0101000100: data <= 15'h00d5; 
        10'b0101000101: data <= 15'h008e; 
        10'b0101000110: data <= 15'h0090; 
        10'b0101000111: data <= 15'h006e; 
        10'b0101001000: data <= 15'h006b; 
        10'b0101001001: data <= 15'h0043; 
        10'b0101001010: data <= 15'h0031; 
        10'b0101001011: data <= 15'h7fef; 
        10'b0101001100: data <= 15'h7fcf; 
        10'b0101001101: data <= 15'h7fff; 
        10'b0101001110: data <= 15'h0005; 
        10'b0101001111: data <= 15'h0016; 
        10'b0101010000: data <= 15'h0011; 
        10'b0101010001: data <= 15'h7fff; 
        10'b0101010010: data <= 15'h000c; 
        10'b0101010011: data <= 15'h002c; 
        10'b0101010100: data <= 15'h0031; 
        10'b0101010101: data <= 15'h0008; 
        10'b0101010110: data <= 15'h000b; 
        10'b0101010111: data <= 15'h002f; 
        10'b0101011000: data <= 15'h0020; 
        10'b0101011001: data <= 15'h7ffe; 
        10'b0101011010: data <= 15'h7fda; 
        10'b0101011011: data <= 15'h7f9a; 
        10'b0101011100: data <= 15'h7f28; 
        10'b0101011101: data <= 15'h7eb1; 
        10'b0101011110: data <= 15'h7f06; 
        10'b0101011111: data <= 15'h0005; 
        10'b0101100000: data <= 15'h008d; 
        10'b0101100001: data <= 15'h0080; 
        10'b0101100010: data <= 15'h0032; 
        10'b0101100011: data <= 15'h0012; 
        10'b0101100100: data <= 15'h0003; 
        10'b0101100101: data <= 15'h7fee; 
        10'b0101100110: data <= 15'h7fef; 
        10'b0101100111: data <= 15'h7fe2; 
        10'b0101101000: data <= 15'h7fea; 
        10'b0101101001: data <= 15'h0014; 
        10'b0101101010: data <= 15'h000e; 
        10'b0101101011: data <= 15'h0000; 
        10'b0101101100: data <= 15'h0012; 
        10'b0101101101: data <= 15'h000b; 
        10'b0101101110: data <= 15'h0013; 
        10'b0101101111: data <= 15'h0028; 
        10'b0101110000: data <= 15'h000f; 
        10'b0101110001: data <= 15'h0006; 
        10'b0101110010: data <= 15'h7ff3; 
        10'b0101110011: data <= 15'h0009; 
        10'b0101110100: data <= 15'h7ffa; 
        10'b0101110101: data <= 15'h7fdf; 
        10'b0101110110: data <= 15'h7f95; 
        10'b0101110111: data <= 15'h7f1e; 
        10'b0101111000: data <= 15'h7e73; 
        10'b0101111001: data <= 15'h7e44; 
        10'b0101111010: data <= 15'h7f13; 
        10'b0101111011: data <= 15'h7fe1; 
        10'b0101111100: data <= 15'h0048; 
        10'b0101111101: data <= 15'h002f; 
        10'b0101111110: data <= 15'h000a; 
        10'b0101111111: data <= 15'h0015; 
        10'b0110000000: data <= 15'h7fd5; 
        10'b0110000001: data <= 15'h7fc8; 
        10'b0110000010: data <= 15'h7ff3; 
        10'b0110000011: data <= 15'h0004; 
        10'b0110000100: data <= 15'h7ff5; 
        10'b0110000101: data <= 15'h7ff8; 
        10'b0110000110: data <= 15'h000b; 
        10'b0110000111: data <= 15'h7ff5; 
        10'b0110001000: data <= 15'h7ffb; 
        10'b0110001001: data <= 15'h000a; 
        10'b0110001010: data <= 15'h0024; 
        10'b0110001011: data <= 15'h002c; 
        10'b0110001100: data <= 15'h001c; 
        10'b0110001101: data <= 15'h0021; 
        10'b0110001110: data <= 15'h7ff5; 
        10'b0110001111: data <= 15'h7fe9; 
        10'b0110010000: data <= 15'h7fce; 
        10'b0110010001: data <= 15'h7f8a; 
        10'b0110010010: data <= 15'h7f53; 
        10'b0110010011: data <= 15'h7ef4; 
        10'b0110010100: data <= 15'h7ea8; 
        10'b0110010101: data <= 15'h7ede; 
        10'b0110010110: data <= 15'h7f96; 
        10'b0110010111: data <= 15'h0002; 
        10'b0110011000: data <= 15'h0016; 
        10'b0110011001: data <= 15'h002e; 
        10'b0110011010: data <= 15'h0083; 
        10'b0110011011: data <= 15'h008d; 
        10'b0110011100: data <= 15'h0055; 
        10'b0110011101: data <= 15'h0036; 
        10'b0110011110: data <= 15'h0037; 
        10'b0110011111: data <= 15'h002f; 
        10'b0110100000: data <= 15'h0010; 
        10'b0110100001: data <= 15'h0005; 
        10'b0110100010: data <= 15'h7ff8; 
        10'b0110100011: data <= 15'h7ff9; 
        10'b0110100100: data <= 15'h000c; 
        10'b0110100101: data <= 15'h0011; 
        10'b0110100110: data <= 15'h0006; 
        10'b0110100111: data <= 15'h0011; 
        10'b0110101000: data <= 15'h0011; 
        10'b0110101001: data <= 15'h7fd0; 
        10'b0110101010: data <= 15'h7feb; 
        10'b0110101011: data <= 15'h7fe3; 
        10'b0110101100: data <= 15'h7f81; 
        10'b0110101101: data <= 15'h7f66; 
        10'b0110101110: data <= 15'h7f34; 
        10'b0110101111: data <= 15'h7f16; 
        10'b0110110000: data <= 15'h7f01; 
        10'b0110110001: data <= 15'h7f44; 
        10'b0110110010: data <= 15'h7f92; 
        10'b0110110011: data <= 15'h0003; 
        10'b0110110100: data <= 15'h000c; 
        10'b0110110101: data <= 15'h00b3; 
        10'b0110110110: data <= 15'h00d1; 
        10'b0110110111: data <= 15'h00ac; 
        10'b0110111000: data <= 15'h0099; 
        10'b0110111001: data <= 15'h0084; 
        10'b0110111010: data <= 15'h0055; 
        10'b0110111011: data <= 15'h0026; 
        10'b0110111100: data <= 15'h7ffe; 
        10'b0110111101: data <= 15'h7ff5; 
        10'b0110111110: data <= 15'h0003; 
        10'b0110111111: data <= 15'h0012; 
        10'b0111000000: data <= 15'h000b; 
        10'b0111000001: data <= 15'h0017; 
        10'b0111000010: data <= 15'h7ffe; 
        10'b0111000011: data <= 15'h0018; 
        10'b0111000100: data <= 15'h0013; 
        10'b0111000101: data <= 15'h7feb; 
        10'b0111000110: data <= 15'h7fe2; 
        10'b0111000111: data <= 15'h7ffc; 
        10'b0111001000: data <= 15'h7f9a; 
        10'b0111001001: data <= 15'h7f8d; 
        10'b0111001010: data <= 15'h7f47; 
        10'b0111001011: data <= 15'h7f24; 
        10'b0111001100: data <= 15'h7f76; 
        10'b0111001101: data <= 15'h7fb3; 
        10'b0111001110: data <= 15'h7f90; 
        10'b0111001111: data <= 15'h003a; 
        10'b0111010000: data <= 15'h0046; 
        10'b0111010001: data <= 15'h0097; 
        10'b0111010010: data <= 15'h0082; 
        10'b0111010011: data <= 15'h0088; 
        10'b0111010100: data <= 15'h006c; 
        10'b0111010101: data <= 15'h0052; 
        10'b0111010110: data <= 15'h0010; 
        10'b0111010111: data <= 15'h7fde; 
        10'b0111011000: data <= 15'h7feb; 
        10'b0111011001: data <= 15'h7ff4; 
        10'b0111011010: data <= 15'h000d; 
        10'b0111011011: data <= 15'h0016; 
        10'b0111011100: data <= 15'h0001; 
        10'b0111011101: data <= 15'h0003; 
        10'b0111011110: data <= 15'h000e; 
        10'b0111011111: data <= 15'h7fff; 
        10'b0111100000: data <= 15'h0005; 
        10'b0111100001: data <= 15'h7ff2; 
        10'b0111100010: data <= 15'h7fbb; 
        10'b0111100011: data <= 15'h7fa6; 
        10'b0111100100: data <= 15'h7f8e; 
        10'b0111100101: data <= 15'h7fa2; 
        10'b0111100110: data <= 15'h7f84; 
        10'b0111100111: data <= 15'h7fa4; 
        10'b0111101000: data <= 15'h7fe3; 
        10'b0111101001: data <= 15'h0017; 
        10'b0111101010: data <= 15'h000d; 
        10'b0111101011: data <= 15'h0017; 
        10'b0111101100: data <= 15'h7ff2; 
        10'b0111101101: data <= 15'h0024; 
        10'b0111101110: data <= 15'h0020; 
        10'b0111101111: data <= 15'h0017; 
        10'b0111110000: data <= 15'h000c; 
        10'b0111110001: data <= 15'h7fed; 
        10'b0111110010: data <= 15'h7fd6; 
        10'b0111110011: data <= 15'h7fed; 
        10'b0111110100: data <= 15'h7ff0; 
        10'b0111110101: data <= 15'h7ff3; 
        10'b0111110110: data <= 15'h7ff9; 
        10'b0111110111: data <= 15'h7ffa; 
        10'b0111111000: data <= 15'h7ffa; 
        10'b0111111001: data <= 15'h7ffe; 
        10'b0111111010: data <= 15'h0010; 
        10'b0111111011: data <= 15'h0005; 
        10'b0111111100: data <= 15'h7fe4; 
        10'b0111111101: data <= 15'h7fbe; 
        10'b0111111110: data <= 15'h7f93; 
        10'b0111111111: data <= 15'h7f78; 
        10'b1000000000: data <= 15'h7f82; 
        10'b1000000001: data <= 15'h7f8a; 
        10'b1000000010: data <= 15'h7f68; 
        10'b1000000011: data <= 15'h7fcc; 
        10'b1000000100: data <= 15'h7ff0; 
        10'b1000000101: data <= 15'h0002; 
        10'b1000000110: data <= 15'h002b; 
        10'b1000000111: data <= 15'h7fd3; 
        10'b1000001000: data <= 15'h7fc9; 
        10'b1000001001: data <= 15'h7fe1; 
        10'b1000001010: data <= 15'h7fba; 
        10'b1000001011: data <= 15'h7fd5; 
        10'b1000001100: data <= 15'h7fb8; 
        10'b1000001101: data <= 15'h7f92; 
        10'b1000001110: data <= 15'h7faf; 
        10'b1000001111: data <= 15'h7fcd; 
        10'b1000010000: data <= 15'h7fd8; 
        10'b1000010001: data <= 15'h0004; 
        10'b1000010010: data <= 15'h7ffc; 
        10'b1000010011: data <= 15'h0001; 
        10'b1000010100: data <= 15'h0016; 
        10'b1000010101: data <= 15'h0017; 
        10'b1000010110: data <= 15'h0015; 
        10'b1000010111: data <= 15'h000b; 
        10'b1000011000: data <= 15'h7fed; 
        10'b1000011001: data <= 15'h7faa; 
        10'b1000011010: data <= 15'h7f76; 
        10'b1000011011: data <= 15'h7f6c; 
        10'b1000011100: data <= 15'h7f68; 
        10'b1000011101: data <= 15'h7f67; 
        10'b1000011110: data <= 15'h7f99; 
        10'b1000011111: data <= 15'h7fb6; 
        10'b1000100000: data <= 15'h7fd4; 
        10'b1000100001: data <= 15'h0013; 
        10'b1000100010: data <= 15'h003c; 
        10'b1000100011: data <= 15'h7fc1; 
        10'b1000100100: data <= 15'h7fc2; 
        10'b1000100101: data <= 15'h7fb2; 
        10'b1000100110: data <= 15'h7f84; 
        10'b1000100111: data <= 15'h7f8b; 
        10'b1000101000: data <= 15'h7f70; 
        10'b1000101001: data <= 15'h7f7b; 
        10'b1000101010: data <= 15'h7f9b; 
        10'b1000101011: data <= 15'h7fba; 
        10'b1000101100: data <= 15'h7fdd; 
        10'b1000101101: data <= 15'h7ff3; 
        10'b1000101110: data <= 15'h0016; 
        10'b1000101111: data <= 15'h7ff6; 
        10'b1000110000: data <= 15'h7ff4; 
        10'b1000110001: data <= 15'h7ffb; 
        10'b1000110010: data <= 15'h0009; 
        10'b1000110011: data <= 15'h7ffc; 
        10'b1000110100: data <= 15'h7fea; 
        10'b1000110101: data <= 15'h7fbe; 
        10'b1000110110: data <= 15'h7f75; 
        10'b1000110111: data <= 15'h7f6f; 
        10'b1000111000: data <= 15'h7f78; 
        10'b1000111001: data <= 15'h7f7b; 
        10'b1000111010: data <= 15'h7fa3; 
        10'b1000111011: data <= 15'h7fa0; 
        10'b1000111100: data <= 15'h0007; 
        10'b1000111101: data <= 15'h000a; 
        10'b1000111110: data <= 15'h0020; 
        10'b1000111111: data <= 15'h7fab; 
        10'b1001000000: data <= 15'h7f96; 
        10'b1001000001: data <= 15'h7f76; 
        10'b1001000010: data <= 15'h7f41; 
        10'b1001000011: data <= 15'h7f87; 
        10'b1001000100: data <= 15'h7f59; 
        10'b1001000101: data <= 15'h7f81; 
        10'b1001000110: data <= 15'h7fa4; 
        10'b1001000111: data <= 15'h7fd9; 
        10'b1001001000: data <= 15'h7fe6; 
        10'b1001001001: data <= 15'h0014; 
        10'b1001001010: data <= 15'h0013; 
        10'b1001001011: data <= 15'h000d; 
        10'b1001001100: data <= 15'h0012; 
        10'b1001001101: data <= 15'h0013; 
        10'b1001001110: data <= 15'h0004; 
        10'b1001001111: data <= 15'h7fe8; 
        10'b1001010000: data <= 15'h7ff4; 
        10'b1001010001: data <= 15'h7fc5; 
        10'b1001010010: data <= 15'h7fbb; 
        10'b1001010011: data <= 15'h7f9c; 
        10'b1001010100: data <= 15'h7fa6; 
        10'b1001010101: data <= 15'h7fca; 
        10'b1001010110: data <= 15'h7fb4; 
        10'b1001010111: data <= 15'h7fc2; 
        10'b1001011000: data <= 15'h7fe4; 
        10'b1001011001: data <= 15'h0004; 
        10'b1001011010: data <= 15'h7fef; 
        10'b1001011011: data <= 15'h7fc7; 
        10'b1001011100: data <= 15'h7fbe; 
        10'b1001011101: data <= 15'h7f78; 
        10'b1001011110: data <= 15'h7f78; 
        10'b1001011111: data <= 15'h7f78; 
        10'b1001100000: data <= 15'h7f71; 
        10'b1001100001: data <= 15'h7f87; 
        10'b1001100010: data <= 15'h7fb9; 
        10'b1001100011: data <= 15'h7fca; 
        10'b1001100100: data <= 15'h7ffe; 
        10'b1001100101: data <= 15'h0008; 
        10'b1001100110: data <= 15'h0012; 
        10'b1001100111: data <= 15'h7ffc; 
        10'b1001101000: data <= 15'h0006; 
        10'b1001101001: data <= 15'h0001; 
        10'b1001101010: data <= 15'h0005; 
        10'b1001101011: data <= 15'h7ff1; 
        10'b1001101100: data <= 15'h7ff9; 
        10'b1001101101: data <= 15'h0009; 
        10'b1001101110: data <= 15'h7fea; 
        10'b1001101111: data <= 15'h000b; 
        10'b1001110000: data <= 15'h0011; 
        10'b1001110001: data <= 15'h7fe5; 
        10'b1001110010: data <= 15'h7fcc; 
        10'b1001110011: data <= 15'h7fa7; 
        10'b1001110100: data <= 15'h7fad; 
        10'b1001110101: data <= 15'h7fde; 
        10'b1001110110: data <= 15'h000a; 
        10'b1001110111: data <= 15'h000a; 
        10'b1001111000: data <= 15'h7fcc; 
        10'b1001111001: data <= 15'h7fc0; 
        10'b1001111010: data <= 15'h7f93; 
        10'b1001111011: data <= 15'h7f93; 
        10'b1001111100: data <= 15'h7f85; 
        10'b1001111101: data <= 15'h7f94; 
        10'b1001111110: data <= 15'h7fc9; 
        10'b1001111111: data <= 15'h7fee; 
        10'b1010000000: data <= 15'h000c; 
        10'b1010000001: data <= 15'h7ff4; 
        10'b1010000010: data <= 15'h0006; 
        10'b1010000011: data <= 15'h0000; 
        10'b1010000100: data <= 15'h0008; 
        10'b1010000101: data <= 15'h0011; 
        10'b1010000110: data <= 15'h7ff3; 
        10'b1010000111: data <= 15'h7ff4; 
        10'b1010001000: data <= 15'h0017; 
        10'b1010001001: data <= 15'h001e; 
        10'b1010001010: data <= 15'h0042; 
        10'b1010001011: data <= 15'h0057; 
        10'b1010001100: data <= 15'h002a; 
        10'b1010001101: data <= 15'h0008; 
        10'b1010001110: data <= 15'h7fe6; 
        10'b1010001111: data <= 15'h7fc5; 
        10'b1010010000: data <= 15'h7fcf; 
        10'b1010010001: data <= 15'h0003; 
        10'b1010010010: data <= 15'h0022; 
        10'b1010010011: data <= 15'h001f; 
        10'b1010010100: data <= 15'h7ff3; 
        10'b1010010101: data <= 15'h7fed; 
        10'b1010010110: data <= 15'h7fba; 
        10'b1010010111: data <= 15'h7f9f; 
        10'b1010011000: data <= 15'h7f9c; 
        10'b1010011001: data <= 15'h7fb2; 
        10'b1010011010: data <= 15'h7fc0; 
        10'b1010011011: data <= 15'h7fd6; 
        10'b1010011100: data <= 15'h7fee; 
        10'b1010011101: data <= 15'h0001; 
        10'b1010011110: data <= 15'h0001; 
        10'b1010011111: data <= 15'h7ff9; 
        10'b1010100000: data <= 15'h0000; 
        10'b1010100001: data <= 15'h7ffe; 
        10'b1010100010: data <= 15'h0006; 
        10'b1010100011: data <= 15'h000f; 
        10'b1010100100: data <= 15'h001f; 
        10'b1010100101: data <= 15'h0048; 
        10'b1010100110: data <= 15'h006d; 
        10'b1010100111: data <= 15'h007b; 
        10'b1010101000: data <= 15'h0068; 
        10'b1010101001: data <= 15'h0036; 
        10'b1010101010: data <= 15'h0074; 
        10'b1010101011: data <= 15'h0044; 
        10'b1010101100: data <= 15'h003b; 
        10'b1010101101: data <= 15'h0054; 
        10'b1010101110: data <= 15'h0033; 
        10'b1010101111: data <= 15'h004a; 
        10'b1010110000: data <= 15'h002c; 
        10'b1010110001: data <= 15'h0022; 
        10'b1010110010: data <= 15'h7ffe; 
        10'b1010110011: data <= 15'h7fe0; 
        10'b1010110100: data <= 15'h7fde; 
        10'b1010110101: data <= 15'h7fd7; 
        10'b1010110110: data <= 15'h7fd1; 
        10'b1010110111: data <= 15'h7fd6; 
        10'b1010111000: data <= 15'h0006; 
        10'b1010111001: data <= 15'h7ffd; 
        10'b1010111010: data <= 15'h7ff5; 
        10'b1010111011: data <= 15'h000d; 
        10'b1010111100: data <= 15'h7ff5; 
        10'b1010111101: data <= 15'h000a; 
        10'b1010111110: data <= 15'h0013; 
        10'b1010111111: data <= 15'h0012; 
        10'b1011000000: data <= 15'h000a; 
        10'b1011000001: data <= 15'h0024; 
        10'b1011000010: data <= 15'h0035; 
        10'b1011000011: data <= 15'h0052; 
        10'b1011000100: data <= 15'h007f; 
        10'b1011000101: data <= 15'h007c; 
        10'b1011000110: data <= 15'h0093; 
        10'b1011000111: data <= 15'h0088; 
        10'b1011001000: data <= 15'h007a; 
        10'b1011001001: data <= 15'h0060; 
        10'b1011001010: data <= 15'h0062; 
        10'b1011001011: data <= 15'h0068; 
        10'b1011001100: data <= 15'h0057; 
        10'b1011001101: data <= 15'h0052; 
        10'b1011001110: data <= 15'h0042; 
        10'b1011001111: data <= 15'h0017; 
        10'b1011010000: data <= 15'h7fe4; 
        10'b1011010001: data <= 15'h0004; 
        10'b1011010010: data <= 15'h7ff2; 
        10'b1011010011: data <= 15'h7ff6; 
        10'b1011010100: data <= 15'h7ffd; 
        10'b1011010101: data <= 15'h0006; 
        10'b1011010110: data <= 15'h0019; 
        10'b1011010111: data <= 15'h0010; 
        10'b1011011000: data <= 15'h7ff7; 
        10'b1011011001: data <= 15'h0005; 
        10'b1011011010: data <= 15'h0017; 
        10'b1011011011: data <= 15'h7ffc; 
        10'b1011011100: data <= 15'h7ff8; 
        10'b1011011101: data <= 15'h0016; 
        10'b1011011110: data <= 15'h0002; 
        10'b1011011111: data <= 15'h0014; 
        10'b1011100000: data <= 15'h0013; 
        10'b1011100001: data <= 15'h0003; 
        10'b1011100010: data <= 15'h001c; 
        10'b1011100011: data <= 15'h0029; 
        10'b1011100100: data <= 15'h000c; 
        10'b1011100101: data <= 15'h0023; 
        10'b1011100110: data <= 15'h004b; 
        10'b1011100111: data <= 15'h005c; 
        10'b1011101000: data <= 15'h0049; 
        10'b1011101001: data <= 15'h005d; 
        10'b1011101010: data <= 15'h0035; 
        10'b1011101011: data <= 15'h0019; 
        10'b1011101100: data <= 15'h0001; 
        10'b1011101101: data <= 15'h000a; 
        10'b1011101110: data <= 15'h7ffd; 
        10'b1011101111: data <= 15'h0005; 
        10'b1011110000: data <= 15'h0001; 
        10'b1011110001: data <= 15'h7ffa; 
        10'b1011110010: data <= 15'h7fff; 
        10'b1011110011: data <= 15'h7ffd; 
        10'b1011110100: data <= 15'h7ff4; 
        10'b1011110101: data <= 15'h0009; 
        10'b1011110110: data <= 15'h0006; 
        10'b1011110111: data <= 15'h000c; 
        10'b1011111000: data <= 15'h0010; 
        10'b1011111001: data <= 15'h000a; 
        10'b1011111010: data <= 15'h0004; 
        10'b1011111011: data <= 15'h0002; 
        10'b1011111100: data <= 15'h001a; 
        10'b1011111101: data <= 15'h0010; 
        10'b1011111110: data <= 15'h0005; 
        10'b1011111111: data <= 15'h0010; 
        10'b1100000000: data <= 15'h0008; 
        10'b1100000001: data <= 15'h001e; 
        10'b1100000010: data <= 15'h0012; 
        10'b1100000011: data <= 15'h000e; 
        10'b1100000100: data <= 15'h002a; 
        10'b1100000101: data <= 15'h000e; 
        10'b1100000110: data <= 15'h000d; 
        10'b1100000111: data <= 15'h001d; 
        10'b1100001000: data <= 15'h0003; 
        10'b1100001001: data <= 15'h7ffb; 
        10'b1100001010: data <= 15'h0018; 
        10'b1100001011: data <= 15'h000d; 
        10'b1100001100: data <= 15'h0006; 
        10'b1100001101: data <= 15'h7ffc; 
        10'b1100001110: data <= 15'h7ff6; 
        10'b1100001111: data <= 15'h0010; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 10) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 16'h0003; 
        10'b0000000001: data <= 16'h0004; 
        10'b0000000010: data <= 16'h001e; 
        10'b0000000011: data <= 16'h000c; 
        10'b0000000100: data <= 16'h0032; 
        10'b0000000101: data <= 16'hffea; 
        10'b0000000110: data <= 16'hfff1; 
        10'b0000000111: data <= 16'h0010; 
        10'b0000001000: data <= 16'h0026; 
        10'b0000001001: data <= 16'h0025; 
        10'b0000001010: data <= 16'hffeb; 
        10'b0000001011: data <= 16'h000a; 
        10'b0000001100: data <= 16'h000b; 
        10'b0000001101: data <= 16'hfffa; 
        10'b0000001110: data <= 16'h0028; 
        10'b0000001111: data <= 16'h000b; 
        10'b0000010000: data <= 16'h0001; 
        10'b0000010001: data <= 16'hffff; 
        10'b0000010010: data <= 16'h0004; 
        10'b0000010011: data <= 16'h000e; 
        10'b0000010100: data <= 16'h001a; 
        10'b0000010101: data <= 16'h0030; 
        10'b0000010110: data <= 16'hfff3; 
        10'b0000010111: data <= 16'h0024; 
        10'b0000011000: data <= 16'hfffb; 
        10'b0000011001: data <= 16'h001a; 
        10'b0000011010: data <= 16'hfffe; 
        10'b0000011011: data <= 16'h0000; 
        10'b0000011100: data <= 16'h002e; 
        10'b0000011101: data <= 16'hfff6; 
        10'b0000011110: data <= 16'h000a; 
        10'b0000011111: data <= 16'h002d; 
        10'b0000100000: data <= 16'h0011; 
        10'b0000100001: data <= 16'h0002; 
        10'b0000100010: data <= 16'h002d; 
        10'b0000100011: data <= 16'h000e; 
        10'b0000100100: data <= 16'h0004; 
        10'b0000100101: data <= 16'hfff8; 
        10'b0000100110: data <= 16'hfffa; 
        10'b0000100111: data <= 16'hffe9; 
        10'b0000101000: data <= 16'h0026; 
        10'b0000101001: data <= 16'hfffd; 
        10'b0000101010: data <= 16'h002e; 
        10'b0000101011: data <= 16'hfff4; 
        10'b0000101100: data <= 16'h0014; 
        10'b0000101101: data <= 16'h0023; 
        10'b0000101110: data <= 16'h0027; 
        10'b0000101111: data <= 16'h001f; 
        10'b0000110000: data <= 16'h0001; 
        10'b0000110001: data <= 16'h001f; 
        10'b0000110010: data <= 16'hffff; 
        10'b0000110011: data <= 16'h0031; 
        10'b0000110100: data <= 16'h0025; 
        10'b0000110101: data <= 16'hfff2; 
        10'b0000110110: data <= 16'hfff3; 
        10'b0000110111: data <= 16'h0014; 
        10'b0000111000: data <= 16'h002b; 
        10'b0000111001: data <= 16'h002b; 
        10'b0000111010: data <= 16'h0022; 
        10'b0000111011: data <= 16'hfffa; 
        10'b0000111100: data <= 16'h0027; 
        10'b0000111101: data <= 16'hffee; 
        10'b0000111110: data <= 16'hfff1; 
        10'b0000111111: data <= 16'h001e; 
        10'b0001000000: data <= 16'h001a; 
        10'b0001000001: data <= 16'hfff1; 
        10'b0001000010: data <= 16'hfffd; 
        10'b0001000011: data <= 16'h0013; 
        10'b0001000100: data <= 16'hfffb; 
        10'b0001000101: data <= 16'hfff6; 
        10'b0001000110: data <= 16'h000c; 
        10'b0001000111: data <= 16'h0027; 
        10'b0001001000: data <= 16'h0020; 
        10'b0001001001: data <= 16'h0006; 
        10'b0001001010: data <= 16'h000f; 
        10'b0001001011: data <= 16'h002c; 
        10'b0001001100: data <= 16'h0026; 
        10'b0001001101: data <= 16'h002b; 
        10'b0001001110: data <= 16'hffea; 
        10'b0001001111: data <= 16'h0022; 
        10'b0001010000: data <= 16'h000d; 
        10'b0001010001: data <= 16'h001e; 
        10'b0001010010: data <= 16'h001a; 
        10'b0001010011: data <= 16'h0026; 
        10'b0001010100: data <= 16'hfffd; 
        10'b0001010101: data <= 16'h0003; 
        10'b0001010110: data <= 16'h0028; 
        10'b0001010111: data <= 16'hfffa; 
        10'b0001011000: data <= 16'h0004; 
        10'b0001011001: data <= 16'hfffd; 
        10'b0001011010: data <= 16'hfff1; 
        10'b0001011011: data <= 16'h001a; 
        10'b0001011100: data <= 16'h0000; 
        10'b0001011101: data <= 16'h001a; 
        10'b0001011110: data <= 16'hffeb; 
        10'b0001011111: data <= 16'h0005; 
        10'b0001100000: data <= 16'h0015; 
        10'b0001100001: data <= 16'hffe3; 
        10'b0001100010: data <= 16'h0018; 
        10'b0001100011: data <= 16'hffed; 
        10'b0001100100: data <= 16'hffd6; 
        10'b0001100101: data <= 16'hffde; 
        10'b0001100110: data <= 16'hffe3; 
        10'b0001100111: data <= 16'hffec; 
        10'b0001101000: data <= 16'hfffb; 
        10'b0001101001: data <= 16'hffee; 
        10'b0001101010: data <= 16'h0010; 
        10'b0001101011: data <= 16'hfffe; 
        10'b0001101100: data <= 16'h0013; 
        10'b0001101101: data <= 16'h0031; 
        10'b0001101110: data <= 16'hfff0; 
        10'b0001101111: data <= 16'h0014; 
        10'b0001110000: data <= 16'h002f; 
        10'b0001110001: data <= 16'hffef; 
        10'b0001110010: data <= 16'h001a; 
        10'b0001110011: data <= 16'hffec; 
        10'b0001110100: data <= 16'h000b; 
        10'b0001110101: data <= 16'hfff7; 
        10'b0001110110: data <= 16'h0002; 
        10'b0001110111: data <= 16'hffed; 
        10'b0001111000: data <= 16'h000f; 
        10'b0001111001: data <= 16'hfff9; 
        10'b0001111010: data <= 16'hffd2; 
        10'b0001111011: data <= 16'hffa7; 
        10'b0001111100: data <= 16'hffa2; 
        10'b0001111101: data <= 16'hffa6; 
        10'b0001111110: data <= 16'hff95; 
        10'b0001111111: data <= 16'hff50; 
        10'b0010000000: data <= 16'hff98; 
        10'b0010000001: data <= 16'hffb2; 
        10'b0010000010: data <= 16'hffbc; 
        10'b0010000011: data <= 16'hffee; 
        10'b0010000100: data <= 16'hffcd; 
        10'b0010000101: data <= 16'h0018; 
        10'b0010000110: data <= 16'h0004; 
        10'b0010000111: data <= 16'hffe7; 
        10'b0010001000: data <= 16'h002d; 
        10'b0010001001: data <= 16'hfffe; 
        10'b0010001010: data <= 16'h002c; 
        10'b0010001011: data <= 16'h002b; 
        10'b0010001100: data <= 16'h0028; 
        10'b0010001101: data <= 16'h0002; 
        10'b0010001110: data <= 16'h0027; 
        10'b0010001111: data <= 16'hfff5; 
        10'b0010010000: data <= 16'hffe2; 
        10'b0010010001: data <= 16'hfffb; 
        10'b0010010010: data <= 16'hffe9; 
        10'b0010010011: data <= 16'hfff7; 
        10'b0010010100: data <= 16'hffe4; 
        10'b0010010101: data <= 16'hffc0; 
        10'b0010010110: data <= 16'hff63; 
        10'b0010010111: data <= 16'hff3f; 
        10'b0010011000: data <= 16'hff0d; 
        10'b0010011001: data <= 16'hfee3; 
        10'b0010011010: data <= 16'hfe9d; 
        10'b0010011011: data <= 16'hfe9f; 
        10'b0010011100: data <= 16'hfe8e; 
        10'b0010011101: data <= 16'hfeba; 
        10'b0010011110: data <= 16'hfeeb; 
        10'b0010011111: data <= 16'hff2e; 
        10'b0010100000: data <= 16'hff6b; 
        10'b0010100001: data <= 16'hffcb; 
        10'b0010100010: data <= 16'hffae; 
        10'b0010100011: data <= 16'hfff6; 
        10'b0010100100: data <= 16'h0024; 
        10'b0010100101: data <= 16'h001d; 
        10'b0010100110: data <= 16'hfff9; 
        10'b0010100111: data <= 16'h0002; 
        10'b0010101000: data <= 16'h0022; 
        10'b0010101001: data <= 16'h002e; 
        10'b0010101010: data <= 16'h0003; 
        10'b0010101011: data <= 16'h0007; 
        10'b0010101100: data <= 16'h0032; 
        10'b0010101101: data <= 16'h003b; 
        10'b0010101110: data <= 16'h0045; 
        10'b0010101111: data <= 16'h0068; 
        10'b0010110000: data <= 16'h009b; 
        10'b0010110001: data <= 16'h007c; 
        10'b0010110010: data <= 16'h0084; 
        10'b0010110011: data <= 16'h0018; 
        10'b0010110100: data <= 16'hff96; 
        10'b0010110101: data <= 16'hff22; 
        10'b0010110110: data <= 16'hff19; 
        10'b0010110111: data <= 16'hff88; 
        10'b0010111000: data <= 16'hffb7; 
        10'b0010111001: data <= 16'hffa9; 
        10'b0010111010: data <= 16'hff97; 
        10'b0010111011: data <= 16'hff86; 
        10'b0010111100: data <= 16'hff48; 
        10'b0010111101: data <= 16'hffbb; 
        10'b0010111110: data <= 16'hff7f; 
        10'b0010111111: data <= 16'hffa2; 
        10'b0011000000: data <= 16'hffc1; 
        10'b0011000001: data <= 16'hffeb; 
        10'b0011000010: data <= 16'hffea; 
        10'b0011000011: data <= 16'h0005; 
        10'b0011000100: data <= 16'h001f; 
        10'b0011000101: data <= 16'h002e; 
        10'b0011000110: data <= 16'h0026; 
        10'b0011000111: data <= 16'h005a; 
        10'b0011001000: data <= 16'h006d; 
        10'b0011001001: data <= 16'h0062; 
        10'b0011001010: data <= 16'h008e; 
        10'b0011001011: data <= 16'h00d9; 
        10'b0011001100: data <= 16'h012a; 
        10'b0011001101: data <= 16'h00ec; 
        10'b0011001110: data <= 16'h00a3; 
        10'b0011001111: data <= 16'h00b3; 
        10'b0011010000: data <= 16'h00bf; 
        10'b0011010001: data <= 16'h0025; 
        10'b0011010010: data <= 16'h001b; 
        10'b0011010011: data <= 16'h0044; 
        10'b0011010100: data <= 16'h00c9; 
        10'b0011010101: data <= 16'h00e0; 
        10'b0011010110: data <= 16'h0098; 
        10'b0011010111: data <= 16'h007a; 
        10'b0011011000: data <= 16'h001e; 
        10'b0011011001: data <= 16'hffde; 
        10'b0011011010: data <= 16'h0010; 
        10'b0011011011: data <= 16'hffdc; 
        10'b0011011100: data <= 16'hffde; 
        10'b0011011101: data <= 16'hfffe; 
        10'b0011011110: data <= 16'h0018; 
        10'b0011011111: data <= 16'hfff7; 
        10'b0011100000: data <= 16'hffe9; 
        10'b0011100001: data <= 16'h0030; 
        10'b0011100010: data <= 16'h0013; 
        10'b0011100011: data <= 16'h004c; 
        10'b0011100100: data <= 16'h009a; 
        10'b0011100101: data <= 16'h008b; 
        10'b0011100110: data <= 16'h00ba; 
        10'b0011100111: data <= 16'h014e; 
        10'b0011101000: data <= 16'h00e1; 
        10'b0011101001: data <= 16'h009b; 
        10'b0011101010: data <= 16'h00c5; 
        10'b0011101011: data <= 16'h0108; 
        10'b0011101100: data <= 16'h00fb; 
        10'b0011101101: data <= 16'h007e; 
        10'b0011101110: data <= 16'h004a; 
        10'b0011101111: data <= 16'h0066; 
        10'b0011110000: data <= 16'h00b2; 
        10'b0011110001: data <= 16'h0111; 
        10'b0011110010: data <= 16'h00bb; 
        10'b0011110011: data <= 16'h00a0; 
        10'b0011110100: data <= 16'h0080; 
        10'b0011110101: data <= 16'h0003; 
        10'b0011110110: data <= 16'h004e; 
        10'b0011110111: data <= 16'h0042; 
        10'b0011111000: data <= 16'hffd1; 
        10'b0011111001: data <= 16'hffea; 
        10'b0011111010: data <= 16'h001a; 
        10'b0011111011: data <= 16'h0028; 
        10'b0011111100: data <= 16'h0015; 
        10'b0011111101: data <= 16'h0027; 
        10'b0011111110: data <= 16'h0034; 
        10'b0011111111: data <= 16'h006e; 
        10'b0100000000: data <= 16'h0097; 
        10'b0100000001: data <= 16'h00ab; 
        10'b0100000010: data <= 16'h003f; 
        10'b0100000011: data <= 16'h0054; 
        10'b0100000100: data <= 16'h005f; 
        10'b0100000101: data <= 16'h003f; 
        10'b0100000110: data <= 16'h009a; 
        10'b0100000111: data <= 16'h00bc; 
        10'b0100001000: data <= 16'h00f0; 
        10'b0100001001: data <= 16'h00c3; 
        10'b0100001010: data <= 16'h0118; 
        10'b0100001011: data <= 16'h0158; 
        10'b0100001100: data <= 16'h013d; 
        10'b0100001101: data <= 16'h0162; 
        10'b0100001110: data <= 16'h00e7; 
        10'b0100001111: data <= 16'h00eb; 
        10'b0100010000: data <= 16'h00c6; 
        10'b0100010001: data <= 16'h00a5; 
        10'b0100010010: data <= 16'h004e; 
        10'b0100010011: data <= 16'hffe4; 
        10'b0100010100: data <= 16'hffd0; 
        10'b0100010101: data <= 16'hffe8; 
        10'b0100010110: data <= 16'h0015; 
        10'b0100010111: data <= 16'hfff5; 
        10'b0100011000: data <= 16'h0008; 
        10'b0100011001: data <= 16'h002a; 
        10'b0100011010: data <= 16'h002f; 
        10'b0100011011: data <= 16'h0088; 
        10'b0100011100: data <= 16'h009c; 
        10'b0100011101: data <= 16'h0082; 
        10'b0100011110: data <= 16'h0018; 
        10'b0100011111: data <= 16'h0027; 
        10'b0100100000: data <= 16'hffcb; 
        10'b0100100001: data <= 16'hfffe; 
        10'b0100100010: data <= 16'h005f; 
        10'b0100100011: data <= 16'h00a8; 
        10'b0100100100: data <= 16'h0075; 
        10'b0100100101: data <= 16'h0110; 
        10'b0100100110: data <= 16'h015d; 
        10'b0100100111: data <= 16'h01ad; 
        10'b0100101000: data <= 16'h01e9; 
        10'b0100101001: data <= 16'h016a; 
        10'b0100101010: data <= 16'h011d; 
        10'b0100101011: data <= 16'h0129; 
        10'b0100101100: data <= 16'h0104; 
        10'b0100101101: data <= 16'h00dd; 
        10'b0100101110: data <= 16'h0062; 
        10'b0100101111: data <= 16'hffd8; 
        10'b0100110000: data <= 16'hffbe; 
        10'b0100110001: data <= 16'hffe5; 
        10'b0100110010: data <= 16'h0005; 
        10'b0100110011: data <= 16'hfff6; 
        10'b0100110100: data <= 16'h0025; 
        10'b0100110101: data <= 16'h001a; 
        10'b0100110110: data <= 16'h002f; 
        10'b0100110111: data <= 16'h008c; 
        10'b0100111000: data <= 16'h00a8; 
        10'b0100111001: data <= 16'h0053; 
        10'b0100111010: data <= 16'h001e; 
        10'b0100111011: data <= 16'h001b; 
        10'b0100111100: data <= 16'h0008; 
        10'b0100111101: data <= 16'h0065; 
        10'b0100111110: data <= 16'h0034; 
        10'b0100111111: data <= 16'h0042; 
        10'b0101000000: data <= 16'h006d; 
        10'b0101000001: data <= 16'h006c; 
        10'b0101000010: data <= 16'h0070; 
        10'b0101000011: data <= 16'h0148; 
        10'b0101000100: data <= 16'h01aa; 
        10'b0101000101: data <= 16'h011c; 
        10'b0101000110: data <= 16'h011f; 
        10'b0101000111: data <= 16'h00dd; 
        10'b0101001000: data <= 16'h00d6; 
        10'b0101001001: data <= 16'h0087; 
        10'b0101001010: data <= 16'h0061; 
        10'b0101001011: data <= 16'hffde; 
        10'b0101001100: data <= 16'hff9d; 
        10'b0101001101: data <= 16'hfffd; 
        10'b0101001110: data <= 16'h0009; 
        10'b0101001111: data <= 16'h002b; 
        10'b0101010000: data <= 16'h0021; 
        10'b0101010001: data <= 16'hfffe; 
        10'b0101010010: data <= 16'h0017; 
        10'b0101010011: data <= 16'h0058; 
        10'b0101010100: data <= 16'h0063; 
        10'b0101010101: data <= 16'h0010; 
        10'b0101010110: data <= 16'h0016; 
        10'b0101010111: data <= 16'h005e; 
        10'b0101011000: data <= 16'h0040; 
        10'b0101011001: data <= 16'hfffc; 
        10'b0101011010: data <= 16'hffb3; 
        10'b0101011011: data <= 16'hff34; 
        10'b0101011100: data <= 16'hfe50; 
        10'b0101011101: data <= 16'hfd63; 
        10'b0101011110: data <= 16'hfe0b; 
        10'b0101011111: data <= 16'h000b; 
        10'b0101100000: data <= 16'h011b; 
        10'b0101100001: data <= 16'h0101; 
        10'b0101100010: data <= 16'h0065; 
        10'b0101100011: data <= 16'h0024; 
        10'b0101100100: data <= 16'h0007; 
        10'b0101100101: data <= 16'hffdb; 
        10'b0101100110: data <= 16'hffde; 
        10'b0101100111: data <= 16'hffc4; 
        10'b0101101000: data <= 16'hffd4; 
        10'b0101101001: data <= 16'h0029; 
        10'b0101101010: data <= 16'h001d; 
        10'b0101101011: data <= 16'h0000; 
        10'b0101101100: data <= 16'h0024; 
        10'b0101101101: data <= 16'h0015; 
        10'b0101101110: data <= 16'h0027; 
        10'b0101101111: data <= 16'h0050; 
        10'b0101110000: data <= 16'h001e; 
        10'b0101110001: data <= 16'h000d; 
        10'b0101110010: data <= 16'hffe6; 
        10'b0101110011: data <= 16'h0011; 
        10'b0101110100: data <= 16'hfff4; 
        10'b0101110101: data <= 16'hffbe; 
        10'b0101110110: data <= 16'hff29; 
        10'b0101110111: data <= 16'hfe3c; 
        10'b0101111000: data <= 16'hfce6; 
        10'b0101111001: data <= 16'hfc89; 
        10'b0101111010: data <= 16'hfe25; 
        10'b0101111011: data <= 16'hffc2; 
        10'b0101111100: data <= 16'h0090; 
        10'b0101111101: data <= 16'h005d; 
        10'b0101111110: data <= 16'h0014; 
        10'b0101111111: data <= 16'h002a; 
        10'b0110000000: data <= 16'hffa9; 
        10'b0110000001: data <= 16'hff91; 
        10'b0110000010: data <= 16'hffe6; 
        10'b0110000011: data <= 16'h0008; 
        10'b0110000100: data <= 16'hffeb; 
        10'b0110000101: data <= 16'hffef; 
        10'b0110000110: data <= 16'h0017; 
        10'b0110000111: data <= 16'hffea; 
        10'b0110001000: data <= 16'hfff6; 
        10'b0110001001: data <= 16'h0013; 
        10'b0110001010: data <= 16'h0047; 
        10'b0110001011: data <= 16'h0059; 
        10'b0110001100: data <= 16'h0038; 
        10'b0110001101: data <= 16'h0041; 
        10'b0110001110: data <= 16'hffea; 
        10'b0110001111: data <= 16'hffd2; 
        10'b0110010000: data <= 16'hff9b; 
        10'b0110010001: data <= 16'hff14; 
        10'b0110010010: data <= 16'hfea5; 
        10'b0110010011: data <= 16'hfde8; 
        10'b0110010100: data <= 16'hfd51; 
        10'b0110010101: data <= 16'hfdbc; 
        10'b0110010110: data <= 16'hff2b; 
        10'b0110010111: data <= 16'h0005; 
        10'b0110011000: data <= 16'h002c; 
        10'b0110011001: data <= 16'h005c; 
        10'b0110011010: data <= 16'h0107; 
        10'b0110011011: data <= 16'h011a; 
        10'b0110011100: data <= 16'h00aa; 
        10'b0110011101: data <= 16'h006d; 
        10'b0110011110: data <= 16'h006d; 
        10'b0110011111: data <= 16'h005f; 
        10'b0110100000: data <= 16'h0020; 
        10'b0110100001: data <= 16'h000a; 
        10'b0110100010: data <= 16'hfff1; 
        10'b0110100011: data <= 16'hfff2; 
        10'b0110100100: data <= 16'h0017; 
        10'b0110100101: data <= 16'h0022; 
        10'b0110100110: data <= 16'h000c; 
        10'b0110100111: data <= 16'h0022; 
        10'b0110101000: data <= 16'h0022; 
        10'b0110101001: data <= 16'hffa1; 
        10'b0110101010: data <= 16'hffd6; 
        10'b0110101011: data <= 16'hffc5; 
        10'b0110101100: data <= 16'hff03; 
        10'b0110101101: data <= 16'hfecd; 
        10'b0110101110: data <= 16'hfe68; 
        10'b0110101111: data <= 16'hfe2c; 
        10'b0110110000: data <= 16'hfe02; 
        10'b0110110001: data <= 16'hfe88; 
        10'b0110110010: data <= 16'hff25; 
        10'b0110110011: data <= 16'h0007; 
        10'b0110110100: data <= 16'h0018; 
        10'b0110110101: data <= 16'h0165; 
        10'b0110110110: data <= 16'h01a2; 
        10'b0110110111: data <= 16'h0159; 
        10'b0110111000: data <= 16'h0132; 
        10'b0110111001: data <= 16'h0107; 
        10'b0110111010: data <= 16'h00aa; 
        10'b0110111011: data <= 16'h004d; 
        10'b0110111100: data <= 16'hfffd; 
        10'b0110111101: data <= 16'hffeb; 
        10'b0110111110: data <= 16'h0006; 
        10'b0110111111: data <= 16'h0025; 
        10'b0111000000: data <= 16'h0017; 
        10'b0111000001: data <= 16'h002d; 
        10'b0111000010: data <= 16'hfffc; 
        10'b0111000011: data <= 16'h0030; 
        10'b0111000100: data <= 16'h0025; 
        10'b0111000101: data <= 16'hffd5; 
        10'b0111000110: data <= 16'hffc4; 
        10'b0111000111: data <= 16'hfff7; 
        10'b0111001000: data <= 16'hff34; 
        10'b0111001001: data <= 16'hff1a; 
        10'b0111001010: data <= 16'hfe8e; 
        10'b0111001011: data <= 16'hfe48; 
        10'b0111001100: data <= 16'hfeec; 
        10'b0111001101: data <= 16'hff66; 
        10'b0111001110: data <= 16'hff20; 
        10'b0111001111: data <= 16'h0073; 
        10'b0111010000: data <= 16'h008b; 
        10'b0111010001: data <= 16'h012e; 
        10'b0111010010: data <= 16'h0103; 
        10'b0111010011: data <= 16'h010f; 
        10'b0111010100: data <= 16'h00d8; 
        10'b0111010101: data <= 16'h00a4; 
        10'b0111010110: data <= 16'h0020; 
        10'b0111010111: data <= 16'hffbc; 
        10'b0111011000: data <= 16'hffd6; 
        10'b0111011001: data <= 16'hffe8; 
        10'b0111011010: data <= 16'h001a; 
        10'b0111011011: data <= 16'h002d; 
        10'b0111011100: data <= 16'h0001; 
        10'b0111011101: data <= 16'h0006; 
        10'b0111011110: data <= 16'h001b; 
        10'b0111011111: data <= 16'hfffe; 
        10'b0111100000: data <= 16'h0009; 
        10'b0111100001: data <= 16'hffe5; 
        10'b0111100010: data <= 16'hff77; 
        10'b0111100011: data <= 16'hff4b; 
        10'b0111100100: data <= 16'hff1d; 
        10'b0111100101: data <= 16'hff45; 
        10'b0111100110: data <= 16'hff08; 
        10'b0111100111: data <= 16'hff48; 
        10'b0111101000: data <= 16'hffc5; 
        10'b0111101001: data <= 16'h002e; 
        10'b0111101010: data <= 16'h001a; 
        10'b0111101011: data <= 16'h002e; 
        10'b0111101100: data <= 16'hffe5; 
        10'b0111101101: data <= 16'h0049; 
        10'b0111101110: data <= 16'h0041; 
        10'b0111101111: data <= 16'h002e; 
        10'b0111110000: data <= 16'h0018; 
        10'b0111110001: data <= 16'hffda; 
        10'b0111110010: data <= 16'hffac; 
        10'b0111110011: data <= 16'hffda; 
        10'b0111110100: data <= 16'hffdf; 
        10'b0111110101: data <= 16'hffe6; 
        10'b0111110110: data <= 16'hfff2; 
        10'b0111110111: data <= 16'hfff4; 
        10'b0111111000: data <= 16'hfff3; 
        10'b0111111001: data <= 16'hfffc; 
        10'b0111111010: data <= 16'h001f; 
        10'b0111111011: data <= 16'h000a; 
        10'b0111111100: data <= 16'hffc8; 
        10'b0111111101: data <= 16'hff7c; 
        10'b0111111110: data <= 16'hff25; 
        10'b0111111111: data <= 16'hfef0; 
        10'b1000000000: data <= 16'hff03; 
        10'b1000000001: data <= 16'hff14; 
        10'b1000000010: data <= 16'hfed0; 
        10'b1000000011: data <= 16'hff98; 
        10'b1000000100: data <= 16'hffe0; 
        10'b1000000101: data <= 16'h0004; 
        10'b1000000110: data <= 16'h0055; 
        10'b1000000111: data <= 16'hffa6; 
        10'b1000001000: data <= 16'hff91; 
        10'b1000001001: data <= 16'hffc3; 
        10'b1000001010: data <= 16'hff74; 
        10'b1000001011: data <= 16'hffaa; 
        10'b1000001100: data <= 16'hff70; 
        10'b1000001101: data <= 16'hff23; 
        10'b1000001110: data <= 16'hff5e; 
        10'b1000001111: data <= 16'hff9a; 
        10'b1000010000: data <= 16'hffb0; 
        10'b1000010001: data <= 16'h0008; 
        10'b1000010010: data <= 16'hfff7; 
        10'b1000010011: data <= 16'h0002; 
        10'b1000010100: data <= 16'h002b; 
        10'b1000010101: data <= 16'h002e; 
        10'b1000010110: data <= 16'h002a; 
        10'b1000010111: data <= 16'h0015; 
        10'b1000011000: data <= 16'hffda; 
        10'b1000011001: data <= 16'hff54; 
        10'b1000011010: data <= 16'hfeed; 
        10'b1000011011: data <= 16'hfed9; 
        10'b1000011100: data <= 16'hfed1; 
        10'b1000011101: data <= 16'hfecf; 
        10'b1000011110: data <= 16'hff31; 
        10'b1000011111: data <= 16'hff6b; 
        10'b1000100000: data <= 16'hffa7; 
        10'b1000100001: data <= 16'h0027; 
        10'b1000100010: data <= 16'h0079; 
        10'b1000100011: data <= 16'hff82; 
        10'b1000100100: data <= 16'hff85; 
        10'b1000100101: data <= 16'hff65; 
        10'b1000100110: data <= 16'hff09; 
        10'b1000100111: data <= 16'hff16; 
        10'b1000101000: data <= 16'hfee0; 
        10'b1000101001: data <= 16'hfef6; 
        10'b1000101010: data <= 16'hff35; 
        10'b1000101011: data <= 16'hff74; 
        10'b1000101100: data <= 16'hffb9; 
        10'b1000101101: data <= 16'hffe6; 
        10'b1000101110: data <= 16'h002c; 
        10'b1000101111: data <= 16'hffec; 
        10'b1000110000: data <= 16'hffe9; 
        10'b1000110001: data <= 16'hfff6; 
        10'b1000110010: data <= 16'h0012; 
        10'b1000110011: data <= 16'hfff9; 
        10'b1000110100: data <= 16'hffd5; 
        10'b1000110101: data <= 16'hff7b; 
        10'b1000110110: data <= 16'hfeeb; 
        10'b1000110111: data <= 16'hfedf; 
        10'b1000111000: data <= 16'hfeef; 
        10'b1000111001: data <= 16'hfef5; 
        10'b1000111010: data <= 16'hff46; 
        10'b1000111011: data <= 16'hff40; 
        10'b1000111100: data <= 16'h000e; 
        10'b1000111101: data <= 16'h0013; 
        10'b1000111110: data <= 16'h0040; 
        10'b1000111111: data <= 16'hff57; 
        10'b1001000000: data <= 16'hff2d; 
        10'b1001000001: data <= 16'hfeec; 
        10'b1001000010: data <= 16'hfe83; 
        10'b1001000011: data <= 16'hff0d; 
        10'b1001000100: data <= 16'hfeb2; 
        10'b1001000101: data <= 16'hff01; 
        10'b1001000110: data <= 16'hff48; 
        10'b1001000111: data <= 16'hffb2; 
        10'b1001001000: data <= 16'hffcc; 
        10'b1001001001: data <= 16'h0028; 
        10'b1001001010: data <= 16'h0026; 
        10'b1001001011: data <= 16'h001a; 
        10'b1001001100: data <= 16'h0024; 
        10'b1001001101: data <= 16'h0025; 
        10'b1001001110: data <= 16'h0008; 
        10'b1001001111: data <= 16'hffcf; 
        10'b1001010000: data <= 16'hffe7; 
        10'b1001010001: data <= 16'hff8a; 
        10'b1001010010: data <= 16'hff75; 
        10'b1001010011: data <= 16'hff38; 
        10'b1001010100: data <= 16'hff4c; 
        10'b1001010101: data <= 16'hff95; 
        10'b1001010110: data <= 16'hff68; 
        10'b1001010111: data <= 16'hff84; 
        10'b1001011000: data <= 16'hffc8; 
        10'b1001011001: data <= 16'h0008; 
        10'b1001011010: data <= 16'hffdf; 
        10'b1001011011: data <= 16'hff8e; 
        10'b1001011100: data <= 16'hff7d; 
        10'b1001011101: data <= 16'hfef0; 
        10'b1001011110: data <= 16'hfef1; 
        10'b1001011111: data <= 16'hfef0; 
        10'b1001100000: data <= 16'hfee2; 
        10'b1001100001: data <= 16'hff0e; 
        10'b1001100010: data <= 16'hff72; 
        10'b1001100011: data <= 16'hff94; 
        10'b1001100100: data <= 16'hfffb; 
        10'b1001100101: data <= 16'h0011; 
        10'b1001100110: data <= 16'h0024; 
        10'b1001100111: data <= 16'hfff8; 
        10'b1001101000: data <= 16'h000c; 
        10'b1001101001: data <= 16'h0003; 
        10'b1001101010: data <= 16'h000a; 
        10'b1001101011: data <= 16'hffe2; 
        10'b1001101100: data <= 16'hfff2; 
        10'b1001101101: data <= 16'h0012; 
        10'b1001101110: data <= 16'hffd5; 
        10'b1001101111: data <= 16'h0016; 
        10'b1001110000: data <= 16'h0022; 
        10'b1001110001: data <= 16'hffc9; 
        10'b1001110010: data <= 16'hff98; 
        10'b1001110011: data <= 16'hff4e; 
        10'b1001110100: data <= 16'hff5a; 
        10'b1001110101: data <= 16'hffbd; 
        10'b1001110110: data <= 16'h0014; 
        10'b1001110111: data <= 16'h0014; 
        10'b1001111000: data <= 16'hff99; 
        10'b1001111001: data <= 16'hff80; 
        10'b1001111010: data <= 16'hff26; 
        10'b1001111011: data <= 16'hff26; 
        10'b1001111100: data <= 16'hff0a; 
        10'b1001111101: data <= 16'hff29; 
        10'b1001111110: data <= 16'hff93; 
        10'b1001111111: data <= 16'hffdb; 
        10'b1010000000: data <= 16'h0018; 
        10'b1010000001: data <= 16'hffe9; 
        10'b1010000010: data <= 16'h000b; 
        10'b1010000011: data <= 16'h0001; 
        10'b1010000100: data <= 16'h0011; 
        10'b1010000101: data <= 16'h0022; 
        10'b1010000110: data <= 16'hffe6; 
        10'b1010000111: data <= 16'hffe8; 
        10'b1010001000: data <= 16'h002d; 
        10'b1010001001: data <= 16'h003c; 
        10'b1010001010: data <= 16'h0083; 
        10'b1010001011: data <= 16'h00af; 
        10'b1010001100: data <= 16'h0054; 
        10'b1010001101: data <= 16'h0011; 
        10'b1010001110: data <= 16'hffcd; 
        10'b1010001111: data <= 16'hff89; 
        10'b1010010000: data <= 16'hff9f; 
        10'b1010010001: data <= 16'h0007; 
        10'b1010010010: data <= 16'h0044; 
        10'b1010010011: data <= 16'h003f; 
        10'b1010010100: data <= 16'hffe6; 
        10'b1010010101: data <= 16'hffd9; 
        10'b1010010110: data <= 16'hff74; 
        10'b1010010111: data <= 16'hff3d; 
        10'b1010011000: data <= 16'hff39; 
        10'b1010011001: data <= 16'hff64; 
        10'b1010011010: data <= 16'hff80; 
        10'b1010011011: data <= 16'hffac; 
        10'b1010011100: data <= 16'hffdb; 
        10'b1010011101: data <= 16'h0003; 
        10'b1010011110: data <= 16'h0002; 
        10'b1010011111: data <= 16'hfff2; 
        10'b1010100000: data <= 16'h0000; 
        10'b1010100001: data <= 16'hfffb; 
        10'b1010100010: data <= 16'h000c; 
        10'b1010100011: data <= 16'h001d; 
        10'b1010100100: data <= 16'h003f; 
        10'b1010100101: data <= 16'h0090; 
        10'b1010100110: data <= 16'h00da; 
        10'b1010100111: data <= 16'h00f6; 
        10'b1010101000: data <= 16'h00d1; 
        10'b1010101001: data <= 16'h006c; 
        10'b1010101010: data <= 16'h00e8; 
        10'b1010101011: data <= 16'h0089; 
        10'b1010101100: data <= 16'h0077; 
        10'b1010101101: data <= 16'h00a7; 
        10'b1010101110: data <= 16'h0067; 
        10'b1010101111: data <= 16'h0094; 
        10'b1010110000: data <= 16'h0058; 
        10'b1010110001: data <= 16'h0045; 
        10'b1010110010: data <= 16'hfffc; 
        10'b1010110011: data <= 16'hffc0; 
        10'b1010110100: data <= 16'hffbc; 
        10'b1010110101: data <= 16'hffad; 
        10'b1010110110: data <= 16'hffa3; 
        10'b1010110111: data <= 16'hffab; 
        10'b1010111000: data <= 16'h000d; 
        10'b1010111001: data <= 16'hfff9; 
        10'b1010111010: data <= 16'hffea; 
        10'b1010111011: data <= 16'h0019; 
        10'b1010111100: data <= 16'hffe9; 
        10'b1010111101: data <= 16'h0015; 
        10'b1010111110: data <= 16'h0026; 
        10'b1010111111: data <= 16'h0023; 
        10'b1011000000: data <= 16'h0014; 
        10'b1011000001: data <= 16'h0048; 
        10'b1011000010: data <= 16'h006a; 
        10'b1011000011: data <= 16'h00a4; 
        10'b1011000100: data <= 16'h00fe; 
        10'b1011000101: data <= 16'h00f8; 
        10'b1011000110: data <= 16'h0125; 
        10'b1011000111: data <= 16'h0111; 
        10'b1011001000: data <= 16'h00f3; 
        10'b1011001001: data <= 16'h00c1; 
        10'b1011001010: data <= 16'h00c5; 
        10'b1011001011: data <= 16'h00d1; 
        10'b1011001100: data <= 16'h00af; 
        10'b1011001101: data <= 16'h00a3; 
        10'b1011001110: data <= 16'h0084; 
        10'b1011001111: data <= 16'h002d; 
        10'b1011010000: data <= 16'hffc9; 
        10'b1011010001: data <= 16'h0007; 
        10'b1011010010: data <= 16'hffe5; 
        10'b1011010011: data <= 16'hffec; 
        10'b1011010100: data <= 16'hfffa; 
        10'b1011010101: data <= 16'h000d; 
        10'b1011010110: data <= 16'h0032; 
        10'b1011010111: data <= 16'h0020; 
        10'b1011011000: data <= 16'hffee; 
        10'b1011011001: data <= 16'h000a; 
        10'b1011011010: data <= 16'h002f; 
        10'b1011011011: data <= 16'hfff8; 
        10'b1011011100: data <= 16'hfff0; 
        10'b1011011101: data <= 16'h002c; 
        10'b1011011110: data <= 16'h0003; 
        10'b1011011111: data <= 16'h0028; 
        10'b1011100000: data <= 16'h0026; 
        10'b1011100001: data <= 16'h0005; 
        10'b1011100010: data <= 16'h0037; 
        10'b1011100011: data <= 16'h0051; 
        10'b1011100100: data <= 16'h0017; 
        10'b1011100101: data <= 16'h0046; 
        10'b1011100110: data <= 16'h0096; 
        10'b1011100111: data <= 16'h00b9; 
        10'b1011101000: data <= 16'h0092; 
        10'b1011101001: data <= 16'h00bb; 
        10'b1011101010: data <= 16'h006b; 
        10'b1011101011: data <= 16'h0032; 
        10'b1011101100: data <= 16'h0002; 
        10'b1011101101: data <= 16'h0013; 
        10'b1011101110: data <= 16'hfffb; 
        10'b1011101111: data <= 16'h000b; 
        10'b1011110000: data <= 16'h0002; 
        10'b1011110001: data <= 16'hfff3; 
        10'b1011110010: data <= 16'hfffd; 
        10'b1011110011: data <= 16'hfffa; 
        10'b1011110100: data <= 16'hffe9; 
        10'b1011110101: data <= 16'h0013; 
        10'b1011110110: data <= 16'h000d; 
        10'b1011110111: data <= 16'h0018; 
        10'b1011111000: data <= 16'h0020; 
        10'b1011111001: data <= 16'h0013; 
        10'b1011111010: data <= 16'h0008; 
        10'b1011111011: data <= 16'h0003; 
        10'b1011111100: data <= 16'h0035; 
        10'b1011111101: data <= 16'h0020; 
        10'b1011111110: data <= 16'h000a; 
        10'b1011111111: data <= 16'h0021; 
        10'b1100000000: data <= 16'h0010; 
        10'b1100000001: data <= 16'h003d; 
        10'b1100000010: data <= 16'h0024; 
        10'b1100000011: data <= 16'h001c; 
        10'b1100000100: data <= 16'h0054; 
        10'b1100000101: data <= 16'h001d; 
        10'b1100000110: data <= 16'h0019; 
        10'b1100000111: data <= 16'h003b; 
        10'b1100001000: data <= 16'h0007; 
        10'b1100001001: data <= 16'hfff6; 
        10'b1100001010: data <= 16'h0030; 
        10'b1100001011: data <= 16'h001a; 
        10'b1100001100: data <= 16'h000c; 
        10'b1100001101: data <= 16'hfff7; 
        10'b1100001110: data <= 16'hffec; 
        10'b1100001111: data <= 16'h0020; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 11) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 17'h00006; 
        10'b0000000001: data <= 17'h00008; 
        10'b0000000010: data <= 17'h0003d; 
        10'b0000000011: data <= 17'h00017; 
        10'b0000000100: data <= 17'h00063; 
        10'b0000000101: data <= 17'h1ffd4; 
        10'b0000000110: data <= 17'h1ffe3; 
        10'b0000000111: data <= 17'h00020; 
        10'b0000001000: data <= 17'h0004c; 
        10'b0000001001: data <= 17'h0004b; 
        10'b0000001010: data <= 17'h1ffd6; 
        10'b0000001011: data <= 17'h00014; 
        10'b0000001100: data <= 17'h00015; 
        10'b0000001101: data <= 17'h1fff5; 
        10'b0000001110: data <= 17'h00050; 
        10'b0000001111: data <= 17'h00015; 
        10'b0000010000: data <= 17'h00002; 
        10'b0000010001: data <= 17'h1fffd; 
        10'b0000010010: data <= 17'h00008; 
        10'b0000010011: data <= 17'h0001c; 
        10'b0000010100: data <= 17'h00033; 
        10'b0000010101: data <= 17'h00061; 
        10'b0000010110: data <= 17'h1ffe6; 
        10'b0000010111: data <= 17'h00047; 
        10'b0000011000: data <= 17'h1fff6; 
        10'b0000011001: data <= 17'h00033; 
        10'b0000011010: data <= 17'h1fffc; 
        10'b0000011011: data <= 17'h00000; 
        10'b0000011100: data <= 17'h0005b; 
        10'b0000011101: data <= 17'h1ffec; 
        10'b0000011110: data <= 17'h00015; 
        10'b0000011111: data <= 17'h0005a; 
        10'b0000100000: data <= 17'h00023; 
        10'b0000100001: data <= 17'h00003; 
        10'b0000100010: data <= 17'h00059; 
        10'b0000100011: data <= 17'h0001c; 
        10'b0000100100: data <= 17'h00009; 
        10'b0000100101: data <= 17'h1fff1; 
        10'b0000100110: data <= 17'h1fff4; 
        10'b0000100111: data <= 17'h1ffd1; 
        10'b0000101000: data <= 17'h0004d; 
        10'b0000101001: data <= 17'h1fffa; 
        10'b0000101010: data <= 17'h0005c; 
        10'b0000101011: data <= 17'h1ffe8; 
        10'b0000101100: data <= 17'h00028; 
        10'b0000101101: data <= 17'h00045; 
        10'b0000101110: data <= 17'h0004e; 
        10'b0000101111: data <= 17'h0003e; 
        10'b0000110000: data <= 17'h00002; 
        10'b0000110001: data <= 17'h0003d; 
        10'b0000110010: data <= 17'h1fffe; 
        10'b0000110011: data <= 17'h00061; 
        10'b0000110100: data <= 17'h0004b; 
        10'b0000110101: data <= 17'h1ffe5; 
        10'b0000110110: data <= 17'h1ffe6; 
        10'b0000110111: data <= 17'h00028; 
        10'b0000111000: data <= 17'h00056; 
        10'b0000111001: data <= 17'h00055; 
        10'b0000111010: data <= 17'h00043; 
        10'b0000111011: data <= 17'h1fff4; 
        10'b0000111100: data <= 17'h0004e; 
        10'b0000111101: data <= 17'h1ffdb; 
        10'b0000111110: data <= 17'h1ffe2; 
        10'b0000111111: data <= 17'h0003d; 
        10'b0001000000: data <= 17'h00033; 
        10'b0001000001: data <= 17'h1ffe2; 
        10'b0001000010: data <= 17'h1fff9; 
        10'b0001000011: data <= 17'h00026; 
        10'b0001000100: data <= 17'h1fff5; 
        10'b0001000101: data <= 17'h1ffec; 
        10'b0001000110: data <= 17'h00018; 
        10'b0001000111: data <= 17'h0004e; 
        10'b0001001000: data <= 17'h0003f; 
        10'b0001001001: data <= 17'h0000c; 
        10'b0001001010: data <= 17'h0001f; 
        10'b0001001011: data <= 17'h00058; 
        10'b0001001100: data <= 17'h0004b; 
        10'b0001001101: data <= 17'h00057; 
        10'b0001001110: data <= 17'h1ffd4; 
        10'b0001001111: data <= 17'h00044; 
        10'b0001010000: data <= 17'h0001a; 
        10'b0001010001: data <= 17'h0003c; 
        10'b0001010010: data <= 17'h00033; 
        10'b0001010011: data <= 17'h0004c; 
        10'b0001010100: data <= 17'h1fff9; 
        10'b0001010101: data <= 17'h00005; 
        10'b0001010110: data <= 17'h0004f; 
        10'b0001010111: data <= 17'h1fff4; 
        10'b0001011000: data <= 17'h00009; 
        10'b0001011001: data <= 17'h1fffb; 
        10'b0001011010: data <= 17'h1ffe3; 
        10'b0001011011: data <= 17'h00033; 
        10'b0001011100: data <= 17'h00000; 
        10'b0001011101: data <= 17'h00034; 
        10'b0001011110: data <= 17'h1ffd6; 
        10'b0001011111: data <= 17'h0000a; 
        10'b0001100000: data <= 17'h00029; 
        10'b0001100001: data <= 17'h1ffc7; 
        10'b0001100010: data <= 17'h0002f; 
        10'b0001100011: data <= 17'h1ffd9; 
        10'b0001100100: data <= 17'h1ffac; 
        10'b0001100101: data <= 17'h1ffbb; 
        10'b0001100110: data <= 17'h1ffc5; 
        10'b0001100111: data <= 17'h1ffd8; 
        10'b0001101000: data <= 17'h1fff6; 
        10'b0001101001: data <= 17'h1ffdc; 
        10'b0001101010: data <= 17'h00020; 
        10'b0001101011: data <= 17'h1fffc; 
        10'b0001101100: data <= 17'h00026; 
        10'b0001101101: data <= 17'h00062; 
        10'b0001101110: data <= 17'h1ffe0; 
        10'b0001101111: data <= 17'h00028; 
        10'b0001110000: data <= 17'h0005f; 
        10'b0001110001: data <= 17'h1ffde; 
        10'b0001110010: data <= 17'h00035; 
        10'b0001110011: data <= 17'h1ffd8; 
        10'b0001110100: data <= 17'h00016; 
        10'b0001110101: data <= 17'h1ffee; 
        10'b0001110110: data <= 17'h00004; 
        10'b0001110111: data <= 17'h1ffd9; 
        10'b0001111000: data <= 17'h0001d; 
        10'b0001111001: data <= 17'h1fff2; 
        10'b0001111010: data <= 17'h1ffa3; 
        10'b0001111011: data <= 17'h1ff4d; 
        10'b0001111100: data <= 17'h1ff44; 
        10'b0001111101: data <= 17'h1ff4d; 
        10'b0001111110: data <= 17'h1ff2b; 
        10'b0001111111: data <= 17'h1fea1; 
        10'b0010000000: data <= 17'h1ff31; 
        10'b0010000001: data <= 17'h1ff64; 
        10'b0010000010: data <= 17'h1ff78; 
        10'b0010000011: data <= 17'h1ffdb; 
        10'b0010000100: data <= 17'h1ff9b; 
        10'b0010000101: data <= 17'h0002f; 
        10'b0010000110: data <= 17'h00007; 
        10'b0010000111: data <= 17'h1ffcf; 
        10'b0010001000: data <= 17'h0005a; 
        10'b0010001001: data <= 17'h1fffd; 
        10'b0010001010: data <= 17'h00058; 
        10'b0010001011: data <= 17'h00055; 
        10'b0010001100: data <= 17'h00051; 
        10'b0010001101: data <= 17'h00003; 
        10'b0010001110: data <= 17'h0004e; 
        10'b0010001111: data <= 17'h1ffeb; 
        10'b0010010000: data <= 17'h1ffc3; 
        10'b0010010001: data <= 17'h1fff6; 
        10'b0010010010: data <= 17'h1ffd1; 
        10'b0010010011: data <= 17'h1ffef; 
        10'b0010010100: data <= 17'h1ffc9; 
        10'b0010010101: data <= 17'h1ff80; 
        10'b0010010110: data <= 17'h1fec5; 
        10'b0010010111: data <= 17'h1fe7e; 
        10'b0010011000: data <= 17'h1fe1a; 
        10'b0010011001: data <= 17'h1fdc6; 
        10'b0010011010: data <= 17'h1fd39; 
        10'b0010011011: data <= 17'h1fd3e; 
        10'b0010011100: data <= 17'h1fd1c; 
        10'b0010011101: data <= 17'h1fd73; 
        10'b0010011110: data <= 17'h1fdd7; 
        10'b0010011111: data <= 17'h1fe5b; 
        10'b0010100000: data <= 17'h1fed5; 
        10'b0010100001: data <= 17'h1ff95; 
        10'b0010100010: data <= 17'h1ff5b; 
        10'b0010100011: data <= 17'h1ffeb; 
        10'b0010100100: data <= 17'h00048; 
        10'b0010100101: data <= 17'h0003a; 
        10'b0010100110: data <= 17'h1fff1; 
        10'b0010100111: data <= 17'h00003; 
        10'b0010101000: data <= 17'h00043; 
        10'b0010101001: data <= 17'h0005c; 
        10'b0010101010: data <= 17'h00006; 
        10'b0010101011: data <= 17'h0000f; 
        10'b0010101100: data <= 17'h00063; 
        10'b0010101101: data <= 17'h00076; 
        10'b0010101110: data <= 17'h0008a; 
        10'b0010101111: data <= 17'h000d0; 
        10'b0010110000: data <= 17'h00135; 
        10'b0010110001: data <= 17'h000f8; 
        10'b0010110010: data <= 17'h00107; 
        10'b0010110011: data <= 17'h0002f; 
        10'b0010110100: data <= 17'h1ff2d; 
        10'b0010110101: data <= 17'h1fe45; 
        10'b0010110110: data <= 17'h1fe31; 
        10'b0010110111: data <= 17'h1ff10; 
        10'b0010111000: data <= 17'h1ff6e; 
        10'b0010111001: data <= 17'h1ff53; 
        10'b0010111010: data <= 17'h1ff2e; 
        10'b0010111011: data <= 17'h1ff0d; 
        10'b0010111100: data <= 17'h1fe90; 
        10'b0010111101: data <= 17'h1ff76; 
        10'b0010111110: data <= 17'h1fefe; 
        10'b0010111111: data <= 17'h1ff44; 
        10'b0011000000: data <= 17'h1ff82; 
        10'b0011000001: data <= 17'h1ffd6; 
        10'b0011000010: data <= 17'h1ffd4; 
        10'b0011000011: data <= 17'h0000a; 
        10'b0011000100: data <= 17'h0003d; 
        10'b0011000101: data <= 17'h0005d; 
        10'b0011000110: data <= 17'h0004c; 
        10'b0011000111: data <= 17'h000b4; 
        10'b0011001000: data <= 17'h000da; 
        10'b0011001001: data <= 17'h000c4; 
        10'b0011001010: data <= 17'h0011c; 
        10'b0011001011: data <= 17'h001b3; 
        10'b0011001100: data <= 17'h00253; 
        10'b0011001101: data <= 17'h001d8; 
        10'b0011001110: data <= 17'h00145; 
        10'b0011001111: data <= 17'h00166; 
        10'b0011010000: data <= 17'h0017e; 
        10'b0011010001: data <= 17'h00049; 
        10'b0011010010: data <= 17'h00036; 
        10'b0011010011: data <= 17'h00089; 
        10'b0011010100: data <= 17'h00193; 
        10'b0011010101: data <= 17'h001c0; 
        10'b0011010110: data <= 17'h00130; 
        10'b0011010111: data <= 17'h000f3; 
        10'b0011011000: data <= 17'h0003b; 
        10'b0011011001: data <= 17'h1ffbd; 
        10'b0011011010: data <= 17'h00020; 
        10'b0011011011: data <= 17'h1ffb7; 
        10'b0011011100: data <= 17'h1ffbc; 
        10'b0011011101: data <= 17'h1fffc; 
        10'b0011011110: data <= 17'h00030; 
        10'b0011011111: data <= 17'h1ffee; 
        10'b0011100000: data <= 17'h1ffd1; 
        10'b0011100001: data <= 17'h00061; 
        10'b0011100010: data <= 17'h00025; 
        10'b0011100011: data <= 17'h00098; 
        10'b0011100100: data <= 17'h00134; 
        10'b0011100101: data <= 17'h00116; 
        10'b0011100110: data <= 17'h00174; 
        10'b0011100111: data <= 17'h0029b; 
        10'b0011101000: data <= 17'h001c1; 
        10'b0011101001: data <= 17'h00135; 
        10'b0011101010: data <= 17'h0018a; 
        10'b0011101011: data <= 17'h0020f; 
        10'b0011101100: data <= 17'h001f5; 
        10'b0011101101: data <= 17'h000fc; 
        10'b0011101110: data <= 17'h00093; 
        10'b0011101111: data <= 17'h000cd; 
        10'b0011110000: data <= 17'h00163; 
        10'b0011110001: data <= 17'h00222; 
        10'b0011110010: data <= 17'h00176; 
        10'b0011110011: data <= 17'h00141; 
        10'b0011110100: data <= 17'h00100; 
        10'b0011110101: data <= 17'h00006; 
        10'b0011110110: data <= 17'h0009b; 
        10'b0011110111: data <= 17'h00084; 
        10'b0011111000: data <= 17'h1ffa2; 
        10'b0011111001: data <= 17'h1ffd3; 
        10'b0011111010: data <= 17'h00034; 
        10'b0011111011: data <= 17'h00050; 
        10'b0011111100: data <= 17'h00029; 
        10'b0011111101: data <= 17'h0004d; 
        10'b0011111110: data <= 17'h00068; 
        10'b0011111111: data <= 17'h000db; 
        10'b0100000000: data <= 17'h0012e; 
        10'b0100000001: data <= 17'h00157; 
        10'b0100000010: data <= 17'h0007e; 
        10'b0100000011: data <= 17'h000a7; 
        10'b0100000100: data <= 17'h000be; 
        10'b0100000101: data <= 17'h0007d; 
        10'b0100000110: data <= 17'h00133; 
        10'b0100000111: data <= 17'h00178; 
        10'b0100001000: data <= 17'h001e0; 
        10'b0100001001: data <= 17'h00186; 
        10'b0100001010: data <= 17'h0022f; 
        10'b0100001011: data <= 17'h002b0; 
        10'b0100001100: data <= 17'h0027a; 
        10'b0100001101: data <= 17'h002c4; 
        10'b0100001110: data <= 17'h001ce; 
        10'b0100001111: data <= 17'h001d7; 
        10'b0100010000: data <= 17'h0018c; 
        10'b0100010001: data <= 17'h0014a; 
        10'b0100010010: data <= 17'h0009c; 
        10'b0100010011: data <= 17'h1ffc7; 
        10'b0100010100: data <= 17'h1ffa0; 
        10'b0100010101: data <= 17'h1ffd1; 
        10'b0100010110: data <= 17'h0002a; 
        10'b0100010111: data <= 17'h1ffeb; 
        10'b0100011000: data <= 17'h00010; 
        10'b0100011001: data <= 17'h00054; 
        10'b0100011010: data <= 17'h0005d; 
        10'b0100011011: data <= 17'h00111; 
        10'b0100011100: data <= 17'h00138; 
        10'b0100011101: data <= 17'h00104; 
        10'b0100011110: data <= 17'h00030; 
        10'b0100011111: data <= 17'h0004e; 
        10'b0100100000: data <= 17'h1ff97; 
        10'b0100100001: data <= 17'h1fffc; 
        10'b0100100010: data <= 17'h000bf; 
        10'b0100100011: data <= 17'h0014f; 
        10'b0100100100: data <= 17'h000e9; 
        10'b0100100101: data <= 17'h0021f; 
        10'b0100100110: data <= 17'h002bb; 
        10'b0100100111: data <= 17'h0035a; 
        10'b0100101000: data <= 17'h003d1; 
        10'b0100101001: data <= 17'h002d4; 
        10'b0100101010: data <= 17'h0023a; 
        10'b0100101011: data <= 17'h00251; 
        10'b0100101100: data <= 17'h00209; 
        10'b0100101101: data <= 17'h001bb; 
        10'b0100101110: data <= 17'h000c4; 
        10'b0100101111: data <= 17'h1ffb0; 
        10'b0100110000: data <= 17'h1ff7c; 
        10'b0100110001: data <= 17'h1ffca; 
        10'b0100110010: data <= 17'h0000a; 
        10'b0100110011: data <= 17'h1ffec; 
        10'b0100110100: data <= 17'h0004a; 
        10'b0100110101: data <= 17'h00034; 
        10'b0100110110: data <= 17'h0005e; 
        10'b0100110111: data <= 17'h00117; 
        10'b0100111000: data <= 17'h00150; 
        10'b0100111001: data <= 17'h000a7; 
        10'b0100111010: data <= 17'h0003d; 
        10'b0100111011: data <= 17'h00036; 
        10'b0100111100: data <= 17'h00010; 
        10'b0100111101: data <= 17'h000ca; 
        10'b0100111110: data <= 17'h00068; 
        10'b0100111111: data <= 17'h00083; 
        10'b0101000000: data <= 17'h000d9; 
        10'b0101000001: data <= 17'h000d7; 
        10'b0101000010: data <= 17'h000e0; 
        10'b0101000011: data <= 17'h00291; 
        10'b0101000100: data <= 17'h00355; 
        10'b0101000101: data <= 17'h00238; 
        10'b0101000110: data <= 17'h0023e; 
        10'b0101000111: data <= 17'h001b9; 
        10'b0101001000: data <= 17'h001ad; 
        10'b0101001001: data <= 17'h0010e; 
        10'b0101001010: data <= 17'h000c3; 
        10'b0101001011: data <= 17'h1ffbc; 
        10'b0101001100: data <= 17'h1ff3b; 
        10'b0101001101: data <= 17'h1fffa; 
        10'b0101001110: data <= 17'h00013; 
        10'b0101001111: data <= 17'h00056; 
        10'b0101010000: data <= 17'h00042; 
        10'b0101010001: data <= 17'h1fffb; 
        10'b0101010010: data <= 17'h0002f; 
        10'b0101010011: data <= 17'h000b0; 
        10'b0101010100: data <= 17'h000c5; 
        10'b0101010101: data <= 17'h00020; 
        10'b0101010110: data <= 17'h0002c; 
        10'b0101010111: data <= 17'h000bc; 
        10'b0101011000: data <= 17'h00081; 
        10'b0101011001: data <= 17'h1fff9; 
        10'b0101011010: data <= 17'h1ff66; 
        10'b0101011011: data <= 17'h1fe67; 
        10'b0101011100: data <= 17'h1fc9f; 
        10'b0101011101: data <= 17'h1fac6; 
        10'b0101011110: data <= 17'h1fc16; 
        10'b0101011111: data <= 17'h00016; 
        10'b0101100000: data <= 17'h00236; 
        10'b0101100001: data <= 17'h00201; 
        10'b0101100010: data <= 17'h000ca; 
        10'b0101100011: data <= 17'h00049; 
        10'b0101100100: data <= 17'h0000e; 
        10'b0101100101: data <= 17'h1ffb6; 
        10'b0101100110: data <= 17'h1ffbd; 
        10'b0101100111: data <= 17'h1ff87; 
        10'b0101101000: data <= 17'h1ffa9; 
        10'b0101101001: data <= 17'h00052; 
        10'b0101101010: data <= 17'h00039; 
        10'b0101101011: data <= 17'h00001; 
        10'b0101101100: data <= 17'h00047; 
        10'b0101101101: data <= 17'h0002a; 
        10'b0101101110: data <= 17'h0004d; 
        10'b0101101111: data <= 17'h000a0; 
        10'b0101110000: data <= 17'h0003b; 
        10'b0101110001: data <= 17'h00019; 
        10'b0101110010: data <= 17'h1ffcc; 
        10'b0101110011: data <= 17'h00022; 
        10'b0101110100: data <= 17'h1ffe8; 
        10'b0101110101: data <= 17'h1ff7d; 
        10'b0101110110: data <= 17'h1fe53; 
        10'b0101110111: data <= 17'h1fc77; 
        10'b0101111000: data <= 17'h1f9cc; 
        10'b0101111001: data <= 17'h1f912; 
        10'b0101111010: data <= 17'h1fc4b; 
        10'b0101111011: data <= 17'h1ff84; 
        10'b0101111100: data <= 17'h00121; 
        10'b0101111101: data <= 17'h000ba; 
        10'b0101111110: data <= 17'h00028; 
        10'b0101111111: data <= 17'h00055; 
        10'b0110000000: data <= 17'h1ff52; 
        10'b0110000001: data <= 17'h1ff21; 
        10'b0110000010: data <= 17'h1ffcc; 
        10'b0110000011: data <= 17'h00010; 
        10'b0110000100: data <= 17'h1ffd6; 
        10'b0110000101: data <= 17'h1ffde; 
        10'b0110000110: data <= 17'h0002d; 
        10'b0110000111: data <= 17'h1ffd4; 
        10'b0110001000: data <= 17'h1ffed; 
        10'b0110001001: data <= 17'h00026; 
        10'b0110001010: data <= 17'h0008f; 
        10'b0110001011: data <= 17'h000b2; 
        10'b0110001100: data <= 17'h00071; 
        10'b0110001101: data <= 17'h00083; 
        10'b0110001110: data <= 17'h1ffd5; 
        10'b0110001111: data <= 17'h1ffa5; 
        10'b0110010000: data <= 17'h1ff37; 
        10'b0110010001: data <= 17'h1fe28; 
        10'b0110010010: data <= 17'h1fd4b; 
        10'b0110010011: data <= 17'h1fbd0; 
        10'b0110010100: data <= 17'h1faa1; 
        10'b0110010101: data <= 17'h1fb78; 
        10'b0110010110: data <= 17'h1fe57; 
        10'b0110010111: data <= 17'h0000a; 
        10'b0110011000: data <= 17'h00058; 
        10'b0110011001: data <= 17'h000b7; 
        10'b0110011010: data <= 17'h0020d; 
        10'b0110011011: data <= 17'h00235; 
        10'b0110011100: data <= 17'h00154; 
        10'b0110011101: data <= 17'h000d9; 
        10'b0110011110: data <= 17'h000da; 
        10'b0110011111: data <= 17'h000bd; 
        10'b0110100000: data <= 17'h00040; 
        10'b0110100001: data <= 17'h00013; 
        10'b0110100010: data <= 17'h1ffe2; 
        10'b0110100011: data <= 17'h1ffe5; 
        10'b0110100100: data <= 17'h0002e; 
        10'b0110100101: data <= 17'h00044; 
        10'b0110100110: data <= 17'h00019; 
        10'b0110100111: data <= 17'h00043; 
        10'b0110101000: data <= 17'h00043; 
        10'b0110101001: data <= 17'h1ff42; 
        10'b0110101010: data <= 17'h1ffab; 
        10'b0110101011: data <= 17'h1ff8a; 
        10'b0110101100: data <= 17'h1fe06; 
        10'b0110101101: data <= 17'h1fd9a; 
        10'b0110101110: data <= 17'h1fccf; 
        10'b0110101111: data <= 17'h1fc58; 
        10'b0110110000: data <= 17'h1fc05; 
        10'b0110110001: data <= 17'h1fd11; 
        10'b0110110010: data <= 17'h1fe49; 
        10'b0110110011: data <= 17'h0000d; 
        10'b0110110100: data <= 17'h00030; 
        10'b0110110101: data <= 17'h002cb; 
        10'b0110110110: data <= 17'h00345; 
        10'b0110110111: data <= 17'h002b2; 
        10'b0110111000: data <= 17'h00264; 
        10'b0110111001: data <= 17'h0020f; 
        10'b0110111010: data <= 17'h00154; 
        10'b0110111011: data <= 17'h0009a; 
        10'b0110111100: data <= 17'h1fffa; 
        10'b0110111101: data <= 17'h1ffd6; 
        10'b0110111110: data <= 17'h0000b; 
        10'b0110111111: data <= 17'h00049; 
        10'b0111000000: data <= 17'h0002e; 
        10'b0111000001: data <= 17'h0005b; 
        10'b0111000010: data <= 17'h1fff9; 
        10'b0111000011: data <= 17'h0005f; 
        10'b0111000100: data <= 17'h0004b; 
        10'b0111000101: data <= 17'h1ffab; 
        10'b0111000110: data <= 17'h1ff88; 
        10'b0111000111: data <= 17'h1ffef; 
        10'b0111001000: data <= 17'h1fe69; 
        10'b0111001001: data <= 17'h1fe34; 
        10'b0111001010: data <= 17'h1fd1b; 
        10'b0111001011: data <= 17'h1fc90; 
        10'b0111001100: data <= 17'h1fdd8; 
        10'b0111001101: data <= 17'h1fecb; 
        10'b0111001110: data <= 17'h1fe40; 
        10'b0111001111: data <= 17'h000e6; 
        10'b0111010000: data <= 17'h00117; 
        10'b0111010001: data <= 17'h0025d; 
        10'b0111010010: data <= 17'h00206; 
        10'b0111010011: data <= 17'h0021f; 
        10'b0111010100: data <= 17'h001b0; 
        10'b0111010101: data <= 17'h00149; 
        10'b0111010110: data <= 17'h00041; 
        10'b0111010111: data <= 17'h1ff79; 
        10'b0111011000: data <= 17'h1ffac; 
        10'b0111011001: data <= 17'h1ffd0; 
        10'b0111011010: data <= 17'h00033; 
        10'b0111011011: data <= 17'h00059; 
        10'b0111011100: data <= 17'h00003; 
        10'b0111011101: data <= 17'h0000c; 
        10'b0111011110: data <= 17'h00037; 
        10'b0111011111: data <= 17'h1fffc; 
        10'b0111100000: data <= 17'h00012; 
        10'b0111100001: data <= 17'h1ffca; 
        10'b0111100010: data <= 17'h1feed; 
        10'b0111100011: data <= 17'h1fe96; 
        10'b0111100100: data <= 17'h1fe3a; 
        10'b0111100101: data <= 17'h1fe89; 
        10'b0111100110: data <= 17'h1fe0f; 
        10'b0111100111: data <= 17'h1fe8f; 
        10'b0111101000: data <= 17'h1ff8a; 
        10'b0111101001: data <= 17'h0005c; 
        10'b0111101010: data <= 17'h00034; 
        10'b0111101011: data <= 17'h0005c; 
        10'b0111101100: data <= 17'h1ffca; 
        10'b0111101101: data <= 17'h00091; 
        10'b0111101110: data <= 17'h00082; 
        10'b0111101111: data <= 17'h0005c; 
        10'b0111110000: data <= 17'h00031; 
        10'b0111110001: data <= 17'h1ffb5; 
        10'b0111110010: data <= 17'h1ff59; 
        10'b0111110011: data <= 17'h1ffb5; 
        10'b0111110100: data <= 17'h1ffbf; 
        10'b0111110101: data <= 17'h1ffcd; 
        10'b0111110110: data <= 17'h1ffe4; 
        10'b0111110111: data <= 17'h1ffe7; 
        10'b0111111000: data <= 17'h1ffe7; 
        10'b0111111001: data <= 17'h1fff8; 
        10'b0111111010: data <= 17'h0003e; 
        10'b0111111011: data <= 17'h00013; 
        10'b0111111100: data <= 17'h1ff91; 
        10'b0111111101: data <= 17'h1fef7; 
        10'b0111111110: data <= 17'h1fe4b; 
        10'b0111111111: data <= 17'h1fde0; 
        10'b1000000000: data <= 17'h1fe07; 
        10'b1000000001: data <= 17'h1fe27; 
        10'b1000000010: data <= 17'h1fda0; 
        10'b1000000011: data <= 17'h1ff2f; 
        10'b1000000100: data <= 17'h1ffc1; 
        10'b1000000101: data <= 17'h00007; 
        10'b1000000110: data <= 17'h000ab; 
        10'b1000000111: data <= 17'h1ff4c; 
        10'b1000001000: data <= 17'h1ff22; 
        10'b1000001001: data <= 17'h1ff86; 
        10'b1000001010: data <= 17'h1fee9; 
        10'b1000001011: data <= 17'h1ff55; 
        10'b1000001100: data <= 17'h1fee1; 
        10'b1000001101: data <= 17'h1fe46; 
        10'b1000001110: data <= 17'h1febd; 
        10'b1000001111: data <= 17'h1ff34; 
        10'b1000010000: data <= 17'h1ff60; 
        10'b1000010001: data <= 17'h00011; 
        10'b1000010010: data <= 17'h1ffee; 
        10'b1000010011: data <= 17'h00004; 
        10'b1000010100: data <= 17'h00057; 
        10'b1000010101: data <= 17'h0005d; 
        10'b1000010110: data <= 17'h00055; 
        10'b1000010111: data <= 17'h0002a; 
        10'b1000011000: data <= 17'h1ffb5; 
        10'b1000011001: data <= 17'h1fea8; 
        10'b1000011010: data <= 17'h1fdd9; 
        10'b1000011011: data <= 17'h1fdb1; 
        10'b1000011100: data <= 17'h1fda1; 
        10'b1000011101: data <= 17'h1fd9e; 
        10'b1000011110: data <= 17'h1fe63; 
        10'b1000011111: data <= 17'h1fed6; 
        10'b1000100000: data <= 17'h1ff4e; 
        10'b1000100001: data <= 17'h0004d; 
        10'b1000100010: data <= 17'h000f2; 
        10'b1000100011: data <= 17'h1ff04; 
        10'b1000100100: data <= 17'h1ff0a; 
        10'b1000100101: data <= 17'h1fec9; 
        10'b1000100110: data <= 17'h1fe12; 
        10'b1000100111: data <= 17'h1fe2c; 
        10'b1000101000: data <= 17'h1fdbf; 
        10'b1000101001: data <= 17'h1fdec; 
        10'b1000101010: data <= 17'h1fe6b; 
        10'b1000101011: data <= 17'h1fee9; 
        10'b1000101100: data <= 17'h1ff72; 
        10'b1000101101: data <= 17'h1ffcb; 
        10'b1000101110: data <= 17'h00059; 
        10'b1000101111: data <= 17'h1ffd8; 
        10'b1000110000: data <= 17'h1ffd2; 
        10'b1000110001: data <= 17'h1ffeb; 
        10'b1000110010: data <= 17'h00024; 
        10'b1000110011: data <= 17'h1fff1; 
        10'b1000110100: data <= 17'h1ffa9; 
        10'b1000110101: data <= 17'h1fef7; 
        10'b1000110110: data <= 17'h1fdd5; 
        10'b1000110111: data <= 17'h1fdbd; 
        10'b1000111000: data <= 17'h1fdde; 
        10'b1000111001: data <= 17'h1fdeb; 
        10'b1000111010: data <= 17'h1fe8c; 
        10'b1000111011: data <= 17'h1fe81; 
        10'b1000111100: data <= 17'h0001c; 
        10'b1000111101: data <= 17'h00026; 
        10'b1000111110: data <= 17'h00080; 
        10'b1000111111: data <= 17'h1feae; 
        10'b1001000000: data <= 17'h1fe59; 
        10'b1001000001: data <= 17'h1fdd8; 
        10'b1001000010: data <= 17'h1fd06; 
        10'b1001000011: data <= 17'h1fe1b; 
        10'b1001000100: data <= 17'h1fd64; 
        10'b1001000101: data <= 17'h1fe02; 
        10'b1001000110: data <= 17'h1fe8f; 
        10'b1001000111: data <= 17'h1ff63; 
        10'b1001001000: data <= 17'h1ff97; 
        10'b1001001001: data <= 17'h0004f; 
        10'b1001001010: data <= 17'h0004b; 
        10'b1001001011: data <= 17'h00033; 
        10'b1001001100: data <= 17'h00047; 
        10'b1001001101: data <= 17'h0004b; 
        10'b1001001110: data <= 17'h00011; 
        10'b1001001111: data <= 17'h1ff9e; 
        10'b1001010000: data <= 17'h1ffcf; 
        10'b1001010001: data <= 17'h1ff13; 
        10'b1001010010: data <= 17'h1feeb; 
        10'b1001010011: data <= 17'h1fe70; 
        10'b1001010100: data <= 17'h1fe98; 
        10'b1001010101: data <= 17'h1ff2a; 
        10'b1001010110: data <= 17'h1fecf; 
        10'b1001010111: data <= 17'h1ff08; 
        10'b1001011000: data <= 17'h1ff91; 
        10'b1001011001: data <= 17'h0000f; 
        10'b1001011010: data <= 17'h1ffbd; 
        10'b1001011011: data <= 17'h1ff1c; 
        10'b1001011100: data <= 17'h1fefa; 
        10'b1001011101: data <= 17'h1fddf; 
        10'b1001011110: data <= 17'h1fde1; 
        10'b1001011111: data <= 17'h1fde0; 
        10'b1001100000: data <= 17'h1fdc3; 
        10'b1001100001: data <= 17'h1fe1b; 
        10'b1001100010: data <= 17'h1fee3; 
        10'b1001100011: data <= 17'h1ff29; 
        10'b1001100100: data <= 17'h1fff7; 
        10'b1001100101: data <= 17'h00021; 
        10'b1001100110: data <= 17'h00048; 
        10'b1001100111: data <= 17'h1fff0; 
        10'b1001101000: data <= 17'h00018; 
        10'b1001101001: data <= 17'h00006; 
        10'b1001101010: data <= 17'h00013; 
        10'b1001101011: data <= 17'h1ffc4; 
        10'b1001101100: data <= 17'h1ffe5; 
        10'b1001101101: data <= 17'h00023; 
        10'b1001101110: data <= 17'h1ffa9; 
        10'b1001101111: data <= 17'h0002b; 
        10'b1001110000: data <= 17'h00045; 
        10'b1001110001: data <= 17'h1ff93; 
        10'b1001110010: data <= 17'h1ff30; 
        10'b1001110011: data <= 17'h1fe9c; 
        10'b1001110100: data <= 17'h1feb4; 
        10'b1001110101: data <= 17'h1ff7a; 
        10'b1001110110: data <= 17'h00028; 
        10'b1001110111: data <= 17'h00027; 
        10'b1001111000: data <= 17'h1ff31; 
        10'b1001111001: data <= 17'h1ff00; 
        10'b1001111010: data <= 17'h1fe4c; 
        10'b1001111011: data <= 17'h1fe4c; 
        10'b1001111100: data <= 17'h1fe15; 
        10'b1001111101: data <= 17'h1fe52; 
        10'b1001111110: data <= 17'h1ff26; 
        10'b1001111111: data <= 17'h1ffb6; 
        10'b1010000000: data <= 17'h00030; 
        10'b1010000001: data <= 17'h1ffd2; 
        10'b1010000010: data <= 17'h00017; 
        10'b1010000011: data <= 17'h00001; 
        10'b1010000100: data <= 17'h00022; 
        10'b1010000101: data <= 17'h00044; 
        10'b1010000110: data <= 17'h1ffcc; 
        10'b1010000111: data <= 17'h1ffd0; 
        10'b1010001000: data <= 17'h0005a; 
        10'b1010001001: data <= 17'h00079; 
        10'b1010001010: data <= 17'h00106; 
        10'b1010001011: data <= 17'h0015e; 
        10'b1010001100: data <= 17'h000a7; 
        10'b1010001101: data <= 17'h00021; 
        10'b1010001110: data <= 17'h1ff99; 
        10'b1010001111: data <= 17'h1ff12; 
        10'b1010010000: data <= 17'h1ff3e; 
        10'b1010010001: data <= 17'h0000d; 
        10'b1010010010: data <= 17'h00088; 
        10'b1010010011: data <= 17'h0007e; 
        10'b1010010100: data <= 17'h1ffcc; 
        10'b1010010101: data <= 17'h1ffb2; 
        10'b1010010110: data <= 17'h1fee9; 
        10'b1010010111: data <= 17'h1fe7b; 
        10'b1010011000: data <= 17'h1fe72; 
        10'b1010011001: data <= 17'h1fec9; 
        10'b1010011010: data <= 17'h1feff; 
        10'b1010011011: data <= 17'h1ff59; 
        10'b1010011100: data <= 17'h1ffb6; 
        10'b1010011101: data <= 17'h00006; 
        10'b1010011110: data <= 17'h00005; 
        10'b1010011111: data <= 17'h1ffe4; 
        10'b1010100000: data <= 17'h1ffff; 
        10'b1010100001: data <= 17'h1fff7; 
        10'b1010100010: data <= 17'h00019; 
        10'b1010100011: data <= 17'h0003a; 
        10'b1010100100: data <= 17'h0007d; 
        10'b1010100101: data <= 17'h00120; 
        10'b1010100110: data <= 17'h001b4; 
        10'b1010100111: data <= 17'h001eb; 
        10'b1010101000: data <= 17'h001a1; 
        10'b1010101001: data <= 17'h000d7; 
        10'b1010101010: data <= 17'h001cf; 
        10'b1010101011: data <= 17'h00112; 
        10'b1010101100: data <= 17'h000ed; 
        10'b1010101101: data <= 17'h0014e; 
        10'b1010101110: data <= 17'h000ce; 
        10'b1010101111: data <= 17'h00129; 
        10'b1010110000: data <= 17'h000b0; 
        10'b1010110001: data <= 17'h00089; 
        10'b1010110010: data <= 17'h1fff7; 
        10'b1010110011: data <= 17'h1ff80; 
        10'b1010110100: data <= 17'h1ff78; 
        10'b1010110101: data <= 17'h1ff5b; 
        10'b1010110110: data <= 17'h1ff46; 
        10'b1010110111: data <= 17'h1ff56; 
        10'b1010111000: data <= 17'h0001a; 
        10'b1010111001: data <= 17'h1fff3; 
        10'b1010111010: data <= 17'h1ffd4; 
        10'b1010111011: data <= 17'h00033; 
        10'b1010111100: data <= 17'h1ffd3; 
        10'b1010111101: data <= 17'h00029; 
        10'b1010111110: data <= 17'h0004b; 
        10'b1010111111: data <= 17'h00046; 
        10'b1011000000: data <= 17'h00029; 
        10'b1011000001: data <= 17'h00090; 
        10'b1011000010: data <= 17'h000d4; 
        10'b1011000011: data <= 17'h00148; 
        10'b1011000100: data <= 17'h001fc; 
        10'b1011000101: data <= 17'h001f0; 
        10'b1011000110: data <= 17'h0024b; 
        10'b1011000111: data <= 17'h00222; 
        10'b1011001000: data <= 17'h001e6; 
        10'b1011001001: data <= 17'h00181; 
        10'b1011001010: data <= 17'h0018a; 
        10'b1011001011: data <= 17'h001a1; 
        10'b1011001100: data <= 17'h0015e; 
        10'b1011001101: data <= 17'h00147; 
        10'b1011001110: data <= 17'h00107; 
        10'b1011001111: data <= 17'h0005a; 
        10'b1011010000: data <= 17'h1ff91; 
        10'b1011010001: data <= 17'h0000f; 
        10'b1011010010: data <= 17'h1ffc9; 
        10'b1011010011: data <= 17'h1ffd8; 
        10'b1011010100: data <= 17'h1fff3; 
        10'b1011010101: data <= 17'h00019; 
        10'b1011010110: data <= 17'h00063; 
        10'b1011010111: data <= 17'h00041; 
        10'b1011011000: data <= 17'h1ffdd; 
        10'b1011011001: data <= 17'h00013; 
        10'b1011011010: data <= 17'h0005e; 
        10'b1011011011: data <= 17'h1fff0; 
        10'b1011011100: data <= 17'h1ffe0; 
        10'b1011011101: data <= 17'h00058; 
        10'b1011011110: data <= 17'h00006; 
        10'b1011011111: data <= 17'h00050; 
        10'b1011100000: data <= 17'h0004d; 
        10'b1011100001: data <= 17'h0000b; 
        10'b1011100010: data <= 17'h0006e; 
        10'b1011100011: data <= 17'h000a3; 
        10'b1011100100: data <= 17'h0002f; 
        10'b1011100101: data <= 17'h0008c; 
        10'b1011100110: data <= 17'h0012b; 
        10'b1011100111: data <= 17'h00172; 
        10'b1011101000: data <= 17'h00124; 
        10'b1011101001: data <= 17'h00176; 
        10'b1011101010: data <= 17'h000d5; 
        10'b1011101011: data <= 17'h00065; 
        10'b1011101100: data <= 17'h00003; 
        10'b1011101101: data <= 17'h00027; 
        10'b1011101110: data <= 17'h1fff6; 
        10'b1011101111: data <= 17'h00016; 
        10'b1011110000: data <= 17'h00004; 
        10'b1011110001: data <= 17'h1ffe7; 
        10'b1011110010: data <= 17'h1fffa; 
        10'b1011110011: data <= 17'h1fff3; 
        10'b1011110100: data <= 17'h1ffd2; 
        10'b1011110101: data <= 17'h00026; 
        10'b1011110110: data <= 17'h0001a; 
        10'b1011110111: data <= 17'h0002f; 
        10'b1011111000: data <= 17'h00040; 
        10'b1011111001: data <= 17'h00026; 
        10'b1011111010: data <= 17'h00011; 
        10'b1011111011: data <= 17'h00007; 
        10'b1011111100: data <= 17'h00069; 
        10'b1011111101: data <= 17'h00040; 
        10'b1011111110: data <= 17'h00013; 
        10'b1011111111: data <= 17'h00041; 
        10'b1100000000: data <= 17'h00020; 
        10'b1100000001: data <= 17'h0007a; 
        10'b1100000010: data <= 17'h00048; 
        10'b1100000011: data <= 17'h00037; 
        10'b1100000100: data <= 17'h000a9; 
        10'b1100000101: data <= 17'h00039; 
        10'b1100000110: data <= 17'h00033; 
        10'b1100000111: data <= 17'h00075; 
        10'b1100001000: data <= 17'h0000e; 
        10'b1100001001: data <= 17'h1ffec; 
        10'b1100001010: data <= 17'h00060; 
        10'b1100001011: data <= 17'h00034; 
        10'b1100001100: data <= 17'h00018; 
        10'b1100001101: data <= 17'h1ffef; 
        10'b1100001110: data <= 17'h1ffd9; 
        10'b1100001111: data <= 17'h00040; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 12) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 18'h0000c; 
        10'b0000000001: data <= 18'h00010; 
        10'b0000000010: data <= 18'h00079; 
        10'b0000000011: data <= 18'h0002f; 
        10'b0000000100: data <= 18'h000c6; 
        10'b0000000101: data <= 18'h3ffa8; 
        10'b0000000110: data <= 18'h3ffc5; 
        10'b0000000111: data <= 18'h00040; 
        10'b0000001000: data <= 18'h00098; 
        10'b0000001001: data <= 18'h00095; 
        10'b0000001010: data <= 18'h3ffac; 
        10'b0000001011: data <= 18'h00028; 
        10'b0000001100: data <= 18'h0002b; 
        10'b0000001101: data <= 18'h3ffea; 
        10'b0000001110: data <= 18'h0009f; 
        10'b0000001111: data <= 18'h0002b; 
        10'b0000010000: data <= 18'h00003; 
        10'b0000010001: data <= 18'h3fffa; 
        10'b0000010010: data <= 18'h00011; 
        10'b0000010011: data <= 18'h00037; 
        10'b0000010100: data <= 18'h00066; 
        10'b0000010101: data <= 18'h000c2; 
        10'b0000010110: data <= 18'h3ffcc; 
        10'b0000010111: data <= 18'h0008f; 
        10'b0000011000: data <= 18'h3ffec; 
        10'b0000011001: data <= 18'h00066; 
        10'b0000011010: data <= 18'h3fff8; 
        10'b0000011011: data <= 18'h3ffff; 
        10'b0000011100: data <= 18'h000b7; 
        10'b0000011101: data <= 18'h3ffd9; 
        10'b0000011110: data <= 18'h00029; 
        10'b0000011111: data <= 18'h000b4; 
        10'b0000100000: data <= 18'h00045; 
        10'b0000100001: data <= 18'h00007; 
        10'b0000100010: data <= 18'h000b3; 
        10'b0000100011: data <= 18'h00038; 
        10'b0000100100: data <= 18'h00011; 
        10'b0000100101: data <= 18'h3ffe2; 
        10'b0000100110: data <= 18'h3ffe8; 
        10'b0000100111: data <= 18'h3ffa2; 
        10'b0000101000: data <= 18'h0009a; 
        10'b0000101001: data <= 18'h3fff5; 
        10'b0000101010: data <= 18'h000b8; 
        10'b0000101011: data <= 18'h3ffd0; 
        10'b0000101100: data <= 18'h00050; 
        10'b0000101101: data <= 18'h0008b; 
        10'b0000101110: data <= 18'h0009c; 
        10'b0000101111: data <= 18'h0007c; 
        10'b0000110000: data <= 18'h00004; 
        10'b0000110001: data <= 18'h0007b; 
        10'b0000110010: data <= 18'h3fffc; 
        10'b0000110011: data <= 18'h000c2; 
        10'b0000110100: data <= 18'h00096; 
        10'b0000110101: data <= 18'h3ffca; 
        10'b0000110110: data <= 18'h3ffcb; 
        10'b0000110111: data <= 18'h0004f; 
        10'b0000111000: data <= 18'h000ad; 
        10'b0000111001: data <= 18'h000aa; 
        10'b0000111010: data <= 18'h00086; 
        10'b0000111011: data <= 18'h3ffe7; 
        10'b0000111100: data <= 18'h0009b; 
        10'b0000111101: data <= 18'h3ffb6; 
        10'b0000111110: data <= 18'h3ffc3; 
        10'b0000111111: data <= 18'h0007a; 
        10'b0001000000: data <= 18'h00067; 
        10'b0001000001: data <= 18'h3ffc4; 
        10'b0001000010: data <= 18'h3fff3; 
        10'b0001000011: data <= 18'h0004c; 
        10'b0001000100: data <= 18'h3ffeb; 
        10'b0001000101: data <= 18'h3ffd8; 
        10'b0001000110: data <= 18'h00030; 
        10'b0001000111: data <= 18'h0009c; 
        10'b0001001000: data <= 18'h0007e; 
        10'b0001001001: data <= 18'h00017; 
        10'b0001001010: data <= 18'h0003e; 
        10'b0001001011: data <= 18'h000b1; 
        10'b0001001100: data <= 18'h00096; 
        10'b0001001101: data <= 18'h000ae; 
        10'b0001001110: data <= 18'h3ffa9; 
        10'b0001001111: data <= 18'h00087; 
        10'b0001010000: data <= 18'h00033; 
        10'b0001010001: data <= 18'h00078; 
        10'b0001010010: data <= 18'h00067; 
        10'b0001010011: data <= 18'h00098; 
        10'b0001010100: data <= 18'h3fff2; 
        10'b0001010101: data <= 18'h0000a; 
        10'b0001010110: data <= 18'h0009e; 
        10'b0001010111: data <= 18'h3ffe8; 
        10'b0001011000: data <= 18'h00012; 
        10'b0001011001: data <= 18'h3fff5; 
        10'b0001011010: data <= 18'h3ffc6; 
        10'b0001011011: data <= 18'h00067; 
        10'b0001011100: data <= 18'h00001; 
        10'b0001011101: data <= 18'h00067; 
        10'b0001011110: data <= 18'h3ffab; 
        10'b0001011111: data <= 18'h00015; 
        10'b0001100000: data <= 18'h00053; 
        10'b0001100001: data <= 18'h3ff8e; 
        10'b0001100010: data <= 18'h0005e; 
        10'b0001100011: data <= 18'h3ffb3; 
        10'b0001100100: data <= 18'h3ff58; 
        10'b0001100101: data <= 18'h3ff77; 
        10'b0001100110: data <= 18'h3ff8a; 
        10'b0001100111: data <= 18'h3ffb1; 
        10'b0001101000: data <= 18'h3ffec; 
        10'b0001101001: data <= 18'h3ffb7; 
        10'b0001101010: data <= 18'h00040; 
        10'b0001101011: data <= 18'h3fff8; 
        10'b0001101100: data <= 18'h0004d; 
        10'b0001101101: data <= 18'h000c3; 
        10'b0001101110: data <= 18'h3ffc0; 
        10'b0001101111: data <= 18'h00051; 
        10'b0001110000: data <= 18'h000bd; 
        10'b0001110001: data <= 18'h3ffbb; 
        10'b0001110010: data <= 18'h00069; 
        10'b0001110011: data <= 18'h3ffb0; 
        10'b0001110100: data <= 18'h0002c; 
        10'b0001110101: data <= 18'h3ffdc; 
        10'b0001110110: data <= 18'h00008; 
        10'b0001110111: data <= 18'h3ffb2; 
        10'b0001111000: data <= 18'h0003b; 
        10'b0001111001: data <= 18'h3ffe4; 
        10'b0001111010: data <= 18'h3ff47; 
        10'b0001111011: data <= 18'h3fe9b; 
        10'b0001111100: data <= 18'h3fe89; 
        10'b0001111101: data <= 18'h3fe9a; 
        10'b0001111110: data <= 18'h3fe55; 
        10'b0001111111: data <= 18'h3fd41; 
        10'b0010000000: data <= 18'h3fe61; 
        10'b0010000001: data <= 18'h3fec8; 
        10'b0010000010: data <= 18'h3fef1; 
        10'b0010000011: data <= 18'h3ffb7; 
        10'b0010000100: data <= 18'h3ff35; 
        10'b0010000101: data <= 18'h0005e; 
        10'b0010000110: data <= 18'h0000e; 
        10'b0010000111: data <= 18'h3ff9e; 
        10'b0010001000: data <= 18'h000b3; 
        10'b0010001001: data <= 18'h3fffa; 
        10'b0010001010: data <= 18'h000b0; 
        10'b0010001011: data <= 18'h000aa; 
        10'b0010001100: data <= 18'h000a1; 
        10'b0010001101: data <= 18'h00006; 
        10'b0010001110: data <= 18'h0009b; 
        10'b0010001111: data <= 18'h3ffd6; 
        10'b0010010000: data <= 18'h3ff86; 
        10'b0010010001: data <= 18'h3ffeb; 
        10'b0010010010: data <= 18'h3ffa3; 
        10'b0010010011: data <= 18'h3ffde; 
        10'b0010010100: data <= 18'h3ff92; 
        10'b0010010101: data <= 18'h3ff00; 
        10'b0010010110: data <= 18'h3fd8a; 
        10'b0010010111: data <= 18'h3fcfb; 
        10'b0010011000: data <= 18'h3fc33; 
        10'b0010011001: data <= 18'h3fb8d; 
        10'b0010011010: data <= 18'h3fa72; 
        10'b0010011011: data <= 18'h3fa7d; 
        10'b0010011100: data <= 18'h3fa38; 
        10'b0010011101: data <= 18'h3fae6; 
        10'b0010011110: data <= 18'h3fbae; 
        10'b0010011111: data <= 18'h3fcb6; 
        10'b0010100000: data <= 18'h3fdaa; 
        10'b0010100001: data <= 18'h3ff2b; 
        10'b0010100010: data <= 18'h3feb6; 
        10'b0010100011: data <= 18'h3ffd7; 
        10'b0010100100: data <= 18'h00090; 
        10'b0010100101: data <= 18'h00073; 
        10'b0010100110: data <= 18'h3ffe2; 
        10'b0010100111: data <= 18'h00006; 
        10'b0010101000: data <= 18'h00086; 
        10'b0010101001: data <= 18'h000b8; 
        10'b0010101010: data <= 18'h0000d; 
        10'b0010101011: data <= 18'h0001e; 
        10'b0010101100: data <= 18'h000c7; 
        10'b0010101101: data <= 18'h000ec; 
        10'b0010101110: data <= 18'h00115; 
        10'b0010101111: data <= 18'h001a1; 
        10'b0010110000: data <= 18'h0026a; 
        10'b0010110001: data <= 18'h001ef; 
        10'b0010110010: data <= 18'h0020f; 
        10'b0010110011: data <= 18'h0005f; 
        10'b0010110100: data <= 18'h3fe59; 
        10'b0010110101: data <= 18'h3fc89; 
        10'b0010110110: data <= 18'h3fc62; 
        10'b0010110111: data <= 18'h3fe1f; 
        10'b0010111000: data <= 18'h3fedc; 
        10'b0010111001: data <= 18'h3fea6; 
        10'b0010111010: data <= 18'h3fe5c; 
        10'b0010111011: data <= 18'h3fe1a; 
        10'b0010111100: data <= 18'h3fd20; 
        10'b0010111101: data <= 18'h3feec; 
        10'b0010111110: data <= 18'h3fdfc; 
        10'b0010111111: data <= 18'h3fe89; 
        10'b0011000000: data <= 18'h3ff05; 
        10'b0011000001: data <= 18'h3ffac; 
        10'b0011000010: data <= 18'h3ffa9; 
        10'b0011000011: data <= 18'h00014; 
        10'b0011000100: data <= 18'h0007a; 
        10'b0011000101: data <= 18'h000b9; 
        10'b0011000110: data <= 18'h00098; 
        10'b0011000111: data <= 18'h00168; 
        10'b0011001000: data <= 18'h001b5; 
        10'b0011001001: data <= 18'h00189; 
        10'b0011001010: data <= 18'h00239; 
        10'b0011001011: data <= 18'h00365; 
        10'b0011001100: data <= 18'h004a7; 
        10'b0011001101: data <= 18'h003af; 
        10'b0011001110: data <= 18'h0028b; 
        10'b0011001111: data <= 18'h002cd; 
        10'b0011010000: data <= 18'h002fc; 
        10'b0011010001: data <= 18'h00093; 
        10'b0011010010: data <= 18'h0006c; 
        10'b0011010011: data <= 18'h00111; 
        10'b0011010100: data <= 18'h00326; 
        10'b0011010101: data <= 18'h00380; 
        10'b0011010110: data <= 18'h0025f; 
        10'b0011010111: data <= 18'h001e7; 
        10'b0011011000: data <= 18'h00077; 
        10'b0011011001: data <= 18'h3ff79; 
        10'b0011011010: data <= 18'h0003f; 
        10'b0011011011: data <= 18'h3ff6f; 
        10'b0011011100: data <= 18'h3ff78; 
        10'b0011011101: data <= 18'h3fff9; 
        10'b0011011110: data <= 18'h00060; 
        10'b0011011111: data <= 18'h3ffdc; 
        10'b0011100000: data <= 18'h3ffa3; 
        10'b0011100001: data <= 18'h000c2; 
        10'b0011100010: data <= 18'h0004b; 
        10'b0011100011: data <= 18'h00130; 
        10'b0011100100: data <= 18'h00268; 
        10'b0011100101: data <= 18'h0022b; 
        10'b0011100110: data <= 18'h002e8; 
        10'b0011100111: data <= 18'h00537; 
        10'b0011101000: data <= 18'h00383; 
        10'b0011101001: data <= 18'h0026b; 
        10'b0011101010: data <= 18'h00313; 
        10'b0011101011: data <= 18'h0041f; 
        10'b0011101100: data <= 18'h003eb; 
        10'b0011101101: data <= 18'h001f8; 
        10'b0011101110: data <= 18'h00127; 
        10'b0011101111: data <= 18'h00199; 
        10'b0011110000: data <= 18'h002c7; 
        10'b0011110001: data <= 18'h00445; 
        10'b0011110010: data <= 18'h002ed; 
        10'b0011110011: data <= 18'h00281; 
        10'b0011110100: data <= 18'h00200; 
        10'b0011110101: data <= 18'h0000c; 
        10'b0011110110: data <= 18'h00136; 
        10'b0011110111: data <= 18'h00107; 
        10'b0011111000: data <= 18'h3ff44; 
        10'b0011111001: data <= 18'h3ffa6; 
        10'b0011111010: data <= 18'h00068; 
        10'b0011111011: data <= 18'h000a0; 
        10'b0011111100: data <= 18'h00052; 
        10'b0011111101: data <= 18'h0009a; 
        10'b0011111110: data <= 18'h000cf; 
        10'b0011111111: data <= 18'h001b7; 
        10'b0100000000: data <= 18'h0025b; 
        10'b0100000001: data <= 18'h002ad; 
        10'b0100000010: data <= 18'h000fb; 
        10'b0100000011: data <= 18'h0014e; 
        10'b0100000100: data <= 18'h0017b; 
        10'b0100000101: data <= 18'h000fb; 
        10'b0100000110: data <= 18'h00266; 
        10'b0100000111: data <= 18'h002f1; 
        10'b0100001000: data <= 18'h003c0; 
        10'b0100001001: data <= 18'h0030d; 
        10'b0100001010: data <= 18'h0045f; 
        10'b0100001011: data <= 18'h00561; 
        10'b0100001100: data <= 18'h004f4; 
        10'b0100001101: data <= 18'h00587; 
        10'b0100001110: data <= 18'h0039c; 
        10'b0100001111: data <= 18'h003ad; 
        10'b0100010000: data <= 18'h00317; 
        10'b0100010001: data <= 18'h00294; 
        10'b0100010010: data <= 18'h00138; 
        10'b0100010011: data <= 18'h3ff8e; 
        10'b0100010100: data <= 18'h3ff40; 
        10'b0100010101: data <= 18'h3ffa2; 
        10'b0100010110: data <= 18'h00054; 
        10'b0100010111: data <= 18'h3ffd5; 
        10'b0100011000: data <= 18'h00020; 
        10'b0100011001: data <= 18'h000a8; 
        10'b0100011010: data <= 18'h000bb; 
        10'b0100011011: data <= 18'h00221; 
        10'b0100011100: data <= 18'h00271; 
        10'b0100011101: data <= 18'h00207; 
        10'b0100011110: data <= 18'h00060; 
        10'b0100011111: data <= 18'h0009c; 
        10'b0100100000: data <= 18'h3ff2e; 
        10'b0100100001: data <= 18'h3fff8; 
        10'b0100100010: data <= 18'h0017d; 
        10'b0100100011: data <= 18'h0029f; 
        10'b0100100100: data <= 18'h001d3; 
        10'b0100100101: data <= 18'h0043e; 
        10'b0100100110: data <= 18'h00576; 
        10'b0100100111: data <= 18'h006b5; 
        10'b0100101000: data <= 18'h007a2; 
        10'b0100101001: data <= 18'h005a9; 
        10'b0100101010: data <= 18'h00475; 
        10'b0100101011: data <= 18'h004a3; 
        10'b0100101100: data <= 18'h00412; 
        10'b0100101101: data <= 18'h00376; 
        10'b0100101110: data <= 18'h00188; 
        10'b0100101111: data <= 18'h3ff60; 
        10'b0100110000: data <= 18'h3fef8; 
        10'b0100110001: data <= 18'h3ff95; 
        10'b0100110010: data <= 18'h00014; 
        10'b0100110011: data <= 18'h3ffd8; 
        10'b0100110100: data <= 18'h00094; 
        10'b0100110101: data <= 18'h00068; 
        10'b0100110110: data <= 18'h000bd; 
        10'b0100110111: data <= 18'h0022e; 
        10'b0100111000: data <= 18'h002a1; 
        10'b0100111001: data <= 18'h0014e; 
        10'b0100111010: data <= 18'h00079; 
        10'b0100111011: data <= 18'h0006d; 
        10'b0100111100: data <= 18'h0001f; 
        10'b0100111101: data <= 18'h00194; 
        10'b0100111110: data <= 18'h000d0; 
        10'b0100111111: data <= 18'h00107; 
        10'b0101000000: data <= 18'h001b2; 
        10'b0101000001: data <= 18'h001ae; 
        10'b0101000010: data <= 18'h001c0; 
        10'b0101000011: data <= 18'h00522; 
        10'b0101000100: data <= 18'h006aa; 
        10'b0101000101: data <= 18'h00471; 
        10'b0101000110: data <= 18'h0047c; 
        10'b0101000111: data <= 18'h00373; 
        10'b0101001000: data <= 18'h0035a; 
        10'b0101001001: data <= 18'h0021b; 
        10'b0101001010: data <= 18'h00186; 
        10'b0101001011: data <= 18'h3ff79; 
        10'b0101001100: data <= 18'h3fe76; 
        10'b0101001101: data <= 18'h3fff5; 
        10'b0101001110: data <= 18'h00026; 
        10'b0101001111: data <= 18'h000ad; 
        10'b0101010000: data <= 18'h00084; 
        10'b0101010001: data <= 18'h3fff6; 
        10'b0101010010: data <= 18'h0005e; 
        10'b0101010011: data <= 18'h00160; 
        10'b0101010100: data <= 18'h0018b; 
        10'b0101010101: data <= 18'h00041; 
        10'b0101010110: data <= 18'h00058; 
        10'b0101010111: data <= 18'h00178; 
        10'b0101011000: data <= 18'h00102; 
        10'b0101011001: data <= 18'h3fff1; 
        10'b0101011010: data <= 18'h3fecd; 
        10'b0101011011: data <= 18'h3fcce; 
        10'b0101011100: data <= 18'h3f93f; 
        10'b0101011101: data <= 18'h3f58c; 
        10'b0101011110: data <= 18'h3f82d; 
        10'b0101011111: data <= 18'h0002c; 
        10'b0101100000: data <= 18'h0046b; 
        10'b0101100001: data <= 18'h00403; 
        10'b0101100010: data <= 18'h00194; 
        10'b0101100011: data <= 18'h00091; 
        10'b0101100100: data <= 18'h0001b; 
        10'b0101100101: data <= 18'h3ff6c; 
        10'b0101100110: data <= 18'h3ff7a; 
        10'b0101100111: data <= 18'h3ff0e; 
        10'b0101101000: data <= 18'h3ff52; 
        10'b0101101001: data <= 18'h000a3; 
        10'b0101101010: data <= 18'h00073; 
        10'b0101101011: data <= 18'h00001; 
        10'b0101101100: data <= 18'h0008f; 
        10'b0101101101: data <= 18'h00054; 
        10'b0101101110: data <= 18'h0009a; 
        10'b0101101111: data <= 18'h0013f; 
        10'b0101110000: data <= 18'h00077; 
        10'b0101110001: data <= 18'h00033; 
        10'b0101110010: data <= 18'h3ff97; 
        10'b0101110011: data <= 18'h00045; 
        10'b0101110100: data <= 18'h3ffd0; 
        10'b0101110101: data <= 18'h3fefa; 
        10'b0101110110: data <= 18'h3fca6; 
        10'b0101110111: data <= 18'h3f8ef; 
        10'b0101111000: data <= 18'h3f397; 
        10'b0101111001: data <= 18'h3f224; 
        10'b0101111010: data <= 18'h3f895; 
        10'b0101111011: data <= 18'h3ff07; 
        10'b0101111100: data <= 18'h00242; 
        10'b0101111101: data <= 18'h00174; 
        10'b0101111110: data <= 18'h00051; 
        10'b0101111111: data <= 18'h000a9; 
        10'b0110000000: data <= 18'h3fea4; 
        10'b0110000001: data <= 18'h3fe43; 
        10'b0110000010: data <= 18'h3ff98; 
        10'b0110000011: data <= 18'h00021; 
        10'b0110000100: data <= 18'h3ffab; 
        10'b0110000101: data <= 18'h3ffbc; 
        10'b0110000110: data <= 18'h0005a; 
        10'b0110000111: data <= 18'h3ffa8; 
        10'b0110001000: data <= 18'h3ffda; 
        10'b0110001001: data <= 18'h0004c; 
        10'b0110001010: data <= 18'h0011e; 
        10'b0110001011: data <= 18'h00164; 
        10'b0110001100: data <= 18'h000e2; 
        10'b0110001101: data <= 18'h00106; 
        10'b0110001110: data <= 18'h3ffa9; 
        10'b0110001111: data <= 18'h3ff49; 
        10'b0110010000: data <= 18'h3fe6d; 
        10'b0110010001: data <= 18'h3fc51; 
        10'b0110010010: data <= 18'h3fa95; 
        10'b0110010011: data <= 18'h3f79f; 
        10'b0110010100: data <= 18'h3f543; 
        10'b0110010101: data <= 18'h3f6f1; 
        10'b0110010110: data <= 18'h3fcae; 
        10'b0110010111: data <= 18'h00014; 
        10'b0110011000: data <= 18'h000b1; 
        10'b0110011001: data <= 18'h0016e; 
        10'b0110011010: data <= 18'h0041b; 
        10'b0110011011: data <= 18'h0046a; 
        10'b0110011100: data <= 18'h002a8; 
        10'b0110011101: data <= 18'h001b2; 
        10'b0110011110: data <= 18'h001b5; 
        10'b0110011111: data <= 18'h0017b; 
        10'b0110100000: data <= 18'h00080; 
        10'b0110100001: data <= 18'h00026; 
        10'b0110100010: data <= 18'h3ffc4; 
        10'b0110100011: data <= 18'h3ffc9; 
        10'b0110100100: data <= 18'h0005c; 
        10'b0110100101: data <= 18'h00088; 
        10'b0110100110: data <= 18'h00032; 
        10'b0110100111: data <= 18'h00087; 
        10'b0110101000: data <= 18'h00086; 
        10'b0110101001: data <= 18'h3fe83; 
        10'b0110101010: data <= 18'h3ff56; 
        10'b0110101011: data <= 18'h3ff14; 
        10'b0110101100: data <= 18'h3fc0c; 
        10'b0110101101: data <= 18'h3fb34; 
        10'b0110101110: data <= 18'h3f99f; 
        10'b0110101111: data <= 18'h3f8b1; 
        10'b0110110000: data <= 18'h3f80a; 
        10'b0110110001: data <= 18'h3fa22; 
        10'b0110110010: data <= 18'h3fc93; 
        10'b0110110011: data <= 18'h0001b; 
        10'b0110110100: data <= 18'h00060; 
        10'b0110110101: data <= 18'h00595; 
        10'b0110110110: data <= 18'h00689; 
        10'b0110110111: data <= 18'h00563; 
        10'b0110111000: data <= 18'h004c9; 
        10'b0110111001: data <= 18'h0041d; 
        10'b0110111010: data <= 18'h002a9; 
        10'b0110111011: data <= 18'h00134; 
        10'b0110111100: data <= 18'h3fff3; 
        10'b0110111101: data <= 18'h3ffab; 
        10'b0110111110: data <= 18'h00017; 
        10'b0110111111: data <= 18'h00093; 
        10'b0111000000: data <= 18'h0005b; 
        10'b0111000001: data <= 18'h000b5; 
        10'b0111000010: data <= 18'h3fff1; 
        10'b0111000011: data <= 18'h000be; 
        10'b0111000100: data <= 18'h00096; 
        10'b0111000101: data <= 18'h3ff56; 
        10'b0111000110: data <= 18'h3ff0f; 
        10'b0111000111: data <= 18'h3ffdd; 
        10'b0111001000: data <= 18'h3fcd1; 
        10'b0111001001: data <= 18'h3fc68; 
        10'b0111001010: data <= 18'h3fa37; 
        10'b0111001011: data <= 18'h3f91f; 
        10'b0111001100: data <= 18'h3fbb0; 
        10'b0111001101: data <= 18'h3fd97; 
        10'b0111001110: data <= 18'h3fc81; 
        10'b0111001111: data <= 18'h001cd; 
        10'b0111010000: data <= 18'h0022d; 
        10'b0111010001: data <= 18'h004b9; 
        10'b0111010010: data <= 18'h0040c; 
        10'b0111010011: data <= 18'h0043e; 
        10'b0111010100: data <= 18'h00360; 
        10'b0111010101: data <= 18'h00292; 
        10'b0111010110: data <= 18'h00082; 
        10'b0111010111: data <= 18'h3fef1; 
        10'b0111011000: data <= 18'h3ff58; 
        10'b0111011001: data <= 18'h3ffa0; 
        10'b0111011010: data <= 18'h00067; 
        10'b0111011011: data <= 18'h000b3; 
        10'b0111011100: data <= 18'h00006; 
        10'b0111011101: data <= 18'h00017; 
        10'b0111011110: data <= 18'h0006e; 
        10'b0111011111: data <= 18'h3fff8; 
        10'b0111100000: data <= 18'h00024; 
        10'b0111100001: data <= 18'h3ff93; 
        10'b0111100010: data <= 18'h3fddb; 
        10'b0111100011: data <= 18'h3fd2c; 
        10'b0111100100: data <= 18'h3fc74; 
        10'b0111100101: data <= 18'h3fd12; 
        10'b0111100110: data <= 18'h3fc1e; 
        10'b0111100111: data <= 18'h3fd1e; 
        10'b0111101000: data <= 18'h3ff14; 
        10'b0111101001: data <= 18'h000b8; 
        10'b0111101010: data <= 18'h00068; 
        10'b0111101011: data <= 18'h000b7; 
        10'b0111101100: data <= 18'h3ff93; 
        10'b0111101101: data <= 18'h00123; 
        10'b0111101110: data <= 18'h00103; 
        10'b0111101111: data <= 18'h000b8; 
        10'b0111110000: data <= 18'h00062; 
        10'b0111110001: data <= 18'h3ff69; 
        10'b0111110010: data <= 18'h3feb2; 
        10'b0111110011: data <= 18'h3ff6a; 
        10'b0111110100: data <= 18'h3ff7d; 
        10'b0111110101: data <= 18'h3ff99; 
        10'b0111110110: data <= 18'h3ffc9; 
        10'b0111110111: data <= 18'h3ffce; 
        10'b0111111000: data <= 18'h3ffce; 
        10'b0111111001: data <= 18'h3fff0; 
        10'b0111111010: data <= 18'h0007c; 
        10'b0111111011: data <= 18'h00026; 
        10'b0111111100: data <= 18'h3ff22; 
        10'b0111111101: data <= 18'h3fdef; 
        10'b0111111110: data <= 18'h3fc96; 
        10'b0111111111: data <= 18'h3fbc0; 
        10'b1000000000: data <= 18'h3fc0e; 
        10'b1000000001: data <= 18'h3fc4e; 
        10'b1000000010: data <= 18'h3fb41; 
        10'b1000000011: data <= 18'h3fe5e; 
        10'b1000000100: data <= 18'h3ff82; 
        10'b1000000101: data <= 18'h0000f; 
        10'b1000000110: data <= 18'h00156; 
        10'b1000000111: data <= 18'h3fe97; 
        10'b1000001000: data <= 18'h3fe45; 
        10'b1000001001: data <= 18'h3ff0b; 
        10'b1000001010: data <= 18'h3fdd2; 
        10'b1000001011: data <= 18'h3feaa; 
        10'b1000001100: data <= 18'h3fdc1; 
        10'b1000001101: data <= 18'h3fc8d; 
        10'b1000001110: data <= 18'h3fd7a; 
        10'b1000001111: data <= 18'h3fe68; 
        10'b1000010000: data <= 18'h3febf; 
        10'b1000010001: data <= 18'h00021; 
        10'b1000010010: data <= 18'h3ffdd; 
        10'b1000010011: data <= 18'h00008; 
        10'b1000010100: data <= 18'h000ad; 
        10'b1000010101: data <= 18'h000b9; 
        10'b1000010110: data <= 18'h000aa; 
        10'b1000010111: data <= 18'h00055; 
        10'b1000011000: data <= 18'h3ff6a; 
        10'b1000011001: data <= 18'h3fd50; 
        10'b1000011010: data <= 18'h3fbb3; 
        10'b1000011011: data <= 18'h3fb62; 
        10'b1000011100: data <= 18'h3fb43; 
        10'b1000011101: data <= 18'h3fb3b; 
        10'b1000011110: data <= 18'h3fcc5; 
        10'b1000011111: data <= 18'h3fdad; 
        10'b1000100000: data <= 18'h3fe9c; 
        10'b1000100001: data <= 18'h0009a; 
        10'b1000100010: data <= 18'h001e4; 
        10'b1000100011: data <= 18'h3fe07; 
        10'b1000100100: data <= 18'h3fe13; 
        10'b1000100101: data <= 18'h3fd92; 
        10'b1000100110: data <= 18'h3fc23; 
        10'b1000100111: data <= 18'h3fc57; 
        10'b1000101000: data <= 18'h3fb7f; 
        10'b1000101001: data <= 18'h3fbd7; 
        10'b1000101010: data <= 18'h3fcd5; 
        10'b1000101011: data <= 18'h3fdd2; 
        10'b1000101100: data <= 18'h3fee5; 
        10'b1000101101: data <= 18'h3ff97; 
        10'b1000101110: data <= 18'h000b2; 
        10'b1000101111: data <= 18'h3ffb0; 
        10'b1000110000: data <= 18'h3ffa4; 
        10'b1000110001: data <= 18'h3ffd6; 
        10'b1000110010: data <= 18'h00049; 
        10'b1000110011: data <= 18'h3ffe2; 
        10'b1000110100: data <= 18'h3ff52; 
        10'b1000110101: data <= 18'h3fded; 
        10'b1000110110: data <= 18'h3fbaa; 
        10'b1000110111: data <= 18'h3fb7b; 
        10'b1000111000: data <= 18'h3fbbc; 
        10'b1000111001: data <= 18'h3fbd6; 
        10'b1000111010: data <= 18'h3fd19; 
        10'b1000111011: data <= 18'h3fd01; 
        10'b1000111100: data <= 18'h00038; 
        10'b1000111101: data <= 18'h0004c; 
        10'b1000111110: data <= 18'h00101; 
        10'b1000111111: data <= 18'h3fd5b; 
        10'b1001000000: data <= 18'h3fcb2; 
        10'b1001000001: data <= 18'h3fbaf; 
        10'b1001000010: data <= 18'h3fa0b; 
        10'b1001000011: data <= 18'h3fc36; 
        10'b1001000100: data <= 18'h3fac7; 
        10'b1001000101: data <= 18'h3fc05; 
        10'b1001000110: data <= 18'h3fd1f; 
        10'b1001000111: data <= 18'h3fec6; 
        10'b1001001000: data <= 18'h3ff2f; 
        10'b1001001001: data <= 18'h0009e; 
        10'b1001001010: data <= 18'h00096; 
        10'b1001001011: data <= 18'h00066; 
        10'b1001001100: data <= 18'h0008e; 
        10'b1001001101: data <= 18'h00095; 
        10'b1001001110: data <= 18'h00021; 
        10'b1001001111: data <= 18'h3ff3d; 
        10'b1001010000: data <= 18'h3ff9d; 
        10'b1001010001: data <= 18'h3fe27; 
        10'b1001010010: data <= 18'h3fdd5; 
        10'b1001010011: data <= 18'h3fce1; 
        10'b1001010100: data <= 18'h3fd30; 
        10'b1001010101: data <= 18'h3fe54; 
        10'b1001010110: data <= 18'h3fd9f; 
        10'b1001010111: data <= 18'h3fe0f; 
        10'b1001011000: data <= 18'h3ff22; 
        10'b1001011001: data <= 18'h0001e; 
        10'b1001011010: data <= 18'h3ff7b; 
        10'b1001011011: data <= 18'h3fe38; 
        10'b1001011100: data <= 18'h3fdf3; 
        10'b1001011101: data <= 18'h3fbbe; 
        10'b1001011110: data <= 18'h3fbc3; 
        10'b1001011111: data <= 18'h3fbc0; 
        10'b1001100000: data <= 18'h3fb86; 
        10'b1001100001: data <= 18'h3fc36; 
        10'b1001100010: data <= 18'h3fdc6; 
        10'b1001100011: data <= 18'h3fe51; 
        10'b1001100100: data <= 18'h3ffed; 
        10'b1001100101: data <= 18'h00042; 
        10'b1001100110: data <= 18'h00090; 
        10'b1001100111: data <= 18'h3ffe1; 
        10'b1001101000: data <= 18'h00031; 
        10'b1001101001: data <= 18'h0000b; 
        10'b1001101010: data <= 18'h00026; 
        10'b1001101011: data <= 18'h3ff88; 
        10'b1001101100: data <= 18'h3ffc9; 
        10'b1001101101: data <= 18'h00046; 
        10'b1001101110: data <= 18'h3ff53; 
        10'b1001101111: data <= 18'h00056; 
        10'b1001110000: data <= 18'h00089; 
        10'b1001110001: data <= 18'h3ff25; 
        10'b1001110010: data <= 18'h3fe5f; 
        10'b1001110011: data <= 18'h3fd39; 
        10'b1001110100: data <= 18'h3fd67; 
        10'b1001110101: data <= 18'h3fef4; 
        10'b1001110110: data <= 18'h00050; 
        10'b1001110111: data <= 18'h0004e; 
        10'b1001111000: data <= 18'h3fe63; 
        10'b1001111001: data <= 18'h3fe00; 
        10'b1001111010: data <= 18'h3fc98; 
        10'b1001111011: data <= 18'h3fc98; 
        10'b1001111100: data <= 18'h3fc29; 
        10'b1001111101: data <= 18'h3fca4; 
        10'b1001111110: data <= 18'h3fe4b; 
        10'b1001111111: data <= 18'h3ff6c; 
        10'b1010000000: data <= 18'h0005f; 
        10'b1010000001: data <= 18'h3ffa3; 
        10'b1010000010: data <= 18'h0002d; 
        10'b1010000011: data <= 18'h00003; 
        10'b1010000100: data <= 18'h00043; 
        10'b1010000101: data <= 18'h00088; 
        10'b1010000110: data <= 18'h3ff97; 
        10'b1010000111: data <= 18'h3ffa1; 
        10'b1010001000: data <= 18'h000b4; 
        10'b1010001001: data <= 18'h000f1; 
        10'b1010001010: data <= 18'h0020d; 
        10'b1010001011: data <= 18'h002bc; 
        10'b1010001100: data <= 18'h0014e; 
        10'b1010001101: data <= 18'h00043; 
        10'b1010001110: data <= 18'h3ff32; 
        10'b1010001111: data <= 18'h3fe24; 
        10'b1010010000: data <= 18'h3fe7b; 
        10'b1010010001: data <= 18'h0001b; 
        10'b1010010010: data <= 18'h00111; 
        10'b1010010011: data <= 18'h000fb; 
        10'b1010010100: data <= 18'h3ff97; 
        10'b1010010101: data <= 18'h3ff65; 
        10'b1010010110: data <= 18'h3fdd2; 
        10'b1010010111: data <= 18'h3fcf5; 
        10'b1010011000: data <= 18'h3fce3; 
        10'b1010011001: data <= 18'h3fd92; 
        10'b1010011010: data <= 18'h3fdff; 
        10'b1010011011: data <= 18'h3feb1; 
        10'b1010011100: data <= 18'h3ff6c; 
        10'b1010011101: data <= 18'h0000b; 
        10'b1010011110: data <= 18'h0000a; 
        10'b1010011111: data <= 18'h3ffc9; 
        10'b1010100000: data <= 18'h3ffff; 
        10'b1010100001: data <= 18'h3ffee; 
        10'b1010100010: data <= 18'h00032; 
        10'b1010100011: data <= 18'h00075; 
        10'b1010100100: data <= 18'h000fa; 
        10'b1010100101: data <= 18'h00240; 
        10'b1010100110: data <= 18'h00367; 
        10'b1010100111: data <= 18'h003d6; 
        10'b1010101000: data <= 18'h00342; 
        10'b1010101001: data <= 18'h001ae; 
        10'b1010101010: data <= 18'h0039f; 
        10'b1010101011: data <= 18'h00223; 
        10'b1010101100: data <= 18'h001db; 
        10'b1010101101: data <= 18'h0029d; 
        10'b1010101110: data <= 18'h0019c; 
        10'b1010101111: data <= 18'h00252; 
        10'b1010110000: data <= 18'h00160; 
        10'b1010110001: data <= 18'h00112; 
        10'b1010110010: data <= 18'h3ffee; 
        10'b1010110011: data <= 18'h3ff00; 
        10'b1010110100: data <= 18'h3fef0; 
        10'b1010110101: data <= 18'h3feb6; 
        10'b1010110110: data <= 18'h3fe8b; 
        10'b1010110111: data <= 18'h3fead; 
        10'b1010111000: data <= 18'h00034; 
        10'b1010111001: data <= 18'h3ffe5; 
        10'b1010111010: data <= 18'h3ffa7; 
        10'b1010111011: data <= 18'h00066; 
        10'b1010111100: data <= 18'h3ffa5; 
        10'b1010111101: data <= 18'h00053; 
        10'b1010111110: data <= 18'h00096; 
        10'b1010111111: data <= 18'h0008d; 
        10'b1011000000: data <= 18'h00052; 
        10'b1011000001: data <= 18'h0011f; 
        10'b1011000010: data <= 18'h001a9; 
        10'b1011000011: data <= 18'h00291; 
        10'b1011000100: data <= 18'h003f7; 
        10'b1011000101: data <= 18'h003df; 
        10'b1011000110: data <= 18'h00495; 
        10'b1011000111: data <= 18'h00444; 
        10'b1011001000: data <= 18'h003cd; 
        10'b1011001001: data <= 18'h00303; 
        10'b1011001010: data <= 18'h00313; 
        10'b1011001011: data <= 18'h00342; 
        10'b1011001100: data <= 18'h002bb; 
        10'b1011001101: data <= 18'h0028d; 
        10'b1011001110: data <= 18'h0020f; 
        10'b1011001111: data <= 18'h000b5; 
        10'b1011010000: data <= 18'h3ff22; 
        10'b1011010001: data <= 18'h0001e; 
        10'b1011010010: data <= 18'h3ff92; 
        10'b1011010011: data <= 18'h3ffaf; 
        10'b1011010100: data <= 18'h3ffe6; 
        10'b1011010101: data <= 18'h00032; 
        10'b1011010110: data <= 18'h000c7; 
        10'b1011010111: data <= 18'h00081; 
        10'b1011011000: data <= 18'h3ffb9; 
        10'b1011011001: data <= 18'h00026; 
        10'b1011011010: data <= 18'h000bc; 
        10'b1011011011: data <= 18'h3ffe0; 
        10'b1011011100: data <= 18'h3ffc0; 
        10'b1011011101: data <= 18'h000b0; 
        10'b1011011110: data <= 18'h0000d; 
        10'b1011011111: data <= 18'h000a1; 
        10'b1011100000: data <= 18'h00099; 
        10'b1011100001: data <= 18'h00015; 
        10'b1011100010: data <= 18'h000dd; 
        10'b1011100011: data <= 18'h00145; 
        10'b1011100100: data <= 18'h0005e; 
        10'b1011100101: data <= 18'h00117; 
        10'b1011100110: data <= 18'h00257; 
        10'b1011100111: data <= 18'h002e4; 
        10'b1011101000: data <= 18'h00247; 
        10'b1011101001: data <= 18'h002ec; 
        10'b1011101010: data <= 18'h001aa; 
        10'b1011101011: data <= 18'h000c9; 
        10'b1011101100: data <= 18'h00007; 
        10'b1011101101: data <= 18'h0004d; 
        10'b1011101110: data <= 18'h3ffeb; 
        10'b1011101111: data <= 18'h0002b; 
        10'b1011110000: data <= 18'h00009; 
        10'b1011110001: data <= 18'h3ffce; 
        10'b1011110010: data <= 18'h3fff4; 
        10'b1011110011: data <= 18'h3ffe7; 
        10'b1011110100: data <= 18'h3ffa3; 
        10'b1011110101: data <= 18'h0004c; 
        10'b1011110110: data <= 18'h00033; 
        10'b1011110111: data <= 18'h0005e; 
        10'b1011111000: data <= 18'h00080; 
        10'b1011111001: data <= 18'h0004d; 
        10'b1011111010: data <= 18'h00021; 
        10'b1011111011: data <= 18'h0000e; 
        10'b1011111100: data <= 18'h000d2; 
        10'b1011111101: data <= 18'h00081; 
        10'b1011111110: data <= 18'h00026; 
        10'b1011111111: data <= 18'h00082; 
        10'b1100000000: data <= 18'h0003f; 
        10'b1100000001: data <= 18'h000f3; 
        10'b1100000010: data <= 18'h00091; 
        10'b1100000011: data <= 18'h0006f; 
        10'b1100000100: data <= 18'h00152; 
        10'b1100000101: data <= 18'h00072; 
        10'b1100000110: data <= 18'h00065; 
        10'b1100000111: data <= 18'h000eb; 
        10'b1100001000: data <= 18'h0001c; 
        10'b1100001001: data <= 18'h3ffd8; 
        10'b1100001010: data <= 18'h000bf; 
        10'b1100001011: data <= 18'h00069; 
        10'b1100001100: data <= 18'h00031; 
        10'b1100001101: data <= 18'h3ffdd; 
        10'b1100001110: data <= 18'h3ffb2; 
        10'b1100001111: data <= 18'h0007f; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 13) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 19'h00018; 
        10'b0000000001: data <= 19'h00020; 
        10'b0000000010: data <= 19'h000f3; 
        10'b0000000011: data <= 19'h0005e; 
        10'b0000000100: data <= 19'h0018c; 
        10'b0000000101: data <= 19'h7ff50; 
        10'b0000000110: data <= 19'h7ff8a; 
        10'b0000000111: data <= 19'h00081; 
        10'b0000001000: data <= 19'h00131; 
        10'b0000001001: data <= 19'h0012a; 
        10'b0000001010: data <= 19'h7ff57; 
        10'b0000001011: data <= 19'h00050; 
        10'b0000001100: data <= 19'h00056; 
        10'b0000001101: data <= 19'h7ffd3; 
        10'b0000001110: data <= 19'h0013f; 
        10'b0000001111: data <= 19'h00055; 
        10'b0000010000: data <= 19'h00006; 
        10'b0000010001: data <= 19'h7fff5; 
        10'b0000010010: data <= 19'h00022; 
        10'b0000010011: data <= 19'h0006e; 
        10'b0000010100: data <= 19'h000cd; 
        10'b0000010101: data <= 19'h00184; 
        10'b0000010110: data <= 19'h7ff98; 
        10'b0000010111: data <= 19'h0011d; 
        10'b0000011000: data <= 19'h7ffd8; 
        10'b0000011001: data <= 19'h000cd; 
        10'b0000011010: data <= 19'h7ffef; 
        10'b0000011011: data <= 19'h7ffff; 
        10'b0000011100: data <= 19'h0016d; 
        10'b0000011101: data <= 19'h7ffb2; 
        10'b0000011110: data <= 19'h00052; 
        10'b0000011111: data <= 19'h00168; 
        10'b0000100000: data <= 19'h0008a; 
        10'b0000100001: data <= 19'h0000d; 
        10'b0000100010: data <= 19'h00165; 
        10'b0000100011: data <= 19'h00071; 
        10'b0000100100: data <= 19'h00022; 
        10'b0000100101: data <= 19'h7ffc3; 
        10'b0000100110: data <= 19'h7ffd0; 
        10'b0000100111: data <= 19'h7ff44; 
        10'b0000101000: data <= 19'h00133; 
        10'b0000101001: data <= 19'h7ffea; 
        10'b0000101010: data <= 19'h00171; 
        10'b0000101011: data <= 19'h7ffa0; 
        10'b0000101100: data <= 19'h000a0; 
        10'b0000101101: data <= 19'h00115; 
        10'b0000101110: data <= 19'h00138; 
        10'b0000101111: data <= 19'h000f9; 
        10'b0000110000: data <= 19'h00008; 
        10'b0000110001: data <= 19'h000f5; 
        10'b0000110010: data <= 19'h7fff9; 
        10'b0000110011: data <= 19'h00185; 
        10'b0000110100: data <= 19'h0012c; 
        10'b0000110101: data <= 19'h7ff94; 
        10'b0000110110: data <= 19'h7ff96; 
        10'b0000110111: data <= 19'h0009f; 
        10'b0000111000: data <= 19'h0015a; 
        10'b0000111001: data <= 19'h00155; 
        10'b0000111010: data <= 19'h0010c; 
        10'b0000111011: data <= 19'h7ffce; 
        10'b0000111100: data <= 19'h00137; 
        10'b0000111101: data <= 19'h7ff6c; 
        10'b0000111110: data <= 19'h7ff87; 
        10'b0000111111: data <= 19'h000f3; 
        10'b0001000000: data <= 19'h000cd; 
        10'b0001000001: data <= 19'h7ff88; 
        10'b0001000010: data <= 19'h7ffe5; 
        10'b0001000011: data <= 19'h00097; 
        10'b0001000100: data <= 19'h7ffd6; 
        10'b0001000101: data <= 19'h7ffb0; 
        10'b0001000110: data <= 19'h0005f; 
        10'b0001000111: data <= 19'h00139; 
        10'b0001001000: data <= 19'h000fd; 
        10'b0001001001: data <= 19'h0002f; 
        10'b0001001010: data <= 19'h0007c; 
        10'b0001001011: data <= 19'h00161; 
        10'b0001001100: data <= 19'h0012c; 
        10'b0001001101: data <= 19'h0015b; 
        10'b0001001110: data <= 19'h7ff51; 
        10'b0001001111: data <= 19'h0010f; 
        10'b0001010000: data <= 19'h00067; 
        10'b0001010001: data <= 19'h000ef; 
        10'b0001010010: data <= 19'h000ce; 
        10'b0001010011: data <= 19'h00131; 
        10'b0001010100: data <= 19'h7ffe4; 
        10'b0001010101: data <= 19'h00015; 
        10'b0001010110: data <= 19'h0013d; 
        10'b0001010111: data <= 19'h7ffd0; 
        10'b0001011000: data <= 19'h00024; 
        10'b0001011001: data <= 19'h7ffeb; 
        10'b0001011010: data <= 19'h7ff8b; 
        10'b0001011011: data <= 19'h000ce; 
        10'b0001011100: data <= 19'h00002; 
        10'b0001011101: data <= 19'h000ce; 
        10'b0001011110: data <= 19'h7ff57; 
        10'b0001011111: data <= 19'h0002a; 
        10'b0001100000: data <= 19'h000a6; 
        10'b0001100001: data <= 19'h7ff1c; 
        10'b0001100010: data <= 19'h000bc; 
        10'b0001100011: data <= 19'h7ff65; 
        10'b0001100100: data <= 19'h7feb0; 
        10'b0001100101: data <= 19'h7feed; 
        10'b0001100110: data <= 19'h7ff14; 
        10'b0001100111: data <= 19'h7ff61; 
        10'b0001101000: data <= 19'h7ffd8; 
        10'b0001101001: data <= 19'h7ff6e; 
        10'b0001101010: data <= 19'h0007f; 
        10'b0001101011: data <= 19'h7fff0; 
        10'b0001101100: data <= 19'h0009a; 
        10'b0001101101: data <= 19'h00186; 
        10'b0001101110: data <= 19'h7ff80; 
        10'b0001101111: data <= 19'h000a1; 
        10'b0001110000: data <= 19'h0017a; 
        10'b0001110001: data <= 19'h7ff76; 
        10'b0001110010: data <= 19'h000d3; 
        10'b0001110011: data <= 19'h7ff5f; 
        10'b0001110100: data <= 19'h00058; 
        10'b0001110101: data <= 19'h7ffb7; 
        10'b0001110110: data <= 19'h00011; 
        10'b0001110111: data <= 19'h7ff65; 
        10'b0001111000: data <= 19'h00076; 
        10'b0001111001: data <= 19'h7ffc9; 
        10'b0001111010: data <= 19'h7fe8e; 
        10'b0001111011: data <= 19'h7fd36; 
        10'b0001111100: data <= 19'h7fd12; 
        10'b0001111101: data <= 19'h7fd34; 
        10'b0001111110: data <= 19'h7fcaa; 
        10'b0001111111: data <= 19'h7fa82; 
        10'b0010000000: data <= 19'h7fcc3; 
        10'b0010000001: data <= 19'h7fd8f; 
        10'b0010000010: data <= 19'h7fde1; 
        10'b0010000011: data <= 19'h7ff6d; 
        10'b0010000100: data <= 19'h7fe6b; 
        10'b0010000101: data <= 19'h000bd; 
        10'b0010000110: data <= 19'h0001d; 
        10'b0010000111: data <= 19'h7ff3b; 
        10'b0010001000: data <= 19'h00166; 
        10'b0010001001: data <= 19'h7fff3; 
        10'b0010001010: data <= 19'h0015f; 
        10'b0010001011: data <= 19'h00154; 
        10'b0010001100: data <= 19'h00142; 
        10'b0010001101: data <= 19'h0000d; 
        10'b0010001110: data <= 19'h00137; 
        10'b0010001111: data <= 19'h7ffab; 
        10'b0010010000: data <= 19'h7ff0d; 
        10'b0010010001: data <= 19'h7ffd6; 
        10'b0010010010: data <= 19'h7ff46; 
        10'b0010010011: data <= 19'h7ffbc; 
        10'b0010010100: data <= 19'h7ff23; 
        10'b0010010101: data <= 19'h7fdff; 
        10'b0010010110: data <= 19'h7fb15; 
        10'b0010010111: data <= 19'h7f9f6; 
        10'b0010011000: data <= 19'h7f867; 
        10'b0010011001: data <= 19'h7f719; 
        10'b0010011010: data <= 19'h7f4e4; 
        10'b0010011011: data <= 19'h7f4fa; 
        10'b0010011100: data <= 19'h7f470; 
        10'b0010011101: data <= 19'h7f5cd; 
        10'b0010011110: data <= 19'h7f75b; 
        10'b0010011111: data <= 19'h7f96d; 
        10'b0010100000: data <= 19'h7fb54; 
        10'b0010100001: data <= 19'h7fe55; 
        10'b0010100010: data <= 19'h7fd6c; 
        10'b0010100011: data <= 19'h7ffad; 
        10'b0010100100: data <= 19'h00121; 
        10'b0010100101: data <= 19'h000e6; 
        10'b0010100110: data <= 19'h7ffc5; 
        10'b0010100111: data <= 19'h0000d; 
        10'b0010101000: data <= 19'h0010c; 
        10'b0010101001: data <= 19'h0016f; 
        10'b0010101010: data <= 19'h0001a; 
        10'b0010101011: data <= 19'h0003c; 
        10'b0010101100: data <= 19'h0018d; 
        10'b0010101101: data <= 19'h001d9; 
        10'b0010101110: data <= 19'h0022a; 
        10'b0010101111: data <= 19'h00341; 
        10'b0010110000: data <= 19'h004d4; 
        10'b0010110001: data <= 19'h003de; 
        10'b0010110010: data <= 19'h0041e; 
        10'b0010110011: data <= 19'h000bd; 
        10'b0010110100: data <= 19'h7fcb3; 
        10'b0010110101: data <= 19'h7f912; 
        10'b0010110110: data <= 19'h7f8c5; 
        10'b0010110111: data <= 19'h7fc3f; 
        10'b0010111000: data <= 19'h7fdb8; 
        10'b0010111001: data <= 19'h7fd4b; 
        10'b0010111010: data <= 19'h7fcb8; 
        10'b0010111011: data <= 19'h7fc34; 
        10'b0010111100: data <= 19'h7fa40; 
        10'b0010111101: data <= 19'h7fdd8; 
        10'b0010111110: data <= 19'h7fbf9; 
        10'b0010111111: data <= 19'h7fd11; 
        10'b0011000000: data <= 19'h7fe0a; 
        10'b0011000001: data <= 19'h7ff57; 
        10'b0011000010: data <= 19'h7ff52; 
        10'b0011000011: data <= 19'h00028; 
        10'b0011000100: data <= 19'h000f4; 
        10'b0011000101: data <= 19'h00172; 
        10'b0011000110: data <= 19'h00131; 
        10'b0011000111: data <= 19'h002d0; 
        10'b0011001000: data <= 19'h00369; 
        10'b0011001001: data <= 19'h00311; 
        10'b0011001010: data <= 19'h00471; 
        10'b0011001011: data <= 19'h006cb; 
        10'b0011001100: data <= 19'h0094d; 
        10'b0011001101: data <= 19'h0075f; 
        10'b0011001110: data <= 19'h00516; 
        10'b0011001111: data <= 19'h0059a; 
        10'b0011010000: data <= 19'h005f7; 
        10'b0011010001: data <= 19'h00126; 
        10'b0011010010: data <= 19'h000d9; 
        10'b0011010011: data <= 19'h00223; 
        10'b0011010100: data <= 19'h0064c; 
        10'b0011010101: data <= 19'h00700; 
        10'b0011010110: data <= 19'h004be; 
        10'b0011010111: data <= 19'h003ce; 
        10'b0011011000: data <= 19'h000ed; 
        10'b0011011001: data <= 19'h7fef3; 
        10'b0011011010: data <= 19'h0007e; 
        10'b0011011011: data <= 19'h7fede; 
        10'b0011011100: data <= 19'h7fef0; 
        10'b0011011101: data <= 19'h7fff2; 
        10'b0011011110: data <= 19'h000c0; 
        10'b0011011111: data <= 19'h7ffb8; 
        10'b0011100000: data <= 19'h7ff45; 
        10'b0011100001: data <= 19'h00184; 
        10'b0011100010: data <= 19'h00096; 
        10'b0011100011: data <= 19'h00260; 
        10'b0011100100: data <= 19'h004d0; 
        10'b0011100101: data <= 19'h00457; 
        10'b0011100110: data <= 19'h005cf; 
        10'b0011100111: data <= 19'h00a6e; 
        10'b0011101000: data <= 19'h00705; 
        10'b0011101001: data <= 19'h004d6; 
        10'b0011101010: data <= 19'h00627; 
        10'b0011101011: data <= 19'h0083d; 
        10'b0011101100: data <= 19'h007d5; 
        10'b0011101101: data <= 19'h003f1; 
        10'b0011101110: data <= 19'h0024e; 
        10'b0011101111: data <= 19'h00332; 
        10'b0011110000: data <= 19'h0058e; 
        10'b0011110001: data <= 19'h0088a; 
        10'b0011110010: data <= 19'h005da; 
        10'b0011110011: data <= 19'h00503; 
        10'b0011110100: data <= 19'h00400; 
        10'b0011110101: data <= 19'h00018; 
        10'b0011110110: data <= 19'h0026d; 
        10'b0011110111: data <= 19'h0020f; 
        10'b0011111000: data <= 19'h7fe88; 
        10'b0011111001: data <= 19'h7ff4d; 
        10'b0011111010: data <= 19'h000d0; 
        10'b0011111011: data <= 19'h0013f; 
        10'b0011111100: data <= 19'h000a5; 
        10'b0011111101: data <= 19'h00135; 
        10'b0011111110: data <= 19'h0019f; 
        10'b0011111111: data <= 19'h0036d; 
        10'b0100000000: data <= 19'h004b7; 
        10'b0100000001: data <= 19'h0055b; 
        10'b0100000010: data <= 19'h001f7; 
        10'b0100000011: data <= 19'h0029d; 
        10'b0100000100: data <= 19'h002f6; 
        10'b0100000101: data <= 19'h001f5; 
        10'b0100000110: data <= 19'h004cd; 
        10'b0100000111: data <= 19'h005e1; 
        10'b0100001000: data <= 19'h0077f; 
        10'b0100001001: data <= 19'h00619; 
        10'b0100001010: data <= 19'h008bd; 
        10'b0100001011: data <= 19'h00ac2; 
        10'b0100001100: data <= 19'h009e9; 
        10'b0100001101: data <= 19'h00b0f; 
        10'b0100001110: data <= 19'h00738; 
        10'b0100001111: data <= 19'h0075a; 
        10'b0100010000: data <= 19'h0062f; 
        10'b0100010001: data <= 19'h00528; 
        10'b0100010010: data <= 19'h00271; 
        10'b0100010011: data <= 19'h7ff1d; 
        10'b0100010100: data <= 19'h7fe80; 
        10'b0100010101: data <= 19'h7ff44; 
        10'b0100010110: data <= 19'h000a7; 
        10'b0100010111: data <= 19'h7ffaa; 
        10'b0100011000: data <= 19'h00040; 
        10'b0100011001: data <= 19'h00151; 
        10'b0100011010: data <= 19'h00176; 
        10'b0100011011: data <= 19'h00442; 
        10'b0100011100: data <= 19'h004e1; 
        10'b0100011101: data <= 19'h0040e; 
        10'b0100011110: data <= 19'h000bf; 
        10'b0100011111: data <= 19'h00138; 
        10'b0100100000: data <= 19'h7fe5c; 
        10'b0100100001: data <= 19'h7fff0; 
        10'b0100100010: data <= 19'h002fa; 
        10'b0100100011: data <= 19'h0053e; 
        10'b0100100100: data <= 19'h003a5; 
        10'b0100100101: data <= 19'h0087c; 
        10'b0100100110: data <= 19'h00aeb; 
        10'b0100100111: data <= 19'h00d69; 
        10'b0100101000: data <= 19'h00f45; 
        10'b0100101001: data <= 19'h00b51; 
        10'b0100101010: data <= 19'h008ea; 
        10'b0100101011: data <= 19'h00945; 
        10'b0100101100: data <= 19'h00823; 
        10'b0100101101: data <= 19'h006eb; 
        10'b0100101110: data <= 19'h0030f; 
        10'b0100101111: data <= 19'h7fec0; 
        10'b0100110000: data <= 19'h7fdef; 
        10'b0100110001: data <= 19'h7ff2a; 
        10'b0100110010: data <= 19'h00028; 
        10'b0100110011: data <= 19'h7ffb0; 
        10'b0100110100: data <= 19'h00128; 
        10'b0100110101: data <= 19'h000d0; 
        10'b0100110110: data <= 19'h0017a; 
        10'b0100110111: data <= 19'h0045d; 
        10'b0100111000: data <= 19'h00542; 
        10'b0100111001: data <= 19'h0029b; 
        10'b0100111010: data <= 19'h000f2; 
        10'b0100111011: data <= 19'h000d9; 
        10'b0100111100: data <= 19'h0003e; 
        10'b0100111101: data <= 19'h00328; 
        10'b0100111110: data <= 19'h001a1; 
        10'b0100111111: data <= 19'h0020e; 
        10'b0101000000: data <= 19'h00365; 
        10'b0101000001: data <= 19'h0035d; 
        10'b0101000010: data <= 19'h0037f; 
        10'b0101000011: data <= 19'h00a43; 
        10'b0101000100: data <= 19'h00d54; 
        10'b0101000101: data <= 19'h008e2; 
        10'b0101000110: data <= 19'h008f8; 
        10'b0101000111: data <= 19'h006e5; 
        10'b0101001000: data <= 19'h006b3; 
        10'b0101001001: data <= 19'h00437; 
        10'b0101001010: data <= 19'h0030b; 
        10'b0101001011: data <= 19'h7fef1; 
        10'b0101001100: data <= 19'h7fcec; 
        10'b0101001101: data <= 19'h7ffea; 
        10'b0101001110: data <= 19'h0004b; 
        10'b0101001111: data <= 19'h00159; 
        10'b0101010000: data <= 19'h00108; 
        10'b0101010001: data <= 19'h7ffed; 
        10'b0101010010: data <= 19'h000bc; 
        10'b0101010011: data <= 19'h002bf; 
        10'b0101010100: data <= 19'h00316; 
        10'b0101010101: data <= 19'h00082; 
        10'b0101010110: data <= 19'h000b0; 
        10'b0101010111: data <= 19'h002ef; 
        10'b0101011000: data <= 19'h00203; 
        10'b0101011001: data <= 19'h7ffe2; 
        10'b0101011010: data <= 19'h7fd9a; 
        10'b0101011011: data <= 19'h7f99c; 
        10'b0101011100: data <= 19'h7f27e; 
        10'b0101011101: data <= 19'h7eb18; 
        10'b0101011110: data <= 19'h7f05a; 
        10'b0101011111: data <= 19'h00057; 
        10'b0101100000: data <= 19'h008d7; 
        10'b0101100001: data <= 19'h00806; 
        10'b0101100010: data <= 19'h00328; 
        10'b0101100011: data <= 19'h00122; 
        10'b0101100100: data <= 19'h00036; 
        10'b0101100101: data <= 19'h7fed8; 
        10'b0101100110: data <= 19'h7fef3; 
        10'b0101100111: data <= 19'h7fe1c; 
        10'b0101101000: data <= 19'h7fea3; 
        10'b0101101001: data <= 19'h00146; 
        10'b0101101010: data <= 19'h000e5; 
        10'b0101101011: data <= 19'h00003; 
        10'b0101101100: data <= 19'h0011e; 
        10'b0101101101: data <= 19'h000a8; 
        10'b0101101110: data <= 19'h00134; 
        10'b0101101111: data <= 19'h0027e; 
        10'b0101110000: data <= 19'h000ee; 
        10'b0101110001: data <= 19'h00066; 
        10'b0101110010: data <= 19'h7ff2e; 
        10'b0101110011: data <= 19'h00089; 
        10'b0101110100: data <= 19'h7ffa0; 
        10'b0101110101: data <= 19'h7fdf4; 
        10'b0101110110: data <= 19'h7f94c; 
        10'b0101110111: data <= 19'h7f1dd; 
        10'b0101111000: data <= 19'h7e72f; 
        10'b0101111001: data <= 19'h7e448; 
        10'b0101111010: data <= 19'h7f12b; 
        10'b0101111011: data <= 19'h7fe0e; 
        10'b0101111100: data <= 19'h00483; 
        10'b0101111101: data <= 19'h002e9; 
        10'b0101111110: data <= 19'h000a1; 
        10'b0101111111: data <= 19'h00153; 
        10'b0110000000: data <= 19'h7fd48; 
        10'b0110000001: data <= 19'h7fc86; 
        10'b0110000010: data <= 19'h7ff2f; 
        10'b0110000011: data <= 19'h00042; 
        10'b0110000100: data <= 19'h7ff57; 
        10'b0110000101: data <= 19'h7ff79; 
        10'b0110000110: data <= 19'h000b5; 
        10'b0110000111: data <= 19'h7ff50; 
        10'b0110001000: data <= 19'h7ffb3; 
        10'b0110001001: data <= 19'h00098; 
        10'b0110001010: data <= 19'h0023b; 
        10'b0110001011: data <= 19'h002c8; 
        10'b0110001100: data <= 19'h001c3; 
        10'b0110001101: data <= 19'h0020c; 
        10'b0110001110: data <= 19'h7ff52; 
        10'b0110001111: data <= 19'h7fe93; 
        10'b0110010000: data <= 19'h7fcdb; 
        10'b0110010001: data <= 19'h7f8a1; 
        10'b0110010010: data <= 19'h7f52b; 
        10'b0110010011: data <= 19'h7ef3e; 
        10'b0110010100: data <= 19'h7ea85; 
        10'b0110010101: data <= 19'h7ede2; 
        10'b0110010110: data <= 19'h7f95c; 
        10'b0110010111: data <= 19'h00027; 
        10'b0110011000: data <= 19'h00161; 
        10'b0110011001: data <= 19'h002dc; 
        10'b0110011010: data <= 19'h00836; 
        10'b0110011011: data <= 19'h008d3; 
        10'b0110011100: data <= 19'h0054f; 
        10'b0110011101: data <= 19'h00364; 
        10'b0110011110: data <= 19'h00369; 
        10'b0110011111: data <= 19'h002f5; 
        10'b0110100000: data <= 19'h00100; 
        10'b0110100001: data <= 19'h0004c; 
        10'b0110100010: data <= 19'h7ff87; 
        10'b0110100011: data <= 19'h7ff92; 
        10'b0110100100: data <= 19'h000b8; 
        10'b0110100101: data <= 19'h00110; 
        10'b0110100110: data <= 19'h00064; 
        10'b0110100111: data <= 19'h0010d; 
        10'b0110101000: data <= 19'h0010d; 
        10'b0110101001: data <= 19'h7fd07; 
        10'b0110101010: data <= 19'h7fead; 
        10'b0110101011: data <= 19'h7fe28; 
        10'b0110101100: data <= 19'h7f817; 
        10'b0110101101: data <= 19'h7f667; 
        10'b0110101110: data <= 19'h7f33e; 
        10'b0110101111: data <= 19'h7f162; 
        10'b0110110000: data <= 19'h7f013; 
        10'b0110110001: data <= 19'h7f444; 
        10'b0110110010: data <= 19'h7f925; 
        10'b0110110011: data <= 19'h00036; 
        10'b0110110100: data <= 19'h000bf; 
        10'b0110110101: data <= 19'h00b2b; 
        10'b0110110110: data <= 19'h00d13; 
        10'b0110110111: data <= 19'h00ac6; 
        10'b0110111000: data <= 19'h00991; 
        10'b0110111001: data <= 19'h0083b; 
        10'b0110111010: data <= 19'h00552; 
        10'b0110111011: data <= 19'h00267; 
        10'b0110111100: data <= 19'h7ffe7; 
        10'b0110111101: data <= 19'h7ff56; 
        10'b0110111110: data <= 19'h0002d; 
        10'b0110111111: data <= 19'h00125; 
        10'b0111000000: data <= 19'h000b6; 
        10'b0111000001: data <= 19'h0016b; 
        10'b0111000010: data <= 19'h7ffe2; 
        10'b0111000011: data <= 19'h0017d; 
        10'b0111000100: data <= 19'h0012c; 
        10'b0111000101: data <= 19'h7feab; 
        10'b0111000110: data <= 19'h7fe1e; 
        10'b0111000111: data <= 19'h7ffbb; 
        10'b0111001000: data <= 19'h7f9a2; 
        10'b0111001001: data <= 19'h7f8d0; 
        10'b0111001010: data <= 19'h7f46e; 
        10'b0111001011: data <= 19'h7f23e; 
        10'b0111001100: data <= 19'h7f760; 
        10'b0111001101: data <= 19'h7fb2d; 
        10'b0111001110: data <= 19'h7f902; 
        10'b0111001111: data <= 19'h00399; 
        10'b0111010000: data <= 19'h0045a; 
        10'b0111010001: data <= 19'h00973; 
        10'b0111010010: data <= 19'h00818; 
        10'b0111010011: data <= 19'h0087b; 
        10'b0111010100: data <= 19'h006bf; 
        10'b0111010101: data <= 19'h00524; 
        10'b0111010110: data <= 19'h00103; 
        10'b0111010111: data <= 19'h7fde3; 
        10'b0111011000: data <= 19'h7feb0; 
        10'b0111011001: data <= 19'h7ff41; 
        10'b0111011010: data <= 19'h000ce; 
        10'b0111011011: data <= 19'h00166; 
        10'b0111011100: data <= 19'h0000b; 
        10'b0111011101: data <= 19'h0002e; 
        10'b0111011110: data <= 19'h000dc; 
        10'b0111011111: data <= 19'h7fff1; 
        10'b0111100000: data <= 19'h00048; 
        10'b0111100001: data <= 19'h7ff26; 
        10'b0111100010: data <= 19'h7fbb5; 
        10'b0111100011: data <= 19'h7fa58; 
        10'b0111100100: data <= 19'h7f8e7; 
        10'b0111100101: data <= 19'h7fa24; 
        10'b0111100110: data <= 19'h7f83c; 
        10'b0111100111: data <= 19'h7fa3d; 
        10'b0111101000: data <= 19'h7fe29; 
        10'b0111101001: data <= 19'h00170; 
        10'b0111101010: data <= 19'h000d1; 
        10'b0111101011: data <= 19'h0016e; 
        10'b0111101100: data <= 19'h7ff27; 
        10'b0111101101: data <= 19'h00245; 
        10'b0111101110: data <= 19'h00206; 
        10'b0111101111: data <= 19'h00170; 
        10'b0111110000: data <= 19'h000c3; 
        10'b0111110001: data <= 19'h7fed3; 
        10'b0111110010: data <= 19'h7fd64; 
        10'b0111110011: data <= 19'h7fed3; 
        10'b0111110100: data <= 19'h7fefb; 
        10'b0111110101: data <= 19'h7ff33; 
        10'b0111110110: data <= 19'h7ff92; 
        10'b0111110111: data <= 19'h7ff9d; 
        10'b0111111000: data <= 19'h7ff9b; 
        10'b0111111001: data <= 19'h7ffdf; 
        10'b0111111010: data <= 19'h000f9; 
        10'b0111111011: data <= 19'h0004d; 
        10'b0111111100: data <= 19'h7fe43; 
        10'b0111111101: data <= 19'h7fbde; 
        10'b0111111110: data <= 19'h7f92c; 
        10'b0111111111: data <= 19'h7f77f; 
        10'b1000000000: data <= 19'h7f81b; 
        10'b1000000001: data <= 19'h7f89c; 
        10'b1000000010: data <= 19'h7f682; 
        10'b1000000011: data <= 19'h7fcbc; 
        10'b1000000100: data <= 19'h7ff04; 
        10'b1000000101: data <= 19'h0001e; 
        10'b1000000110: data <= 19'h002ac; 
        10'b1000000111: data <= 19'h7fd2e; 
        10'b1000001000: data <= 19'h7fc8a; 
        10'b1000001001: data <= 19'h7fe16; 
        10'b1000001010: data <= 19'h7fba4; 
        10'b1000001011: data <= 19'h7fd53; 
        10'b1000001100: data <= 19'h7fb82; 
        10'b1000001101: data <= 19'h7f91a; 
        10'b1000001110: data <= 19'h7faf4; 
        10'b1000001111: data <= 19'h7fcd0; 
        10'b1000010000: data <= 19'h7fd7e; 
        10'b1000010001: data <= 19'h00042; 
        10'b1000010010: data <= 19'h7ffb9; 
        10'b1000010011: data <= 19'h0000f; 
        10'b1000010100: data <= 19'h0015a; 
        10'b1000010101: data <= 19'h00173; 
        10'b1000010110: data <= 19'h00153; 
        10'b1000010111: data <= 19'h000a9; 
        10'b1000011000: data <= 19'h7fed4; 
        10'b1000011001: data <= 19'h7faa0; 
        10'b1000011010: data <= 19'h7f765; 
        10'b1000011011: data <= 19'h7f6c5; 
        10'b1000011100: data <= 19'h7f686; 
        10'b1000011101: data <= 19'h7f677; 
        10'b1000011110: data <= 19'h7f98b; 
        10'b1000011111: data <= 19'h7fb5a; 
        10'b1000100000: data <= 19'h7fd38; 
        10'b1000100001: data <= 19'h00135; 
        10'b1000100010: data <= 19'h003c7; 
        10'b1000100011: data <= 19'h7fc0e; 
        10'b1000100100: data <= 19'h7fc27; 
        10'b1000100101: data <= 19'h7fb24; 
        10'b1000100110: data <= 19'h7f847; 
        10'b1000100111: data <= 19'h7f8af; 
        10'b1000101000: data <= 19'h7f6fd; 
        10'b1000101001: data <= 19'h7f7ae; 
        10'b1000101010: data <= 19'h7f9ab; 
        10'b1000101011: data <= 19'h7fba3; 
        10'b1000101100: data <= 19'h7fdca; 
        10'b1000101101: data <= 19'h7ff2e; 
        10'b1000101110: data <= 19'h00163; 
        10'b1000101111: data <= 19'h7ff5f; 
        10'b1000110000: data <= 19'h7ff47; 
        10'b1000110001: data <= 19'h7ffac; 
        10'b1000110010: data <= 19'h00092; 
        10'b1000110011: data <= 19'h7ffc4; 
        10'b1000110100: data <= 19'h7fea4; 
        10'b1000110101: data <= 19'h7fbda; 
        10'b1000110110: data <= 19'h7f755; 
        10'b1000110111: data <= 19'h7f6f5; 
        10'b1000111000: data <= 19'h7f779; 
        10'b1000111001: data <= 19'h7f7ac; 
        10'b1000111010: data <= 19'h7fa31; 
        10'b1000111011: data <= 19'h7fa02; 
        10'b1000111100: data <= 19'h0006f; 
        10'b1000111101: data <= 19'h00098; 
        10'b1000111110: data <= 19'h00201; 
        10'b1000111111: data <= 19'h7fab7; 
        10'b1001000000: data <= 19'h7f965; 
        10'b1001000001: data <= 19'h7f75f; 
        10'b1001000010: data <= 19'h7f416; 
        10'b1001000011: data <= 19'h7f86b; 
        10'b1001000100: data <= 19'h7f58f; 
        10'b1001000101: data <= 19'h7f809; 
        10'b1001000110: data <= 19'h7fa3d; 
        10'b1001000111: data <= 19'h7fd8d; 
        10'b1001001000: data <= 19'h7fe5d; 
        10'b1001001001: data <= 19'h0013c; 
        10'b1001001010: data <= 19'h0012c; 
        10'b1001001011: data <= 19'h000cc; 
        10'b1001001100: data <= 19'h0011d; 
        10'b1001001101: data <= 19'h0012b; 
        10'b1001001110: data <= 19'h00043; 
        10'b1001001111: data <= 19'h7fe7a; 
        10'b1001010000: data <= 19'h7ff3a; 
        10'b1001010001: data <= 19'h7fc4e; 
        10'b1001010010: data <= 19'h7fbab; 
        10'b1001010011: data <= 19'h7f9c1; 
        10'b1001010100: data <= 19'h7fa60; 
        10'b1001010101: data <= 19'h7fca7; 
        10'b1001010110: data <= 19'h7fb3d; 
        10'b1001010111: data <= 19'h7fc1e; 
        10'b1001011000: data <= 19'h7fe44; 
        10'b1001011001: data <= 19'h0003c; 
        10'b1001011010: data <= 19'h7fef5; 
        10'b1001011011: data <= 19'h7fc70; 
        10'b1001011100: data <= 19'h7fbe7; 
        10'b1001011101: data <= 19'h7f77d; 
        10'b1001011110: data <= 19'h7f785; 
        10'b1001011111: data <= 19'h7f781; 
        10'b1001100000: data <= 19'h7f70d; 
        10'b1001100001: data <= 19'h7f86c; 
        10'b1001100010: data <= 19'h7fb8d; 
        10'b1001100011: data <= 19'h7fca2; 
        10'b1001100100: data <= 19'h7ffda; 
        10'b1001100101: data <= 19'h00085; 
        10'b1001100110: data <= 19'h00120; 
        10'b1001100111: data <= 19'h7ffc2; 
        10'b1001101000: data <= 19'h00061; 
        10'b1001101001: data <= 19'h00016; 
        10'b1001101010: data <= 19'h0004c; 
        10'b1001101011: data <= 19'h7ff10; 
        10'b1001101100: data <= 19'h7ff93; 
        10'b1001101101: data <= 19'h0008d; 
        10'b1001101110: data <= 19'h7fea5; 
        10'b1001101111: data <= 19'h000ac; 
        10'b1001110000: data <= 19'h00112; 
        10'b1001110001: data <= 19'h7fe4a; 
        10'b1001110010: data <= 19'h7fcbe; 
        10'b1001110011: data <= 19'h7fa71; 
        10'b1001110100: data <= 19'h7face; 
        10'b1001110101: data <= 19'h7fde8; 
        10'b1001110110: data <= 19'h0009f; 
        10'b1001110111: data <= 19'h0009d; 
        10'b1001111000: data <= 19'h7fcc5; 
        10'b1001111001: data <= 19'h7fc00; 
        10'b1001111010: data <= 19'h7f930; 
        10'b1001111011: data <= 19'h7f930; 
        10'b1001111100: data <= 19'h7f853; 
        10'b1001111101: data <= 19'h7f948; 
        10'b1001111110: data <= 19'h7fc96; 
        10'b1001111111: data <= 19'h7fed9; 
        10'b1010000000: data <= 19'h000be; 
        10'b1010000001: data <= 19'h7ff46; 
        10'b1010000010: data <= 19'h0005b; 
        10'b1010000011: data <= 19'h00006; 
        10'b1010000100: data <= 19'h00086; 
        10'b1010000101: data <= 19'h00110; 
        10'b1010000110: data <= 19'h7ff2e; 
        10'b1010000111: data <= 19'h7ff41; 
        10'b1010001000: data <= 19'h00168; 
        10'b1010001001: data <= 19'h001e2; 
        10'b1010001010: data <= 19'h00419; 
        10'b1010001011: data <= 19'h00577; 
        10'b1010001100: data <= 19'h0029c; 
        10'b1010001101: data <= 19'h00085; 
        10'b1010001110: data <= 19'h7fe64; 
        10'b1010001111: data <= 19'h7fc49; 
        10'b1010010000: data <= 19'h7fcf6; 
        10'b1010010001: data <= 19'h00036; 
        10'b1010010010: data <= 19'h00221; 
        10'b1010010011: data <= 19'h001f6; 
        10'b1010010100: data <= 19'h7ff2e; 
        10'b1010010101: data <= 19'h7fec9; 
        10'b1010010110: data <= 19'h7fba4; 
        10'b1010010111: data <= 19'h7f9eb; 
        10'b1010011000: data <= 19'h7f9c7; 
        10'b1010011001: data <= 19'h7fb24; 
        10'b1010011010: data <= 19'h7fbfe; 
        10'b1010011011: data <= 19'h7fd63; 
        10'b1010011100: data <= 19'h7fed9; 
        10'b1010011101: data <= 19'h00016; 
        10'b1010011110: data <= 19'h00013; 
        10'b1010011111: data <= 19'h7ff92; 
        10'b1010100000: data <= 19'h7fffd; 
        10'b1010100001: data <= 19'h7ffdb; 
        10'b1010100010: data <= 19'h00064; 
        10'b1010100011: data <= 19'h000ea; 
        10'b1010100100: data <= 19'h001f5; 
        10'b1010100101: data <= 19'h00480; 
        10'b1010100110: data <= 19'h006cf; 
        10'b1010100111: data <= 19'h007ac; 
        10'b1010101000: data <= 19'h00684; 
        10'b1010101001: data <= 19'h0035c; 
        10'b1010101010: data <= 19'h0073d; 
        10'b1010101011: data <= 19'h00446; 
        10'b1010101100: data <= 19'h003b5; 
        10'b1010101101: data <= 19'h00539; 
        10'b1010101110: data <= 19'h00337; 
        10'b1010101111: data <= 19'h004a4; 
        10'b1010110000: data <= 19'h002bf; 
        10'b1010110001: data <= 19'h00225; 
        10'b1010110010: data <= 19'h7ffdd; 
        10'b1010110011: data <= 19'h7fe00; 
        10'b1010110100: data <= 19'h7fde0; 
        10'b1010110101: data <= 19'h7fd6c; 
        10'b1010110110: data <= 19'h7fd16; 
        10'b1010110111: data <= 19'h7fd59; 
        10'b1010111000: data <= 19'h00068; 
        10'b1010111001: data <= 19'h7ffca; 
        10'b1010111010: data <= 19'h7ff4e; 
        10'b1010111011: data <= 19'h000cb; 
        10'b1010111100: data <= 19'h7ff4b; 
        10'b1010111101: data <= 19'h000a6; 
        10'b1010111110: data <= 19'h0012c; 
        10'b1010111111: data <= 19'h00119; 
        10'b1011000000: data <= 19'h000a3; 
        10'b1011000001: data <= 19'h0023e; 
        10'b1011000010: data <= 19'h00352; 
        10'b1011000011: data <= 19'h00521; 
        10'b1011000100: data <= 19'h007ee; 
        10'b1011000101: data <= 19'h007be; 
        10'b1011000110: data <= 19'h0092a; 
        10'b1011000111: data <= 19'h00888; 
        10'b1011001000: data <= 19'h0079a; 
        10'b1011001001: data <= 19'h00605; 
        10'b1011001010: data <= 19'h00626; 
        10'b1011001011: data <= 19'h00684; 
        10'b1011001100: data <= 19'h00576; 
        10'b1011001101: data <= 19'h0051b; 
        10'b1011001110: data <= 19'h0041d; 
        10'b1011001111: data <= 19'h00169; 
        10'b1011010000: data <= 19'h7fe44; 
        10'b1011010001: data <= 19'h0003c; 
        10'b1011010010: data <= 19'h7ff25; 
        10'b1011010011: data <= 19'h7ff5f; 
        10'b1011010100: data <= 19'h7ffcd; 
        10'b1011010101: data <= 19'h00064; 
        10'b1011010110: data <= 19'h0018e; 
        10'b1011010111: data <= 19'h00102; 
        10'b1011011000: data <= 19'h7ff73; 
        10'b1011011001: data <= 19'h0004c; 
        10'b1011011010: data <= 19'h00178; 
        10'b1011011011: data <= 19'h7ffc0; 
        10'b1011011100: data <= 19'h7ff80; 
        10'b1011011101: data <= 19'h0015f; 
        10'b1011011110: data <= 19'h00019; 
        10'b1011011111: data <= 19'h00141; 
        10'b1011100000: data <= 19'h00132; 
        10'b1011100001: data <= 19'h0002b; 
        10'b1011100010: data <= 19'h001ba; 
        10'b1011100011: data <= 19'h0028b; 
        10'b1011100100: data <= 19'h000bc; 
        10'b1011100101: data <= 19'h0022f; 
        10'b1011100110: data <= 19'h004ae; 
        10'b1011100111: data <= 19'h005c7; 
        10'b1011101000: data <= 19'h0048f; 
        10'b1011101001: data <= 19'h005d7; 
        10'b1011101010: data <= 19'h00354; 
        10'b1011101011: data <= 19'h00192; 
        10'b1011101100: data <= 19'h0000d; 
        10'b1011101101: data <= 19'h0009b; 
        10'b1011101110: data <= 19'h7ffd6; 
        10'b1011101111: data <= 19'h00056; 
        10'b1011110000: data <= 19'h00011; 
        10'b1011110001: data <= 19'h7ff9c; 
        10'b1011110010: data <= 19'h7ffe8; 
        10'b1011110011: data <= 19'h7ffce; 
        10'b1011110100: data <= 19'h7ff46; 
        10'b1011110101: data <= 19'h00098; 
        10'b1011110110: data <= 19'h00067; 
        10'b1011110111: data <= 19'h000bd; 
        10'b1011111000: data <= 19'h00101; 
        10'b1011111001: data <= 19'h00099; 
        10'b1011111010: data <= 19'h00042; 
        10'b1011111011: data <= 19'h0001c; 
        10'b1011111100: data <= 19'h001a5; 
        10'b1011111101: data <= 19'h00102; 
        10'b1011111110: data <= 19'h0004c; 
        10'b1011111111: data <= 19'h00104; 
        10'b1100000000: data <= 19'h0007e; 
        10'b1100000001: data <= 19'h001e6; 
        10'b1100000010: data <= 19'h00122; 
        10'b1100000011: data <= 19'h000dd; 
        10'b1100000100: data <= 19'h002a4; 
        10'b1100000101: data <= 19'h000e5; 
        10'b1100000110: data <= 19'h000cb; 
        10'b1100000111: data <= 19'h001d5; 
        10'b1100001000: data <= 19'h00038; 
        10'b1100001001: data <= 19'h7ffb1; 
        10'b1100001010: data <= 19'h0017f; 
        10'b1100001011: data <= 19'h000d2; 
        10'b1100001100: data <= 19'h00061; 
        10'b1100001101: data <= 19'h7ffba; 
        10'b1100001110: data <= 19'h7ff63; 
        10'b1100001111: data <= 19'h000ff; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 14) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 20'h00030; 
        10'b0000000001: data <= 20'h00041; 
        10'b0000000010: data <= 20'h001e6; 
        10'b0000000011: data <= 20'h000bb; 
        10'b0000000100: data <= 20'h00318; 
        10'b0000000101: data <= 20'hffea0; 
        10'b0000000110: data <= 20'hfff15; 
        10'b0000000111: data <= 20'h00101; 
        10'b0000001000: data <= 20'h00261; 
        10'b0000001001: data <= 20'h00255; 
        10'b0000001010: data <= 20'hffeaf; 
        10'b0000001011: data <= 20'h0009f; 
        10'b0000001100: data <= 20'h000ac; 
        10'b0000001101: data <= 20'hfffa6; 
        10'b0000001110: data <= 20'h0027d; 
        10'b0000001111: data <= 20'h000ab; 
        10'b0000010000: data <= 20'h0000d; 
        10'b0000010001: data <= 20'hfffea; 
        10'b0000010010: data <= 20'h00043; 
        10'b0000010011: data <= 20'h000dd; 
        10'b0000010100: data <= 20'h0019a; 
        10'b0000010101: data <= 20'h00307; 
        10'b0000010110: data <= 20'hfff30; 
        10'b0000010111: data <= 20'h0023a; 
        10'b0000011000: data <= 20'hfffb1; 
        10'b0000011001: data <= 20'h00199; 
        10'b0000011010: data <= 20'hfffdf; 
        10'b0000011011: data <= 20'hffffe; 
        10'b0000011100: data <= 20'h002da; 
        10'b0000011101: data <= 20'hfff64; 
        10'b0000011110: data <= 20'h000a4; 
        10'b0000011111: data <= 20'h002d0; 
        10'b0000100000: data <= 20'h00114; 
        10'b0000100001: data <= 20'h0001a; 
        10'b0000100010: data <= 20'h002cb; 
        10'b0000100011: data <= 20'h000e1; 
        10'b0000100100: data <= 20'h00045; 
        10'b0000100101: data <= 20'hfff86; 
        10'b0000100110: data <= 20'hfffa1; 
        10'b0000100111: data <= 20'hffe88; 
        10'b0000101000: data <= 20'h00267; 
        10'b0000101001: data <= 20'hfffd3; 
        10'b0000101010: data <= 20'h002e2; 
        10'b0000101011: data <= 20'hfff40; 
        10'b0000101100: data <= 20'h00140; 
        10'b0000101101: data <= 20'h0022a; 
        10'b0000101110: data <= 20'h00270; 
        10'b0000101111: data <= 20'h001f2; 
        10'b0000110000: data <= 20'h00010; 
        10'b0000110001: data <= 20'h001ea; 
        10'b0000110010: data <= 20'hffff1; 
        10'b0000110011: data <= 20'h0030a; 
        10'b0000110100: data <= 20'h00258; 
        10'b0000110101: data <= 20'hfff28; 
        10'b0000110110: data <= 20'hfff2d; 
        10'b0000110111: data <= 20'h0013d; 
        10'b0000111000: data <= 20'h002b4; 
        10'b0000111001: data <= 20'h002aa; 
        10'b0000111010: data <= 20'h00218; 
        10'b0000111011: data <= 20'hfff9d; 
        10'b0000111100: data <= 20'h0026e; 
        10'b0000111101: data <= 20'hffed8; 
        10'b0000111110: data <= 20'hfff0d; 
        10'b0000111111: data <= 20'h001e7; 
        10'b0001000000: data <= 20'h0019a; 
        10'b0001000001: data <= 20'hfff0f; 
        10'b0001000010: data <= 20'hfffcb; 
        10'b0001000011: data <= 20'h0012f; 
        10'b0001000100: data <= 20'hfffac; 
        10'b0001000101: data <= 20'hfff61; 
        10'b0001000110: data <= 20'h000be; 
        10'b0001000111: data <= 20'h00272; 
        10'b0001001000: data <= 20'h001f9; 
        10'b0001001001: data <= 20'h0005e; 
        10'b0001001010: data <= 20'h000f8; 
        10'b0001001011: data <= 20'h002c3; 
        10'b0001001100: data <= 20'h00258; 
        10'b0001001101: data <= 20'h002b7; 
        10'b0001001110: data <= 20'hffea3; 
        10'b0001001111: data <= 20'h0021d; 
        10'b0001010000: data <= 20'h000cd; 
        10'b0001010001: data <= 20'h001de; 
        10'b0001010010: data <= 20'h0019c; 
        10'b0001010011: data <= 20'h00261; 
        10'b0001010100: data <= 20'hfffc8; 
        10'b0001010101: data <= 20'h00029; 
        10'b0001010110: data <= 20'h0027a; 
        10'b0001010111: data <= 20'hfffa0; 
        10'b0001011000: data <= 20'h00047; 
        10'b0001011001: data <= 20'hfffd5; 
        10'b0001011010: data <= 20'hfff17; 
        10'b0001011011: data <= 20'h0019c; 
        10'b0001011100: data <= 20'h00003; 
        10'b0001011101: data <= 20'h0019c; 
        10'b0001011110: data <= 20'hffead; 
        10'b0001011111: data <= 20'h00054; 
        10'b0001100000: data <= 20'h0014c; 
        10'b0001100001: data <= 20'hffe37; 
        10'b0001100010: data <= 20'h00178; 
        10'b0001100011: data <= 20'hffeca; 
        10'b0001100100: data <= 20'hffd61; 
        10'b0001100101: data <= 20'hffdda; 
        10'b0001100110: data <= 20'hffe28; 
        10'b0001100111: data <= 20'hffec3; 
        10'b0001101000: data <= 20'hfffb1; 
        10'b0001101001: data <= 20'hffedd; 
        10'b0001101010: data <= 20'h000ff; 
        10'b0001101011: data <= 20'hfffdf; 
        10'b0001101100: data <= 20'h00133; 
        10'b0001101101: data <= 20'h0030c; 
        10'b0001101110: data <= 20'hfff00; 
        10'b0001101111: data <= 20'h00142; 
        10'b0001110000: data <= 20'h002f5; 
        10'b0001110001: data <= 20'hffeed; 
        10'b0001110010: data <= 20'h001a6; 
        10'b0001110011: data <= 20'hffebf; 
        10'b0001110100: data <= 20'h000b1; 
        10'b0001110101: data <= 20'hfff6e; 
        10'b0001110110: data <= 20'h00022; 
        10'b0001110111: data <= 20'hffec9; 
        10'b0001111000: data <= 20'h000eb; 
        10'b0001111001: data <= 20'hfff91; 
        10'b0001111010: data <= 20'hffd1b; 
        10'b0001111011: data <= 20'hffa6c; 
        10'b0001111100: data <= 20'hffa23; 
        10'b0001111101: data <= 20'hffa68; 
        10'b0001111110: data <= 20'hff955; 
        10'b0001111111: data <= 20'hff505; 
        10'b0010000000: data <= 20'hff985; 
        10'b0010000001: data <= 20'hffb1f; 
        10'b0010000010: data <= 20'hffbc2; 
        10'b0010000011: data <= 20'hffedb; 
        10'b0010000100: data <= 20'hffcd6; 
        10'b0010000101: data <= 20'h0017a; 
        10'b0010000110: data <= 20'h0003a; 
        10'b0010000111: data <= 20'hffe76; 
        10'b0010001000: data <= 20'h002cd; 
        10'b0010001001: data <= 20'hfffe7; 
        10'b0010001010: data <= 20'h002be; 
        10'b0010001011: data <= 20'h002a9; 
        10'b0010001100: data <= 20'h00285; 
        10'b0010001101: data <= 20'h0001a; 
        10'b0010001110: data <= 20'h0026e; 
        10'b0010001111: data <= 20'hfff56; 
        10'b0010010000: data <= 20'hffe19; 
        10'b0010010001: data <= 20'hfffac; 
        10'b0010010010: data <= 20'hffe8b; 
        10'b0010010011: data <= 20'hfff78; 
        10'b0010010100: data <= 20'hffe46; 
        10'b0010010101: data <= 20'hffbfe; 
        10'b0010010110: data <= 20'hff629; 
        10'b0010010111: data <= 20'hff3ed; 
        10'b0010011000: data <= 20'hff0cd; 
        10'b0010011001: data <= 20'hfee32; 
        10'b0010011010: data <= 20'hfe9c9; 
        10'b0010011011: data <= 20'hfe9f3; 
        10'b0010011100: data <= 20'hfe8e1; 
        10'b0010011101: data <= 20'hfeb9a; 
        10'b0010011110: data <= 20'hfeeb7; 
        10'b0010011111: data <= 20'hff2d9; 
        10'b0010100000: data <= 20'hff6a8; 
        10'b0010100001: data <= 20'hffcab; 
        10'b0010100010: data <= 20'hffad9; 
        10'b0010100011: data <= 20'hfff5b; 
        10'b0010100100: data <= 20'h00241; 
        10'b0010100101: data <= 20'h001cd; 
        10'b0010100110: data <= 20'hfff8a; 
        10'b0010100111: data <= 20'h0001a; 
        10'b0010101000: data <= 20'h00218; 
        10'b0010101001: data <= 20'h002de; 
        10'b0010101010: data <= 20'h00034; 
        10'b0010101011: data <= 20'h00077; 
        10'b0010101100: data <= 20'h0031b; 
        10'b0010101101: data <= 20'h003b2; 
        10'b0010101110: data <= 20'h00453; 
        10'b0010101111: data <= 20'h00683; 
        10'b0010110000: data <= 20'h009a9; 
        10'b0010110001: data <= 20'h007bc; 
        10'b0010110010: data <= 20'h0083b; 
        10'b0010110011: data <= 20'h0017b; 
        10'b0010110100: data <= 20'hff966; 
        10'b0010110101: data <= 20'hff224; 
        10'b0010110110: data <= 20'hff18a; 
        10'b0010110111: data <= 20'hff87d; 
        10'b0010111000: data <= 20'hffb70; 
        10'b0010111001: data <= 20'hffa96; 
        10'b0010111010: data <= 20'hff970; 
        10'b0010111011: data <= 20'hff868; 
        10'b0010111100: data <= 20'hff481; 
        10'b0010111101: data <= 20'hffbb0; 
        10'b0010111110: data <= 20'hff7f1; 
        10'b0010111111: data <= 20'hffa23; 
        10'b0011000000: data <= 20'hffc13; 
        10'b0011000001: data <= 20'hffeaf; 
        10'b0011000010: data <= 20'hffea3; 
        10'b0011000011: data <= 20'h00051; 
        10'b0011000100: data <= 20'h001e8; 
        10'b0011000101: data <= 20'h002e4; 
        10'b0011000110: data <= 20'h00261; 
        10'b0011000111: data <= 20'h005a0; 
        10'b0011001000: data <= 20'h006d3; 
        10'b0011001001: data <= 20'h00623; 
        10'b0011001010: data <= 20'h008e3; 
        10'b0011001011: data <= 20'h00d95; 
        10'b0011001100: data <= 20'h0129a; 
        10'b0011001101: data <= 20'h00ebd; 
        10'b0011001110: data <= 20'h00a2b; 
        10'b0011001111: data <= 20'h00b33; 
        10'b0011010000: data <= 20'h00bee; 
        10'b0011010001: data <= 20'h0024b; 
        10'b0011010010: data <= 20'h001b2; 
        10'b0011010011: data <= 20'h00445; 
        10'b0011010100: data <= 20'h00c98; 
        10'b0011010101: data <= 20'h00e00; 
        10'b0011010110: data <= 20'h0097d; 
        10'b0011010111: data <= 20'h0079b; 
        10'b0011011000: data <= 20'h001db; 
        10'b0011011001: data <= 20'hffde5; 
        10'b0011011010: data <= 20'h000fd; 
        10'b0011011011: data <= 20'hffdbb; 
        10'b0011011100: data <= 20'hffde1; 
        10'b0011011101: data <= 20'hfffe3; 
        10'b0011011110: data <= 20'h00180; 
        10'b0011011111: data <= 20'hfff70; 
        10'b0011100000: data <= 20'hffe8a; 
        10'b0011100001: data <= 20'h00308; 
        10'b0011100010: data <= 20'h0012b; 
        10'b0011100011: data <= 20'h004c1; 
        10'b0011100100: data <= 20'h0099f; 
        10'b0011100101: data <= 20'h008ad; 
        10'b0011100110: data <= 20'h00b9e; 
        10'b0011100111: data <= 20'h014db; 
        10'b0011101000: data <= 20'h00e0a; 
        10'b0011101001: data <= 20'h009ac; 
        10'b0011101010: data <= 20'h00c4e; 
        10'b0011101011: data <= 20'h0107b; 
        10'b0011101100: data <= 20'h00faa; 
        10'b0011101101: data <= 20'h007e1; 
        10'b0011101110: data <= 20'h0049b; 
        10'b0011101111: data <= 20'h00665; 
        10'b0011110000: data <= 20'h00b1b; 
        10'b0011110001: data <= 20'h01113; 
        10'b0011110010: data <= 20'h00bb4; 
        10'b0011110011: data <= 20'h00a06; 
        10'b0011110100: data <= 20'h00800; 
        10'b0011110101: data <= 20'h00030; 
        10'b0011110110: data <= 20'h004d9; 
        10'b0011110111: data <= 20'h0041e; 
        10'b0011111000: data <= 20'hffd10; 
        10'b0011111001: data <= 20'hffe99; 
        10'b0011111010: data <= 20'h0019f; 
        10'b0011111011: data <= 20'h0027f; 
        10'b0011111100: data <= 20'h0014a; 
        10'b0011111101: data <= 20'h0026a; 
        10'b0011111110: data <= 20'h0033e; 
        10'b0011111111: data <= 20'h006da; 
        10'b0100000000: data <= 20'h0096e; 
        10'b0100000001: data <= 20'h00ab5; 
        10'b0100000010: data <= 20'h003ee; 
        10'b0100000011: data <= 20'h0053a; 
        10'b0100000100: data <= 20'h005ec; 
        10'b0100000101: data <= 20'h003eb; 
        10'b0100000110: data <= 20'h00999; 
        10'b0100000111: data <= 20'h00bc3; 
        10'b0100001000: data <= 20'h00eff; 
        10'b0100001001: data <= 20'h00c33; 
        10'b0100001010: data <= 20'h0117a; 
        10'b0100001011: data <= 20'h01583; 
        10'b0100001100: data <= 20'h013d1; 
        10'b0100001101: data <= 20'h0161e; 
        10'b0100001110: data <= 20'h00e70; 
        10'b0100001111: data <= 20'h00eb4; 
        10'b0100010000: data <= 20'h00c5e; 
        10'b0100010001: data <= 20'h00a51; 
        10'b0100010010: data <= 20'h004e2; 
        10'b0100010011: data <= 20'hffe39; 
        10'b0100010100: data <= 20'hffcff; 
        10'b0100010101: data <= 20'hffe87; 
        10'b0100010110: data <= 20'h0014e; 
        10'b0100010111: data <= 20'hfff55; 
        10'b0100011000: data <= 20'h00080; 
        10'b0100011001: data <= 20'h002a2; 
        10'b0100011010: data <= 20'h002eb; 
        10'b0100011011: data <= 20'h00885; 
        10'b0100011100: data <= 20'h009c2; 
        10'b0100011101: data <= 20'h0081d; 
        10'b0100011110: data <= 20'h0017f; 
        10'b0100011111: data <= 20'h00271; 
        10'b0100100000: data <= 20'hffcb8; 
        10'b0100100001: data <= 20'hfffe0; 
        10'b0100100010: data <= 20'h005f4; 
        10'b0100100011: data <= 20'h00a7b; 
        10'b0100100100: data <= 20'h0074b; 
        10'b0100100101: data <= 20'h010f9; 
        10'b0100100110: data <= 20'h015d6; 
        10'b0100100111: data <= 20'h01ad2; 
        10'b0100101000: data <= 20'h01e8a; 
        10'b0100101001: data <= 20'h016a2; 
        10'b0100101010: data <= 20'h011d3; 
        10'b0100101011: data <= 20'h0128a; 
        10'b0100101100: data <= 20'h01047; 
        10'b0100101101: data <= 20'h00dd7; 
        10'b0100101110: data <= 20'h0061e; 
        10'b0100101111: data <= 20'hffd81; 
        10'b0100110000: data <= 20'hffbde; 
        10'b0100110001: data <= 20'hffe53; 
        10'b0100110010: data <= 20'h00050; 
        10'b0100110011: data <= 20'hfff60; 
        10'b0100110100: data <= 20'h00251; 
        10'b0100110101: data <= 20'h001a0; 
        10'b0100110110: data <= 20'h002f4; 
        10'b0100110111: data <= 20'h008ba; 
        10'b0100111000: data <= 20'h00a84; 
        10'b0100111001: data <= 20'h00537; 
        10'b0100111010: data <= 20'h001e5; 
        10'b0100111011: data <= 20'h001b3; 
        10'b0100111100: data <= 20'h0007d; 
        10'b0100111101: data <= 20'h00650; 
        10'b0100111110: data <= 20'h00341; 
        10'b0100111111: data <= 20'h0041b; 
        10'b0101000000: data <= 20'h006c9; 
        10'b0101000001: data <= 20'h006b9; 
        10'b0101000010: data <= 20'h006fe; 
        10'b0101000011: data <= 20'h01487; 
        10'b0101000100: data <= 20'h01aa8; 
        10'b0101000101: data <= 20'h011c3; 
        10'b0101000110: data <= 20'h011f0; 
        10'b0101000111: data <= 20'h00dcb; 
        10'b0101001000: data <= 20'h00d67; 
        10'b0101001001: data <= 20'h0086e; 
        10'b0101001010: data <= 20'h00616; 
        10'b0101001011: data <= 20'hffde2; 
        10'b0101001100: data <= 20'hff9d8; 
        10'b0101001101: data <= 20'hfffd4; 
        10'b0101001110: data <= 20'h00097; 
        10'b0101001111: data <= 20'h002b2; 
        10'b0101010000: data <= 20'h00210; 
        10'b0101010001: data <= 20'hfffda; 
        10'b0101010010: data <= 20'h00178; 
        10'b0101010011: data <= 20'h0057f; 
        10'b0101010100: data <= 20'h0062c; 
        10'b0101010101: data <= 20'h00104; 
        10'b0101010110: data <= 20'h00161; 
        10'b0101010111: data <= 20'h005df; 
        10'b0101011000: data <= 20'h00406; 
        10'b0101011001: data <= 20'hfffc4; 
        10'b0101011010: data <= 20'hffb33; 
        10'b0101011011: data <= 20'hff338; 
        10'b0101011100: data <= 20'hfe4fc; 
        10'b0101011101: data <= 20'hfd62f; 
        10'b0101011110: data <= 20'hfe0b3; 
        10'b0101011111: data <= 20'h000ae; 
        10'b0101100000: data <= 20'h011ae; 
        10'b0101100001: data <= 20'h0100b; 
        10'b0101100010: data <= 20'h00650; 
        10'b0101100011: data <= 20'h00245; 
        10'b0101100100: data <= 20'h0006c; 
        10'b0101100101: data <= 20'hffdb0; 
        10'b0101100110: data <= 20'hffde7; 
        10'b0101100111: data <= 20'hffc38; 
        10'b0101101000: data <= 20'hffd47; 
        10'b0101101001: data <= 20'h0028d; 
        10'b0101101010: data <= 20'h001cb; 
        10'b0101101011: data <= 20'h00006; 
        10'b0101101100: data <= 20'h0023c; 
        10'b0101101101: data <= 20'h00151; 
        10'b0101101110: data <= 20'h00269; 
        10'b0101101111: data <= 20'h004fd; 
        10'b0101110000: data <= 20'h001db; 
        10'b0101110001: data <= 20'h000cc; 
        10'b0101110010: data <= 20'hffe5d; 
        10'b0101110011: data <= 20'h00113; 
        10'b0101110100: data <= 20'hfff3f; 
        10'b0101110101: data <= 20'hffbe8; 
        10'b0101110110: data <= 20'hff297; 
        10'b0101110111: data <= 20'hfe3ba; 
        10'b0101111000: data <= 20'hfce5e; 
        10'b0101111001: data <= 20'hfc88f; 
        10'b0101111010: data <= 20'hfe256; 
        10'b0101111011: data <= 20'hffc1c; 
        10'b0101111100: data <= 20'h00906; 
        10'b0101111101: data <= 20'h005d2; 
        10'b0101111110: data <= 20'h00142; 
        10'b0101111111: data <= 20'h002a6; 
        10'b0110000000: data <= 20'hffa91; 
        10'b0110000001: data <= 20'hff90c; 
        10'b0110000010: data <= 20'hffe5e; 
        10'b0110000011: data <= 20'h00083; 
        10'b0110000100: data <= 20'hffeae; 
        10'b0110000101: data <= 20'hffef2; 
        10'b0110000110: data <= 20'h0016a; 
        10'b0110000111: data <= 20'hffea1; 
        10'b0110001000: data <= 20'hfff67; 
        10'b0110001001: data <= 20'h00131; 
        10'b0110001010: data <= 20'h00476; 
        10'b0110001011: data <= 20'h0058f; 
        10'b0110001100: data <= 20'h00386; 
        10'b0110001101: data <= 20'h00418; 
        10'b0110001110: data <= 20'hffea5; 
        10'b0110001111: data <= 20'hffd26; 
        10'b0110010000: data <= 20'hff9b5; 
        10'b0110010001: data <= 20'hff143; 
        10'b0110010010: data <= 20'hfea56; 
        10'b0110010011: data <= 20'hfde7d; 
        10'b0110010100: data <= 20'hfd50b; 
        10'b0110010101: data <= 20'hfdbc3; 
        10'b0110010110: data <= 20'hff2b7; 
        10'b0110010111: data <= 20'h0004f; 
        10'b0110011000: data <= 20'h002c3; 
        10'b0110011001: data <= 20'h005b9; 
        10'b0110011010: data <= 20'h0106b; 
        10'b0110011011: data <= 20'h011a6; 
        10'b0110011100: data <= 20'h00a9e; 
        10'b0110011101: data <= 20'h006c8; 
        10'b0110011110: data <= 20'h006d2; 
        10'b0110011111: data <= 20'h005ea; 
        10'b0110100000: data <= 20'h00200; 
        10'b0110100001: data <= 20'h00098; 
        10'b0110100010: data <= 20'hfff0e; 
        10'b0110100011: data <= 20'hfff24; 
        10'b0110100100: data <= 20'h00171; 
        10'b0110100101: data <= 20'h00220; 
        10'b0110100110: data <= 20'h000c7; 
        10'b0110100111: data <= 20'h0021b; 
        10'b0110101000: data <= 20'h00219; 
        10'b0110101001: data <= 20'hffa0e; 
        10'b0110101010: data <= 20'hffd59; 
        10'b0110101011: data <= 20'hffc51; 
        10'b0110101100: data <= 20'hff02e; 
        10'b0110101101: data <= 20'hfecce; 
        10'b0110101110: data <= 20'hfe67c; 
        10'b0110101111: data <= 20'hfe2c3; 
        10'b0110110000: data <= 20'hfe027; 
        10'b0110110001: data <= 20'hfe887; 
        10'b0110110010: data <= 20'hff24a; 
        10'b0110110011: data <= 20'h0006b; 
        10'b0110110100: data <= 20'h0017f; 
        10'b0110110101: data <= 20'h01655; 
        10'b0110110110: data <= 20'h01a25; 
        10'b0110110111: data <= 20'h0158c; 
        10'b0110111000: data <= 20'h01322; 
        10'b0110111001: data <= 20'h01076; 
        10'b0110111010: data <= 20'h00aa3; 
        10'b0110111011: data <= 20'h004ce; 
        10'b0110111100: data <= 20'hfffcd; 
        10'b0110111101: data <= 20'hffeac; 
        10'b0110111110: data <= 20'h0005b; 
        10'b0110111111: data <= 20'h0024a; 
        10'b0111000000: data <= 20'h0016d; 
        10'b0111000001: data <= 20'h002d5; 
        10'b0111000010: data <= 20'hfffc4; 
        10'b0111000011: data <= 20'h002f9; 
        10'b0111000100: data <= 20'h00257; 
        10'b0111000101: data <= 20'hffd56; 
        10'b0111000110: data <= 20'hffc3c; 
        10'b0111000111: data <= 20'hfff75; 
        10'b0111001000: data <= 20'hff344; 
        10'b0111001001: data <= 20'hff1a0; 
        10'b0111001010: data <= 20'hfe8db; 
        10'b0111001011: data <= 20'hfe47d; 
        10'b0111001100: data <= 20'hfeec1; 
        10'b0111001101: data <= 20'hff65a; 
        10'b0111001110: data <= 20'hff203; 
        10'b0111001111: data <= 20'h00732; 
        10'b0111010000: data <= 20'h008b4; 
        10'b0111010001: data <= 20'h012e5; 
        10'b0111010010: data <= 20'h01030; 
        10'b0111010011: data <= 20'h010f6; 
        10'b0111010100: data <= 20'h00d7f; 
        10'b0111010101: data <= 20'h00a47; 
        10'b0111010110: data <= 20'h00207; 
        10'b0111010111: data <= 20'hffbc5; 
        10'b0111011000: data <= 20'hffd60; 
        10'b0111011001: data <= 20'hffe82; 
        10'b0111011010: data <= 20'h0019b; 
        10'b0111011011: data <= 20'h002cc; 
        10'b0111011100: data <= 20'h00017; 
        10'b0111011101: data <= 20'h0005c; 
        10'b0111011110: data <= 20'h001b8; 
        10'b0111011111: data <= 20'hfffe2; 
        10'b0111100000: data <= 20'h00091; 
        10'b0111100001: data <= 20'hffe4d; 
        10'b0111100010: data <= 20'hff76b; 
        10'b0111100011: data <= 20'hff4b1; 
        10'b0111100100: data <= 20'hff1cf; 
        10'b0111100101: data <= 20'hff449; 
        10'b0111100110: data <= 20'hff078; 
        10'b0111100111: data <= 20'hff47a; 
        10'b0111101000: data <= 20'hffc52; 
        10'b0111101001: data <= 20'h002e0; 
        10'b0111101010: data <= 20'h001a1; 
        10'b0111101011: data <= 20'h002dd; 
        10'b0111101100: data <= 20'hffe4e; 
        10'b0111101101: data <= 20'h0048a; 
        10'b0111101110: data <= 20'h0040c; 
        10'b0111101111: data <= 20'h002e0; 
        10'b0111110000: data <= 20'h00187; 
        10'b0111110001: data <= 20'hffda6; 
        10'b0111110010: data <= 20'hffac7; 
        10'b0111110011: data <= 20'hffda6; 
        10'b0111110100: data <= 20'hffdf5; 
        10'b0111110101: data <= 20'hffe65; 
        10'b0111110110: data <= 20'hfff23; 
        10'b0111110111: data <= 20'hfff39; 
        10'b0111111000: data <= 20'hfff36; 
        10'b0111111001: data <= 20'hfffbf; 
        10'b0111111010: data <= 20'h001f2; 
        10'b0111111011: data <= 20'h0009a; 
        10'b0111111100: data <= 20'hffc86; 
        10'b0111111101: data <= 20'hff7bc; 
        10'b0111111110: data <= 20'hff258; 
        10'b0111111111: data <= 20'hfeefe; 
        10'b1000000000: data <= 20'hff036; 
        10'b1000000001: data <= 20'hff138; 
        10'b1000000010: data <= 20'hfed03; 
        10'b1000000011: data <= 20'hff978; 
        10'b1000000100: data <= 20'hffe07; 
        10'b1000000101: data <= 20'h0003b; 
        10'b1000000110: data <= 20'h00557; 
        10'b1000000111: data <= 20'hffa5c; 
        10'b1000001000: data <= 20'hff913; 
        10'b1000001001: data <= 20'hffc2c; 
        10'b1000001010: data <= 20'hff748; 
        10'b1000001011: data <= 20'hffaa6; 
        10'b1000001100: data <= 20'hff705; 
        10'b1000001101: data <= 20'hff233; 
        10'b1000001110: data <= 20'hff5e8; 
        10'b1000001111: data <= 20'hff9a0; 
        10'b1000010000: data <= 20'hffafd; 
        10'b1000010001: data <= 20'h00085; 
        10'b1000010010: data <= 20'hfff73; 
        10'b1000010011: data <= 20'h0001e; 
        10'b1000010100: data <= 20'h002b4; 
        10'b1000010101: data <= 20'h002e6; 
        10'b1000010110: data <= 20'h002a7; 
        10'b1000010111: data <= 20'h00153; 
        10'b1000011000: data <= 20'hffda7; 
        10'b1000011001: data <= 20'hff540; 
        10'b1000011010: data <= 20'hfeecb; 
        10'b1000011011: data <= 20'hfed8a; 
        10'b1000011100: data <= 20'hfed0b; 
        10'b1000011101: data <= 20'hfeced; 
        10'b1000011110: data <= 20'hff315; 
        10'b1000011111: data <= 20'hff6b4; 
        10'b1000100000: data <= 20'hffa70; 
        10'b1000100001: data <= 20'h00269; 
        10'b1000100010: data <= 20'h0078e; 
        10'b1000100011: data <= 20'hff81d; 
        10'b1000100100: data <= 20'hff84e; 
        10'b1000100101: data <= 20'hff648; 
        10'b1000100110: data <= 20'hff08e; 
        10'b1000100111: data <= 20'hff15e; 
        10'b1000101000: data <= 20'hfedfa; 
        10'b1000101001: data <= 20'hfef5c; 
        10'b1000101010: data <= 20'hff355; 
        10'b1000101011: data <= 20'hff746; 
        10'b1000101100: data <= 20'hffb93; 
        10'b1000101101: data <= 20'hffe5c; 
        10'b1000101110: data <= 20'h002c6; 
        10'b1000101111: data <= 20'hffebe; 
        10'b1000110000: data <= 20'hffe8f; 
        10'b1000110001: data <= 20'hfff59; 
        10'b1000110010: data <= 20'h00124; 
        10'b1000110011: data <= 20'hfff89; 
        10'b1000110100: data <= 20'hffd48; 
        10'b1000110101: data <= 20'hff7b4; 
        10'b1000110110: data <= 20'hfeeaa; 
        10'b1000110111: data <= 20'hfedeb; 
        10'b1000111000: data <= 20'hfeef1; 
        10'b1000111001: data <= 20'hfef57; 
        10'b1000111010: data <= 20'hff462; 
        10'b1000111011: data <= 20'hff404; 
        10'b1000111100: data <= 20'h000de; 
        10'b1000111101: data <= 20'h00131; 
        10'b1000111110: data <= 20'h00402; 
        10'b1000111111: data <= 20'hff56e; 
        10'b1001000000: data <= 20'hff2ca; 
        10'b1001000001: data <= 20'hfeebd; 
        10'b1001000010: data <= 20'hfe82d; 
        10'b1001000011: data <= 20'hff0d6; 
        10'b1001000100: data <= 20'hfeb1e; 
        10'b1001000101: data <= 20'hff013; 
        10'b1001000110: data <= 20'hff47b; 
        10'b1001000111: data <= 20'hffb1a; 
        10'b1001001000: data <= 20'hffcbb; 
        10'b1001001001: data <= 20'h00279; 
        10'b1001001010: data <= 20'h00259; 
        10'b1001001011: data <= 20'h00198; 
        10'b1001001100: data <= 20'h0023a; 
        10'b1001001101: data <= 20'h00255; 
        10'b1001001110: data <= 20'h00086; 
        10'b1001001111: data <= 20'hffcf3; 
        10'b1001010000: data <= 20'hffe74; 
        10'b1001010001: data <= 20'hff89c; 
        10'b1001010010: data <= 20'hff756; 
        10'b1001010011: data <= 20'hff383; 
        10'b1001010100: data <= 20'hff4bf; 
        10'b1001010101: data <= 20'hff94f; 
        10'b1001010110: data <= 20'hff67a; 
        10'b1001010111: data <= 20'hff83d; 
        10'b1001011000: data <= 20'hffc87; 
        10'b1001011001: data <= 20'h00079; 
        10'b1001011010: data <= 20'hffdea; 
        10'b1001011011: data <= 20'hff8e0; 
        10'b1001011100: data <= 20'hff7cd; 
        10'b1001011101: data <= 20'hfeef9; 
        10'b1001011110: data <= 20'hfef0a; 
        10'b1001011111: data <= 20'hfef02; 
        10'b1001100000: data <= 20'hfee1a; 
        10'b1001100001: data <= 20'hff0d9; 
        10'b1001100010: data <= 20'hff719; 
        10'b1001100011: data <= 20'hff944; 
        10'b1001100100: data <= 20'hfffb4; 
        10'b1001100101: data <= 20'h0010a; 
        10'b1001100110: data <= 20'h0023f; 
        10'b1001100111: data <= 20'hfff84; 
        10'b1001101000: data <= 20'h000c2; 
        10'b1001101001: data <= 20'h0002d; 
        10'b1001101010: data <= 20'h00098; 
        10'b1001101011: data <= 20'hffe1f; 
        10'b1001101100: data <= 20'hfff26; 
        10'b1001101101: data <= 20'h0011a; 
        10'b1001101110: data <= 20'hffd4a; 
        10'b1001101111: data <= 20'h00158; 
        10'b1001110000: data <= 20'h00224; 
        10'b1001110001: data <= 20'hffc94; 
        10'b1001110010: data <= 20'hff97d; 
        10'b1001110011: data <= 20'hff4e3; 
        10'b1001110100: data <= 20'hff59d; 
        10'b1001110101: data <= 20'hffbcf; 
        10'b1001110110: data <= 20'h0013e; 
        10'b1001110111: data <= 20'h0013a; 
        10'b1001111000: data <= 20'hff98a; 
        10'b1001111001: data <= 20'hff800; 
        10'b1001111010: data <= 20'hff25f; 
        10'b1001111011: data <= 20'hff261; 
        10'b1001111100: data <= 20'hff0a5; 
        10'b1001111101: data <= 20'hff28f; 
        10'b1001111110: data <= 20'hff92d; 
        10'b1001111111: data <= 20'hffdb1; 
        10'b1010000000: data <= 20'h0017c; 
        10'b1010000001: data <= 20'hffe8c; 
        10'b1010000010: data <= 20'h000b6; 
        10'b1010000011: data <= 20'h0000c; 
        10'b1010000100: data <= 20'h0010d; 
        10'b1010000101: data <= 20'h0021f; 
        10'b1010000110: data <= 20'hffe5d; 
        10'b1010000111: data <= 20'hffe82; 
        10'b1010001000: data <= 20'h002d1; 
        10'b1010001001: data <= 20'h003c5; 
        10'b1010001010: data <= 20'h00832; 
        10'b1010001011: data <= 20'h00aef; 
        10'b1010001100: data <= 20'h00539; 
        10'b1010001101: data <= 20'h0010a; 
        10'b1010001110: data <= 20'hffcc9; 
        10'b1010001111: data <= 20'hff891; 
        10'b1010010000: data <= 20'hff9ec; 
        10'b1010010001: data <= 20'h0006c; 
        10'b1010010010: data <= 20'h00442; 
        10'b1010010011: data <= 20'h003ed; 
        10'b1010010100: data <= 20'hffe5d; 
        10'b1010010101: data <= 20'hffd93; 
        10'b1010010110: data <= 20'hff748; 
        10'b1010010111: data <= 20'hff3d5; 
        10'b1010011000: data <= 20'hff38d; 
        10'b1010011001: data <= 20'hff648; 
        10'b1010011010: data <= 20'hff7fc; 
        10'b1010011011: data <= 20'hffac6; 
        10'b1010011100: data <= 20'hffdb1; 
        10'b1010011101: data <= 20'h0002c; 
        10'b1010011110: data <= 20'h00027; 
        10'b1010011111: data <= 20'hfff24; 
        10'b1010100000: data <= 20'hffffb; 
        10'b1010100001: data <= 20'hfffb7; 
        10'b1010100010: data <= 20'h000c8; 
        10'b1010100011: data <= 20'h001d3; 
        10'b1010100100: data <= 20'h003e9; 
        10'b1010100101: data <= 20'h008ff; 
        10'b1010100110: data <= 20'h00d9e; 
        10'b1010100111: data <= 20'h00f58; 
        10'b1010101000: data <= 20'h00d08; 
        10'b1010101001: data <= 20'h006b8; 
        10'b1010101010: data <= 20'h00e7b; 
        10'b1010101011: data <= 20'h0088d; 
        10'b1010101100: data <= 20'h0076b; 
        10'b1010101101: data <= 20'h00a72; 
        10'b1010101110: data <= 20'h0066e; 
        10'b1010101111: data <= 20'h00947; 
        10'b1010110000: data <= 20'h0057f; 
        10'b1010110001: data <= 20'h0044a; 
        10'b1010110010: data <= 20'hfffba; 
        10'b1010110011: data <= 20'hffc00; 
        10'b1010110100: data <= 20'hffbc0; 
        10'b1010110101: data <= 20'hffad7; 
        10'b1010110110: data <= 20'hffa2c; 
        10'b1010110111: data <= 20'hffab2; 
        10'b1010111000: data <= 20'h000cf; 
        10'b1010111001: data <= 20'hfff95; 
        10'b1010111010: data <= 20'hffe9d; 
        10'b1010111011: data <= 20'h00197; 
        10'b1010111100: data <= 20'hffe95; 
        10'b1010111101: data <= 20'h0014c; 
        10'b1010111110: data <= 20'h00259; 
        10'b1010111111: data <= 20'h00233; 
        10'b1011000000: data <= 20'h00146; 
        10'b1011000001: data <= 20'h0047c; 
        10'b1011000010: data <= 20'h006a4; 
        10'b1011000011: data <= 20'h00a43; 
        10'b1011000100: data <= 20'h00fdd; 
        10'b1011000101: data <= 20'h00f7c; 
        10'b1011000110: data <= 20'h01255; 
        10'b1011000111: data <= 20'h0110f; 
        10'b1011001000: data <= 20'h00f34; 
        10'b1011001001: data <= 20'h00c0a; 
        10'b1011001010: data <= 20'h00c4c; 
        10'b1011001011: data <= 20'h00d08; 
        10'b1011001100: data <= 20'h00aec; 
        10'b1011001101: data <= 20'h00a35; 
        10'b1011001110: data <= 20'h0083a; 
        10'b1011001111: data <= 20'h002d3; 
        10'b1011010000: data <= 20'hffc89; 
        10'b1011010001: data <= 20'h00078; 
        10'b1011010010: data <= 20'hffe49; 
        10'b1011010011: data <= 20'hffebe; 
        10'b1011010100: data <= 20'hfff99; 
        10'b1011010101: data <= 20'h000c9; 
        10'b1011010110: data <= 20'h0031c; 
        10'b1011010111: data <= 20'h00204; 
        10'b1011011000: data <= 20'hffee6; 
        10'b1011011001: data <= 20'h00099; 
        10'b1011011010: data <= 20'h002f0; 
        10'b1011011011: data <= 20'hfff80; 
        10'b1011011100: data <= 20'hfff01; 
        10'b1011011101: data <= 20'h002bf; 
        10'b1011011110: data <= 20'h00033; 
        10'b1011011111: data <= 20'h00282; 
        10'b1011100000: data <= 20'h00264; 
        10'b1011100001: data <= 20'h00056; 
        10'b1011100010: data <= 20'h00373; 
        10'b1011100011: data <= 20'h00516; 
        10'b1011100100: data <= 20'h00177; 
        10'b1011100101: data <= 20'h0045d; 
        10'b1011100110: data <= 20'h0095c; 
        10'b1011100111: data <= 20'h00b8e; 
        10'b1011101000: data <= 20'h0091e; 
        10'b1011101001: data <= 20'h00bae; 
        10'b1011101010: data <= 20'h006a8; 
        10'b1011101011: data <= 20'h00325; 
        10'b1011101100: data <= 20'h0001b; 
        10'b1011101101: data <= 20'h00135; 
        10'b1011101110: data <= 20'hfffad; 
        10'b1011101111: data <= 20'h000ad; 
        10'b1011110000: data <= 20'h00023; 
        10'b1011110001: data <= 20'hfff37; 
        10'b1011110010: data <= 20'hfffd1; 
        10'b1011110011: data <= 20'hfff9c; 
        10'b1011110100: data <= 20'hffe8d; 
        10'b1011110101: data <= 20'h0012f; 
        10'b1011110110: data <= 20'h000ce; 
        10'b1011110111: data <= 20'h0017a; 
        10'b1011111000: data <= 20'h00201; 
        10'b1011111001: data <= 20'h00132; 
        10'b1011111010: data <= 20'h00085; 
        10'b1011111011: data <= 20'h00037; 
        10'b1011111100: data <= 20'h00349; 
        10'b1011111101: data <= 20'h00204; 
        10'b1011111110: data <= 20'h00098; 
        10'b1011111111: data <= 20'h00209; 
        10'b1100000000: data <= 20'h000fc; 
        10'b1100000001: data <= 20'h003cc; 
        10'b1100000010: data <= 20'h00244; 
        10'b1100000011: data <= 20'h001bb; 
        10'b1100000100: data <= 20'h00548; 
        10'b1100000101: data <= 20'h001ca; 
        10'b1100000110: data <= 20'h00195; 
        10'b1100000111: data <= 20'h003aa; 
        10'b1100001000: data <= 20'h0006f; 
        10'b1100001001: data <= 20'hfff62; 
        10'b1100001010: data <= 20'h002fd; 
        10'b1100001011: data <= 20'h001a3; 
        10'b1100001100: data <= 20'h000c3; 
        10'b1100001101: data <= 20'hfff74; 
        10'b1100001110: data <= 20'hffec7; 
        10'b1100001111: data <= 20'h001fd; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 15) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 21'h000060; 
        10'b0000000001: data <= 21'h000082; 
        10'b0000000010: data <= 21'h0003cb; 
        10'b0000000011: data <= 21'h000177; 
        10'b0000000100: data <= 21'h000630; 
        10'b0000000101: data <= 21'h1ffd40; 
        10'b0000000110: data <= 21'h1ffe2a; 
        10'b0000000111: data <= 21'h000202; 
        10'b0000001000: data <= 21'h0004c2; 
        10'b0000001001: data <= 21'h0004a9; 
        10'b0000001010: data <= 21'h1ffd5e; 
        10'b0000001011: data <= 21'h00013e; 
        10'b0000001100: data <= 21'h000158; 
        10'b0000001101: data <= 21'h1fff4c; 
        10'b0000001110: data <= 21'h0004fb; 
        10'b0000001111: data <= 21'h000155; 
        10'b0000010000: data <= 21'h000019; 
        10'b0000010001: data <= 21'h1fffd3; 
        10'b0000010010: data <= 21'h000087; 
        10'b0000010011: data <= 21'h0001b9; 
        10'b0000010100: data <= 21'h000333; 
        10'b0000010101: data <= 21'h00060f; 
        10'b0000010110: data <= 21'h1ffe60; 
        10'b0000010111: data <= 21'h000475; 
        10'b0000011000: data <= 21'h1fff62; 
        10'b0000011001: data <= 21'h000332; 
        10'b0000011010: data <= 21'h1fffbd; 
        10'b0000011011: data <= 21'h1ffffb; 
        10'b0000011100: data <= 21'h0005b4; 
        10'b0000011101: data <= 21'h1ffec8; 
        10'b0000011110: data <= 21'h000148; 
        10'b0000011111: data <= 21'h0005a0; 
        10'b0000100000: data <= 21'h000229; 
        10'b0000100001: data <= 21'h000035; 
        10'b0000100010: data <= 21'h000595; 
        10'b0000100011: data <= 21'h0001c2; 
        10'b0000100100: data <= 21'h000089; 
        10'b0000100101: data <= 21'h1fff0d; 
        10'b0000100110: data <= 21'h1fff41; 
        10'b0000100111: data <= 21'h1ffd11; 
        10'b0000101000: data <= 21'h0004ce; 
        10'b0000101001: data <= 21'h1fffa7; 
        10'b0000101010: data <= 21'h0005c3; 
        10'b0000101011: data <= 21'h1ffe7f; 
        10'b0000101100: data <= 21'h00027f; 
        10'b0000101101: data <= 21'h000455; 
        10'b0000101110: data <= 21'h0004e0; 
        10'b0000101111: data <= 21'h0003e3; 
        10'b0000110000: data <= 21'h000021; 
        10'b0000110001: data <= 21'h0003d5; 
        10'b0000110010: data <= 21'h1fffe3; 
        10'b0000110011: data <= 21'h000613; 
        10'b0000110100: data <= 21'h0004af; 
        10'b0000110101: data <= 21'h1ffe50; 
        10'b0000110110: data <= 21'h1ffe59; 
        10'b0000110111: data <= 21'h00027b; 
        10'b0000111000: data <= 21'h000567; 
        10'b0000111001: data <= 21'h000553; 
        10'b0000111010: data <= 21'h000430; 
        10'b0000111011: data <= 21'h1fff39; 
        10'b0000111100: data <= 21'h0004db; 
        10'b0000111101: data <= 21'h1ffdb0; 
        10'b0000111110: data <= 21'h1ffe1b; 
        10'b0000111111: data <= 21'h0003cd; 
        10'b0001000000: data <= 21'h000334; 
        10'b0001000001: data <= 21'h1ffe1f; 
        10'b0001000010: data <= 21'h1fff95; 
        10'b0001000011: data <= 21'h00025d; 
        10'b0001000100: data <= 21'h1fff58; 
        10'b0001000101: data <= 21'h1ffec2; 
        10'b0001000110: data <= 21'h00017c; 
        10'b0001000111: data <= 21'h0004e4; 
        10'b0001001000: data <= 21'h0003f2; 
        10'b0001001001: data <= 21'h0000bb; 
        10'b0001001010: data <= 21'h0001ef; 
        10'b0001001011: data <= 21'h000586; 
        10'b0001001100: data <= 21'h0004b0; 
        10'b0001001101: data <= 21'h00056d; 
        10'b0001001110: data <= 21'h1ffd45; 
        10'b0001001111: data <= 21'h00043b; 
        10'b0001010000: data <= 21'h00019a; 
        10'b0001010001: data <= 21'h0003bd; 
        10'b0001010010: data <= 21'h000337; 
        10'b0001010011: data <= 21'h0004c3; 
        10'b0001010100: data <= 21'h1fff91; 
        10'b0001010101: data <= 21'h000052; 
        10'b0001010110: data <= 21'h0004f3; 
        10'b0001010111: data <= 21'h1fff3f; 
        10'b0001011000: data <= 21'h00008e; 
        10'b0001011001: data <= 21'h1fffaa; 
        10'b0001011010: data <= 21'h1ffe2d; 
        10'b0001011011: data <= 21'h000338; 
        10'b0001011100: data <= 21'h000006; 
        10'b0001011101: data <= 21'h000338; 
        10'b0001011110: data <= 21'h1ffd5b; 
        10'b0001011111: data <= 21'h0000a8; 
        10'b0001100000: data <= 21'h000297; 
        10'b0001100001: data <= 21'h1ffc6e; 
        10'b0001100010: data <= 21'h0002f0; 
        10'b0001100011: data <= 21'h1ffd94; 
        10'b0001100100: data <= 21'h1ffac1; 
        10'b0001100101: data <= 21'h1ffbb5; 
        10'b0001100110: data <= 21'h1ffc51; 
        10'b0001100111: data <= 21'h1ffd85; 
        10'b0001101000: data <= 21'h1fff62; 
        10'b0001101001: data <= 21'h1ffdba; 
        10'b0001101010: data <= 21'h0001fd; 
        10'b0001101011: data <= 21'h1fffbf; 
        10'b0001101100: data <= 21'h000267; 
        10'b0001101101: data <= 21'h000619; 
        10'b0001101110: data <= 21'h1ffdff; 
        10'b0001101111: data <= 21'h000285; 
        10'b0001110000: data <= 21'h0005e9; 
        10'b0001110001: data <= 21'h1ffdd9; 
        10'b0001110010: data <= 21'h00034c; 
        10'b0001110011: data <= 21'h1ffd7d; 
        10'b0001110100: data <= 21'h000161; 
        10'b0001110101: data <= 21'h1ffedd; 
        10'b0001110110: data <= 21'h000043; 
        10'b0001110111: data <= 21'h1ffd93; 
        10'b0001111000: data <= 21'h0001d7; 
        10'b0001111001: data <= 21'h1fff23; 
        10'b0001111010: data <= 21'h1ffa36; 
        10'b0001111011: data <= 21'h1ff4d7; 
        10'b0001111100: data <= 21'h1ff447; 
        10'b0001111101: data <= 21'h1ff4d0; 
        10'b0001111110: data <= 21'h1ff2aa; 
        10'b0001111111: data <= 21'h1fea0a; 
        10'b0010000000: data <= 21'h1ff30a; 
        10'b0010000001: data <= 21'h1ff63d; 
        10'b0010000010: data <= 21'h1ff784; 
        10'b0010000011: data <= 21'h1ffdb5; 
        10'b0010000100: data <= 21'h1ff9ab; 
        10'b0010000101: data <= 21'h0002f4; 
        10'b0010000110: data <= 21'h000073; 
        10'b0010000111: data <= 21'h1ffced; 
        10'b0010001000: data <= 21'h000599; 
        10'b0010001001: data <= 21'h1fffcd; 
        10'b0010001010: data <= 21'h00057d; 
        10'b0010001011: data <= 21'h000552; 
        10'b0010001100: data <= 21'h00050a; 
        10'b0010001101: data <= 21'h000033; 
        10'b0010001110: data <= 21'h0004dc; 
        10'b0010001111: data <= 21'h1ffead; 
        10'b0010010000: data <= 21'h1ffc33; 
        10'b0010010001: data <= 21'h1fff59; 
        10'b0010010010: data <= 21'h1ffd16; 
        10'b0010010011: data <= 21'h1ffeef; 
        10'b0010010100: data <= 21'h1ffc8d; 
        10'b0010010101: data <= 21'h1ff7fd; 
        10'b0010010110: data <= 21'h1fec53; 
        10'b0010010111: data <= 21'h1fe7da; 
        10'b0010011000: data <= 21'h1fe19b; 
        10'b0010011001: data <= 21'h1fdc64; 
        10'b0010011010: data <= 21'h1fd392; 
        10'b0010011011: data <= 21'h1fd3e7; 
        10'b0010011100: data <= 21'h1fd1c2; 
        10'b0010011101: data <= 21'h1fd734; 
        10'b0010011110: data <= 21'h1fdd6e; 
        10'b0010011111: data <= 21'h1fe5b2; 
        10'b0010100000: data <= 21'h1fed50; 
        10'b0010100001: data <= 21'h1ff955; 
        10'b0010100010: data <= 21'h1ff5b1; 
        10'b0010100011: data <= 21'h1ffeb6; 
        10'b0010100100: data <= 21'h000483; 
        10'b0010100101: data <= 21'h000399; 
        10'b0010100110: data <= 21'h1fff14; 
        10'b0010100111: data <= 21'h000034; 
        10'b0010101000: data <= 21'h000430; 
        10'b0010101001: data <= 21'h0005bc; 
        10'b0010101010: data <= 21'h000067; 
        10'b0010101011: data <= 21'h0000ee; 
        10'b0010101100: data <= 21'h000635; 
        10'b0010101101: data <= 21'h000764; 
        10'b0010101110: data <= 21'h0008a6; 
        10'b0010101111: data <= 21'h000d06; 
        10'b0010110000: data <= 21'h001351; 
        10'b0010110001: data <= 21'h000f79; 
        10'b0010110010: data <= 21'h001077; 
        10'b0010110011: data <= 21'h0002f6; 
        10'b0010110100: data <= 21'h1ff2cb; 
        10'b0010110101: data <= 21'h1fe449; 
        10'b0010110110: data <= 21'h1fe314; 
        10'b0010110111: data <= 21'h1ff0fa; 
        10'b0010111000: data <= 21'h1ff6e1; 
        10'b0010111001: data <= 21'h1ff52c; 
        10'b0010111010: data <= 21'h1ff2e0; 
        10'b0010111011: data <= 21'h1ff0d0; 
        10'b0010111100: data <= 21'h1fe902; 
        10'b0010111101: data <= 21'h1ff760; 
        10'b0010111110: data <= 21'h1fefe2; 
        10'b0010111111: data <= 21'h1ff445; 
        10'b0011000000: data <= 21'h1ff826; 
        10'b0011000001: data <= 21'h1ffd5e; 
        10'b0011000010: data <= 21'h1ffd47; 
        10'b0011000011: data <= 21'h0000a2; 
        10'b0011000100: data <= 21'h0003d1; 
        10'b0011000101: data <= 21'h0005c8; 
        10'b0011000110: data <= 21'h0004c2; 
        10'b0011000111: data <= 21'h000b41; 
        10'b0011001000: data <= 21'h000da5; 
        10'b0011001001: data <= 21'h000c45; 
        10'b0011001010: data <= 21'h0011c5; 
        10'b0011001011: data <= 21'h001b2a; 
        10'b0011001100: data <= 21'h002535; 
        10'b0011001101: data <= 21'h001d7a; 
        10'b0011001110: data <= 21'h001456; 
        10'b0011001111: data <= 21'h001667; 
        10'b0011010000: data <= 21'h0017dd; 
        10'b0011010001: data <= 21'h000496; 
        10'b0011010010: data <= 21'h000363; 
        10'b0011010011: data <= 21'h00088b; 
        10'b0011010100: data <= 21'h00192f; 
        10'b0011010101: data <= 21'h001bff; 
        10'b0011010110: data <= 21'h0012f9; 
        10'b0011010111: data <= 21'h000f36; 
        10'b0011011000: data <= 21'h0003b6; 
        10'b0011011001: data <= 21'h1ffbca; 
        10'b0011011010: data <= 21'h0001fa; 
        10'b0011011011: data <= 21'h1ffb76; 
        10'b0011011100: data <= 21'h1ffbc2; 
        10'b0011011101: data <= 21'h1fffc6; 
        10'b0011011110: data <= 21'h000300; 
        10'b0011011111: data <= 21'h1ffedf; 
        10'b0011100000: data <= 21'h1ffd14; 
        10'b0011100001: data <= 21'h000610; 
        10'b0011100010: data <= 21'h000257; 
        10'b0011100011: data <= 21'h000981; 
        10'b0011100100: data <= 21'h00133e; 
        10'b0011100101: data <= 21'h00115b; 
        10'b0011100110: data <= 21'h00173d; 
        10'b0011100111: data <= 21'h0029b7; 
        10'b0011101000: data <= 21'h001c14; 
        10'b0011101001: data <= 21'h001358; 
        10'b0011101010: data <= 21'h00189c; 
        10'b0011101011: data <= 21'h0020f6; 
        10'b0011101100: data <= 21'h001f54; 
        10'b0011101101: data <= 21'h000fc3; 
        10'b0011101110: data <= 21'h000936; 
        10'b0011101111: data <= 21'h000cc9; 
        10'b0011110000: data <= 21'h001637; 
        10'b0011110001: data <= 21'h002226; 
        10'b0011110010: data <= 21'h001767; 
        10'b0011110011: data <= 21'h00140c; 
        10'b0011110100: data <= 21'h001000; 
        10'b0011110101: data <= 21'h000060; 
        10'b0011110110: data <= 21'h0009b3; 
        10'b0011110111: data <= 21'h00083b; 
        10'b0011111000: data <= 21'h1ffa21; 
        10'b0011111001: data <= 21'h1ffd32; 
        10'b0011111010: data <= 21'h00033f; 
        10'b0011111011: data <= 21'h0004fe; 
        10'b0011111100: data <= 21'h000293; 
        10'b0011111101: data <= 21'h0004d3; 
        10'b0011111110: data <= 21'h00067b; 
        10'b0011111111: data <= 21'h000db4; 
        10'b0100000000: data <= 21'h0012dc; 
        10'b0100000001: data <= 21'h00156b; 
        10'b0100000010: data <= 21'h0007db; 
        10'b0100000011: data <= 21'h000a73; 
        10'b0100000100: data <= 21'h000bd9; 
        10'b0100000101: data <= 21'h0007d5; 
        10'b0100000110: data <= 21'h001333; 
        10'b0100000111: data <= 21'h001786; 
        10'b0100001000: data <= 21'h001dfe; 
        10'b0100001001: data <= 21'h001866; 
        10'b0100001010: data <= 21'h0022f4; 
        10'b0100001011: data <= 21'h002b07; 
        10'b0100001100: data <= 21'h0027a3; 
        10'b0100001101: data <= 21'h002c3c; 
        10'b0100001110: data <= 21'h001ce1; 
        10'b0100001111: data <= 21'h001d69; 
        10'b0100010000: data <= 21'h0018bb; 
        10'b0100010001: data <= 21'h0014a1; 
        10'b0100010010: data <= 21'h0009c4; 
        10'b0100010011: data <= 21'h1ffc73; 
        10'b0100010100: data <= 21'h1ff9ff; 
        10'b0100010101: data <= 21'h1ffd0f; 
        10'b0100010110: data <= 21'h00029c; 
        10'b0100010111: data <= 21'h1ffeaa; 
        10'b0100011000: data <= 21'h0000ff; 
        10'b0100011001: data <= 21'h000543; 
        10'b0100011010: data <= 21'h0005d6; 
        10'b0100011011: data <= 21'h001109; 
        10'b0100011100: data <= 21'h001384; 
        10'b0100011101: data <= 21'h00103a; 
        10'b0100011110: data <= 21'h0002fe; 
        10'b0100011111: data <= 21'h0004e1; 
        10'b0100100000: data <= 21'h1ff970; 
        10'b0100100001: data <= 21'h1fffc0; 
        10'b0100100010: data <= 21'h000be8; 
        10'b0100100011: data <= 21'h0014f7; 
        10'b0100100100: data <= 21'h000e96; 
        10'b0100100101: data <= 21'h0021f2; 
        10'b0100100110: data <= 21'h002bad; 
        10'b0100100111: data <= 21'h0035a4; 
        10'b0100101000: data <= 21'h003d14; 
        10'b0100101001: data <= 21'h002d44; 
        10'b0100101010: data <= 21'h0023a6; 
        10'b0100101011: data <= 21'h002515; 
        10'b0100101100: data <= 21'h00208e; 
        10'b0100101101: data <= 21'h001bae; 
        10'b0100101110: data <= 21'h000c3d; 
        10'b0100101111: data <= 21'h1ffb02; 
        10'b0100110000: data <= 21'h1ff7bd; 
        10'b0100110001: data <= 21'h1ffca6; 
        10'b0100110010: data <= 21'h0000a1; 
        10'b0100110011: data <= 21'h1ffebf; 
        10'b0100110100: data <= 21'h0004a1; 
        10'b0100110101: data <= 21'h000340; 
        10'b0100110110: data <= 21'h0005e7; 
        10'b0100110111: data <= 21'h001173; 
        10'b0100111000: data <= 21'h001507; 
        10'b0100111001: data <= 21'h000a6d; 
        10'b0100111010: data <= 21'h0003ca; 
        10'b0100111011: data <= 21'h000366; 
        10'b0100111100: data <= 21'h0000f9; 
        10'b0100111101: data <= 21'h000ca0; 
        10'b0100111110: data <= 21'h000683; 
        10'b0100111111: data <= 21'h000837; 
        10'b0101000000: data <= 21'h000d92; 
        10'b0101000001: data <= 21'h000d73; 
        10'b0101000010: data <= 21'h000dfc; 
        10'b0101000011: data <= 21'h00290d; 
        10'b0101000100: data <= 21'h00354f; 
        10'b0101000101: data <= 21'h002387; 
        10'b0101000110: data <= 21'h0023e1; 
        10'b0101000111: data <= 21'h001b96; 
        10'b0101001000: data <= 21'h001acd; 
        10'b0101001001: data <= 21'h0010dc; 
        10'b0101001010: data <= 21'h000c2c; 
        10'b0101001011: data <= 21'h1ffbc5; 
        10'b0101001100: data <= 21'h1ff3b0; 
        10'b0101001101: data <= 21'h1fffa8; 
        10'b0101001110: data <= 21'h00012d; 
        10'b0101001111: data <= 21'h000565; 
        10'b0101010000: data <= 21'h000420; 
        10'b0101010001: data <= 21'h1fffb4; 
        10'b0101010010: data <= 21'h0002f0; 
        10'b0101010011: data <= 21'h000afe; 
        10'b0101010100: data <= 21'h000c57; 
        10'b0101010101: data <= 21'h000208; 
        10'b0101010110: data <= 21'h0002c2; 
        10'b0101010111: data <= 21'h000bbe; 
        10'b0101011000: data <= 21'h00080d; 
        10'b0101011001: data <= 21'h1fff88; 
        10'b0101011010: data <= 21'h1ff666; 
        10'b0101011011: data <= 21'h1fe671; 
        10'b0101011100: data <= 21'h1fc9f8; 
        10'b0101011101: data <= 21'h1fac5e; 
        10'b0101011110: data <= 21'h1fc167; 
        10'b0101011111: data <= 21'h00015c; 
        10'b0101100000: data <= 21'h00235b; 
        10'b0101100001: data <= 21'h002017; 
        10'b0101100010: data <= 21'h000ca0; 
        10'b0101100011: data <= 21'h000489; 
        10'b0101100100: data <= 21'h0000d9; 
        10'b0101100101: data <= 21'h1ffb60; 
        10'b0101100110: data <= 21'h1ffbce; 
        10'b0101100111: data <= 21'h1ff870; 
        10'b0101101000: data <= 21'h1ffa8d; 
        10'b0101101001: data <= 21'h00051a; 
        10'b0101101010: data <= 21'h000395; 
        10'b0101101011: data <= 21'h00000b; 
        10'b0101101100: data <= 21'h000478; 
        10'b0101101101: data <= 21'h0002a1; 
        10'b0101101110: data <= 21'h0004d1; 
        10'b0101101111: data <= 21'h0009f9; 
        10'b0101110000: data <= 21'h0003b7; 
        10'b0101110001: data <= 21'h000198; 
        10'b0101110010: data <= 21'h1ffcba; 
        10'b0101110011: data <= 21'h000226; 
        10'b0101110100: data <= 21'h1ffe7e; 
        10'b0101110101: data <= 21'h1ff7cf; 
        10'b0101110110: data <= 21'h1fe52e; 
        10'b0101110111: data <= 21'h1fc775; 
        10'b0101111000: data <= 21'h1f9cbb; 
        10'b0101111001: data <= 21'h1f911e; 
        10'b0101111010: data <= 21'h1fc4ab; 
        10'b0101111011: data <= 21'h1ff838; 
        10'b0101111100: data <= 21'h00120c; 
        10'b0101111101: data <= 21'h000ba4; 
        10'b0101111110: data <= 21'h000285; 
        10'b0101111111: data <= 21'h00054b; 
        10'b0110000000: data <= 21'h1ff521; 
        10'b0110000001: data <= 21'h1ff217; 
        10'b0110000010: data <= 21'h1ffcbc; 
        10'b0110000011: data <= 21'h000107; 
        10'b0110000100: data <= 21'h1ffd5c; 
        10'b0110000101: data <= 21'h1ffde3; 
        10'b0110000110: data <= 21'h0002d3; 
        10'b0110000111: data <= 21'h1ffd42; 
        10'b0110001000: data <= 21'h1ffecd; 
        10'b0110001001: data <= 21'h000262; 
        10'b0110001010: data <= 21'h0008ed; 
        10'b0110001011: data <= 21'h000b1e; 
        10'b0110001100: data <= 21'h00070c; 
        10'b0110001101: data <= 21'h00082f; 
        10'b0110001110: data <= 21'h1ffd4a; 
        10'b0110001111: data <= 21'h1ffa4c; 
        10'b0110010000: data <= 21'h1ff36b; 
        10'b0110010001: data <= 21'h1fe286; 
        10'b0110010010: data <= 21'h1fd4ac; 
        10'b0110010011: data <= 21'h1fbcf9; 
        10'b0110010100: data <= 21'h1faa15; 
        10'b0110010101: data <= 21'h1fb787; 
        10'b0110010110: data <= 21'h1fe56e; 
        10'b0110010111: data <= 21'h00009e; 
        10'b0110011000: data <= 21'h000586; 
        10'b0110011001: data <= 21'h000b72; 
        10'b0110011010: data <= 21'h0020d7; 
        10'b0110011011: data <= 21'h00234c; 
        10'b0110011100: data <= 21'h00153d; 
        10'b0110011101: data <= 21'h000d90; 
        10'b0110011110: data <= 21'h000da5; 
        10'b0110011111: data <= 21'h000bd5; 
        10'b0110100000: data <= 21'h000400; 
        10'b0110100001: data <= 21'h000130; 
        10'b0110100010: data <= 21'h1ffe1c; 
        10'b0110100011: data <= 21'h1ffe49; 
        10'b0110100100: data <= 21'h0002e1; 
        10'b0110100101: data <= 21'h00043f; 
        10'b0110100110: data <= 21'h00018f; 
        10'b0110100111: data <= 21'h000436; 
        10'b0110101000: data <= 21'h000433; 
        10'b0110101001: data <= 21'h1ff41b; 
        10'b0110101010: data <= 21'h1ffab3; 
        10'b0110101011: data <= 21'h1ff8a1; 
        10'b0110101100: data <= 21'h1fe05d; 
        10'b0110101101: data <= 21'h1fd99d; 
        10'b0110101110: data <= 21'h1fccf8; 
        10'b0110101111: data <= 21'h1fc586; 
        10'b0110110000: data <= 21'h1fc04e; 
        10'b0110110001: data <= 21'h1fd10f; 
        10'b0110110010: data <= 21'h1fe495; 
        10'b0110110011: data <= 21'h0000d6; 
        10'b0110110100: data <= 21'h0002fe; 
        10'b0110110101: data <= 21'h002caa; 
        10'b0110110110: data <= 21'h00344b; 
        10'b0110110111: data <= 21'h002b18; 
        10'b0110111000: data <= 21'h002645; 
        10'b0110111001: data <= 21'h0020ec; 
        10'b0110111010: data <= 21'h001547; 
        10'b0110111011: data <= 21'h00099c; 
        10'b0110111100: data <= 21'h1fff9a; 
        10'b0110111101: data <= 21'h1ffd58; 
        10'b0110111110: data <= 21'h0000b6; 
        10'b0110111111: data <= 21'h000494; 
        10'b0111000000: data <= 21'h0002da; 
        10'b0111000001: data <= 21'h0005ab; 
        10'b0111000010: data <= 21'h1fff88; 
        10'b0111000011: data <= 21'h0005f3; 
        10'b0111000100: data <= 21'h0004ae; 
        10'b0111000101: data <= 21'h1ffaac; 
        10'b0111000110: data <= 21'h1ff879; 
        10'b0111000111: data <= 21'h1ffeeb; 
        10'b0111001000: data <= 21'h1fe688; 
        10'b0111001001: data <= 21'h1fe341; 
        10'b0111001010: data <= 21'h1fd1b7; 
        10'b0111001011: data <= 21'h1fc8f9; 
        10'b0111001100: data <= 21'h1fdd81; 
        10'b0111001101: data <= 21'h1fecb4; 
        10'b0111001110: data <= 21'h1fe407; 
        10'b0111001111: data <= 21'h000e64; 
        10'b0111010000: data <= 21'h001169; 
        10'b0111010001: data <= 21'h0025ca; 
        10'b0111010010: data <= 21'h002060; 
        10'b0111010011: data <= 21'h0021ec; 
        10'b0111010100: data <= 21'h001afe; 
        10'b0111010101: data <= 21'h00148e; 
        10'b0111010110: data <= 21'h00040e; 
        10'b0111010111: data <= 21'h1ff78b; 
        10'b0111011000: data <= 21'h1ffac0; 
        10'b0111011001: data <= 21'h1ffd04; 
        10'b0111011010: data <= 21'h000336; 
        10'b0111011011: data <= 21'h000597; 
        10'b0111011100: data <= 21'h00002e; 
        10'b0111011101: data <= 21'h0000b8; 
        10'b0111011110: data <= 21'h00036f; 
        10'b0111011111: data <= 21'h1fffc4; 
        10'b0111100000: data <= 21'h000121; 
        10'b0111100001: data <= 21'h1ffc9a; 
        10'b0111100010: data <= 21'h1feed6; 
        10'b0111100011: data <= 21'h1fe962; 
        10'b0111100100: data <= 21'h1fe39d; 
        10'b0111100101: data <= 21'h1fe892; 
        10'b0111100110: data <= 21'h1fe0f1; 
        10'b0111100111: data <= 21'h1fe8f4; 
        10'b0111101000: data <= 21'h1ff8a3; 
        10'b0111101001: data <= 21'h0005c0; 
        10'b0111101010: data <= 21'h000343; 
        10'b0111101011: data <= 21'h0005ba; 
        10'b0111101100: data <= 21'h1ffc9b; 
        10'b0111101101: data <= 21'h000915; 
        10'b0111101110: data <= 21'h000819; 
        10'b0111101111: data <= 21'h0005c1; 
        10'b0111110000: data <= 21'h00030d; 
        10'b0111110001: data <= 21'h1ffb4b; 
        10'b0111110010: data <= 21'h1ff58f; 
        10'b0111110011: data <= 21'h1ffb4c; 
        10'b0111110100: data <= 21'h1ffbea; 
        10'b0111110101: data <= 21'h1ffccb; 
        10'b0111110110: data <= 21'h1ffe47; 
        10'b0111110111: data <= 21'h1ffe73; 
        10'b0111111000: data <= 21'h1ffe6d; 
        10'b0111111001: data <= 21'h1fff7d; 
        10'b0111111010: data <= 21'h0003e3; 
        10'b0111111011: data <= 21'h000133; 
        10'b0111111100: data <= 21'h1ff90d; 
        10'b0111111101: data <= 21'h1fef77; 
        10'b0111111110: data <= 21'h1fe4af; 
        10'b0111111111: data <= 21'h1fddfc; 
        10'b1000000000: data <= 21'h1fe06d; 
        10'b1000000001: data <= 21'h1fe271; 
        10'b1000000010: data <= 21'h1fda07; 
        10'b1000000011: data <= 21'h1ff2f0; 
        10'b1000000100: data <= 21'h1ffc0e; 
        10'b1000000101: data <= 21'h000077; 
        10'b1000000110: data <= 21'h000aae; 
        10'b1000000111: data <= 21'h1ff4b9; 
        10'b1000001000: data <= 21'h1ff226; 
        10'b1000001001: data <= 21'h1ff859; 
        10'b1000001010: data <= 21'h1fee8f; 
        10'b1000001011: data <= 21'h1ff54c; 
        10'b1000001100: data <= 21'h1fee09; 
        10'b1000001101: data <= 21'h1fe467; 
        10'b1000001110: data <= 21'h1febcf; 
        10'b1000001111: data <= 21'h1ff340; 
        10'b1000010000: data <= 21'h1ff5f9; 
        10'b1000010001: data <= 21'h00010a; 
        10'b1000010010: data <= 21'h1ffee6; 
        10'b1000010011: data <= 21'h00003c; 
        10'b1000010100: data <= 21'h000569; 
        10'b1000010101: data <= 21'h0005cb; 
        10'b1000010110: data <= 21'h00054e; 
        10'b1000010111: data <= 21'h0002a5; 
        10'b1000011000: data <= 21'h1ffb4f; 
        10'b1000011001: data <= 21'h1fea81; 
        10'b1000011010: data <= 21'h1fdd96; 
        10'b1000011011: data <= 21'h1fdb14; 
        10'b1000011100: data <= 21'h1fda17; 
        10'b1000011101: data <= 21'h1fd9db; 
        10'b1000011110: data <= 21'h1fe62b; 
        10'b1000011111: data <= 21'h1fed68; 
        10'b1000100000: data <= 21'h1ff4e0; 
        10'b1000100001: data <= 21'h0004d3; 
        10'b1000100010: data <= 21'h000f1c; 
        10'b1000100011: data <= 21'h1ff039; 
        10'b1000100100: data <= 21'h1ff09c; 
        10'b1000100101: data <= 21'h1fec91; 
        10'b1000100110: data <= 21'h1fe11b; 
        10'b1000100111: data <= 21'h1fe2bc; 
        10'b1000101000: data <= 21'h1fdbf4; 
        10'b1000101001: data <= 21'h1fdeb8; 
        10'b1000101010: data <= 21'h1fe6aa; 
        10'b1000101011: data <= 21'h1fee8c; 
        10'b1000101100: data <= 21'h1ff727; 
        10'b1000101101: data <= 21'h1ffcb8; 
        10'b1000101110: data <= 21'h00058d; 
        10'b1000101111: data <= 21'h1ffd7c; 
        10'b1000110000: data <= 21'h1ffd1d; 
        10'b1000110001: data <= 21'h1ffeb1; 
        10'b1000110010: data <= 21'h000247; 
        10'b1000110011: data <= 21'h1fff12; 
        10'b1000110100: data <= 21'h1ffa90; 
        10'b1000110101: data <= 21'h1fef69; 
        10'b1000110110: data <= 21'h1fdd54; 
        10'b1000110111: data <= 21'h1fdbd5; 
        10'b1000111000: data <= 21'h1fdde2; 
        10'b1000111001: data <= 21'h1fdeae; 
        10'b1000111010: data <= 21'h1fe8c5; 
        10'b1000111011: data <= 21'h1fe808; 
        10'b1000111100: data <= 21'h0001bc; 
        10'b1000111101: data <= 21'h000261; 
        10'b1000111110: data <= 21'h000805; 
        10'b1000111111: data <= 21'h1feadb; 
        10'b1001000000: data <= 21'h1fe593; 
        10'b1001000001: data <= 21'h1fdd7b; 
        10'b1001000010: data <= 21'h1fd05a; 
        10'b1001000011: data <= 21'h1fe1ad; 
        10'b1001000100: data <= 21'h1fd63c; 
        10'b1001000101: data <= 21'h1fe026; 
        10'b1001000110: data <= 21'h1fe8f5; 
        10'b1001000111: data <= 21'h1ff634; 
        10'b1001001000: data <= 21'h1ff975; 
        10'b1001001001: data <= 21'h0004f1; 
        10'b1001001010: data <= 21'h0004b2; 
        10'b1001001011: data <= 21'h000330; 
        10'b1001001100: data <= 21'h000474; 
        10'b1001001101: data <= 21'h0004aa; 
        10'b1001001110: data <= 21'h00010c; 
        10'b1001001111: data <= 21'h1ff9e7; 
        10'b1001010000: data <= 21'h1ffce8; 
        10'b1001010001: data <= 21'h1ff138; 
        10'b1001010010: data <= 21'h1feeac; 
        10'b1001010011: data <= 21'h1fe705; 
        10'b1001010100: data <= 21'h1fe97e; 
        10'b1001010101: data <= 21'h1ff29e; 
        10'b1001010110: data <= 21'h1fecf4; 
        10'b1001010111: data <= 21'h1ff079; 
        10'b1001011000: data <= 21'h1ff90f; 
        10'b1001011001: data <= 21'h0000f1; 
        10'b1001011010: data <= 21'h1ffbd5; 
        10'b1001011011: data <= 21'h1ff1c0; 
        10'b1001011100: data <= 21'h1fef9b; 
        10'b1001011101: data <= 21'h1fddf2; 
        10'b1001011110: data <= 21'h1fde15; 
        10'b1001011111: data <= 21'h1fde03; 
        10'b1001100000: data <= 21'h1fdc34; 
        10'b1001100001: data <= 21'h1fe1b2; 
        10'b1001100010: data <= 21'h1fee32; 
        10'b1001100011: data <= 21'h1ff289; 
        10'b1001100100: data <= 21'h1fff69; 
        10'b1001100101: data <= 21'h000213; 
        10'b1001100110: data <= 21'h00047e; 
        10'b1001100111: data <= 21'h1fff08; 
        10'b1001101000: data <= 21'h000184; 
        10'b1001101001: data <= 21'h00005a; 
        10'b1001101010: data <= 21'h000131; 
        10'b1001101011: data <= 21'h1ffc3f; 
        10'b1001101100: data <= 21'h1ffe4c; 
        10'b1001101101: data <= 21'h000233; 
        10'b1001101110: data <= 21'h1ffa95; 
        10'b1001101111: data <= 21'h0002b0; 
        10'b1001110000: data <= 21'h000448; 
        10'b1001110001: data <= 21'h1ff928; 
        10'b1001110010: data <= 21'h1ff2f9; 
        10'b1001110011: data <= 21'h1fe9c6; 
        10'b1001110100: data <= 21'h1feb3a; 
        10'b1001110101: data <= 21'h1ff79f; 
        10'b1001110110: data <= 21'h00027d; 
        10'b1001110111: data <= 21'h000274; 
        10'b1001111000: data <= 21'h1ff315; 
        10'b1001111001: data <= 21'h1ff001; 
        10'b1001111010: data <= 21'h1fe4bf; 
        10'b1001111011: data <= 21'h1fe4c1; 
        10'b1001111100: data <= 21'h1fe14b; 
        10'b1001111101: data <= 21'h1fe51f; 
        10'b1001111110: data <= 21'h1ff25a; 
        10'b1001111111: data <= 21'h1ffb63; 
        10'b1010000000: data <= 21'h0002f9; 
        10'b1010000001: data <= 21'h1ffd19; 
        10'b1010000010: data <= 21'h00016c; 
        10'b1010000011: data <= 21'h000017; 
        10'b1010000100: data <= 21'h000219; 
        10'b1010000101: data <= 21'h00043f; 
        10'b1010000110: data <= 21'h1ffcb9; 
        10'b1010000111: data <= 21'h1ffd04; 
        10'b1010001000: data <= 21'h0005a2; 
        10'b1010001001: data <= 21'h000789; 
        10'b1010001010: data <= 21'h001065; 
        10'b1010001011: data <= 21'h0015dd; 
        10'b1010001100: data <= 21'h000a71; 
        10'b1010001101: data <= 21'h000214; 
        10'b1010001110: data <= 21'h1ff991; 
        10'b1010001111: data <= 21'h1ff123; 
        10'b1010010000: data <= 21'h1ff3d8; 
        10'b1010010001: data <= 21'h0000d7; 
        10'b1010010010: data <= 21'h000884; 
        10'b1010010011: data <= 21'h0007d9; 
        10'b1010010100: data <= 21'h1ffcba; 
        10'b1010010101: data <= 21'h1ffb26; 
        10'b1010010110: data <= 21'h1fee90; 
        10'b1010010111: data <= 21'h1fe7aa; 
        10'b1010011000: data <= 21'h1fe71a; 
        10'b1010011001: data <= 21'h1fec90; 
        10'b1010011010: data <= 21'h1feff7; 
        10'b1010011011: data <= 21'h1ff58c; 
        10'b1010011100: data <= 21'h1ffb62; 
        10'b1010011101: data <= 21'h000058; 
        10'b1010011110: data <= 21'h00004e; 
        10'b1010011111: data <= 21'h1ffe48; 
        10'b1010100000: data <= 21'h1ffff5; 
        10'b1010100001: data <= 21'h1fff6d; 
        10'b1010100010: data <= 21'h00018f; 
        10'b1010100011: data <= 21'h0003a7; 
        10'b1010100100: data <= 21'h0007d3; 
        10'b1010100101: data <= 21'h0011fe; 
        10'b1010100110: data <= 21'h001b3c; 
        10'b1010100111: data <= 21'h001eb0; 
        10'b1010101000: data <= 21'h001a11; 
        10'b1010101001: data <= 21'h000d71; 
        10'b1010101010: data <= 21'h001cf6; 
        10'b1010101011: data <= 21'h001119; 
        10'b1010101100: data <= 21'h000ed6; 
        10'b1010101101: data <= 21'h0014e5; 
        10'b1010101110: data <= 21'h000cdd; 
        10'b1010101111: data <= 21'h00128f; 
        10'b1010110000: data <= 21'h000afe; 
        10'b1010110001: data <= 21'h000893; 
        10'b1010110010: data <= 21'h1fff73; 
        10'b1010110011: data <= 21'h1ff800; 
        10'b1010110100: data <= 21'h1ff780; 
        10'b1010110101: data <= 21'h1ff5ae; 
        10'b1010110110: data <= 21'h1ff459; 
        10'b1010110111: data <= 21'h1ff564; 
        10'b1010111000: data <= 21'h00019f; 
        10'b1010111001: data <= 21'h1fff2a; 
        10'b1010111010: data <= 21'h1ffd3a; 
        10'b1010111011: data <= 21'h00032e; 
        10'b1010111100: data <= 21'h1ffd2a; 
        10'b1010111101: data <= 21'h000297; 
        10'b1010111110: data <= 21'h0004b2; 
        10'b1010111111: data <= 21'h000465; 
        10'b1011000000: data <= 21'h00028d; 
        10'b1011000001: data <= 21'h0008f8; 
        10'b1011000010: data <= 21'h000d47; 
        10'b1011000011: data <= 21'h001486; 
        10'b1011000100: data <= 21'h001fba; 
        10'b1011000101: data <= 21'h001ef8; 
        10'b1011000110: data <= 21'h0024a9; 
        10'b1011000111: data <= 21'h00221e; 
        10'b1011001000: data <= 21'h001e67; 
        10'b1011001001: data <= 21'h001815; 
        10'b1011001010: data <= 21'h001899; 
        10'b1011001011: data <= 21'h001a11; 
        10'b1011001100: data <= 21'h0015d8; 
        10'b1011001101: data <= 21'h00146a; 
        10'b1011001110: data <= 21'h001074; 
        10'b1011001111: data <= 21'h0005a6; 
        10'b1011010000: data <= 21'h1ff911; 
        10'b1011010001: data <= 21'h0000f0; 
        10'b1011010010: data <= 21'h1ffc93; 
        10'b1011010011: data <= 21'h1ffd7c; 
        10'b1011010100: data <= 21'h1fff33; 
        10'b1011010101: data <= 21'h000192; 
        10'b1011010110: data <= 21'h000637; 
        10'b1011010111: data <= 21'h000409; 
        10'b1011011000: data <= 21'h1ffdcc; 
        10'b1011011001: data <= 21'h000131; 
        10'b1011011010: data <= 21'h0005e0; 
        10'b1011011011: data <= 21'h1fff00; 
        10'b1011011100: data <= 21'h1ffe01; 
        10'b1011011101: data <= 21'h00057d; 
        10'b1011011110: data <= 21'h000065; 
        10'b1011011111: data <= 21'h000504; 
        10'b1011100000: data <= 21'h0004c9; 
        10'b1011100001: data <= 21'h0000ab; 
        10'b1011100010: data <= 21'h0006e6; 
        10'b1011100011: data <= 21'h000a2b; 
        10'b1011100100: data <= 21'h0002ef; 
        10'b1011100101: data <= 21'h0008ba; 
        10'b1011100110: data <= 21'h0012b8; 
        10'b1011100111: data <= 21'h00171d; 
        10'b1011101000: data <= 21'h00123b; 
        10'b1011101001: data <= 21'h00175c; 
        10'b1011101010: data <= 21'h000d50; 
        10'b1011101011: data <= 21'h00064a; 
        10'b1011101100: data <= 21'h000035; 
        10'b1011101101: data <= 21'h00026b; 
        10'b1011101110: data <= 21'h1fff5a; 
        10'b1011101111: data <= 21'h000159; 
        10'b1011110000: data <= 21'h000045; 
        10'b1011110001: data <= 21'h1ffe6e; 
        10'b1011110010: data <= 21'h1fffa1; 
        10'b1011110011: data <= 21'h1fff37; 
        10'b1011110100: data <= 21'h1ffd1a; 
        10'b1011110101: data <= 21'h00025e; 
        10'b1011110110: data <= 21'h00019c; 
        10'b1011110111: data <= 21'h0002f3; 
        10'b1011111000: data <= 21'h000402; 
        10'b1011111001: data <= 21'h000265; 
        10'b1011111010: data <= 21'h000109; 
        10'b1011111011: data <= 21'h00006e; 
        10'b1011111100: data <= 21'h000692; 
        10'b1011111101: data <= 21'h000408; 
        10'b1011111110: data <= 21'h000130; 
        10'b1011111111: data <= 21'h000412; 
        10'b1100000000: data <= 21'h0001f9; 
        10'b1100000001: data <= 21'h000799; 
        10'b1100000010: data <= 21'h000488; 
        10'b1100000011: data <= 21'h000375; 
        10'b1100000100: data <= 21'h000a8f; 
        10'b1100000101: data <= 21'h000394; 
        10'b1100000110: data <= 21'h00032b; 
        10'b1100000111: data <= 21'h000754; 
        10'b1100001000: data <= 21'h0000df; 
        10'b1100001001: data <= 21'h1ffec3; 
        10'b1100001010: data <= 21'h0005fb; 
        10'b1100001011: data <= 21'h000347; 
        10'b1100001100: data <= 21'h000185; 
        10'b1100001101: data <= 21'h1ffee8; 
        10'b1100001110: data <= 21'h1ffd8e; 
        10'b1100001111: data <= 21'h0003fb; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 16) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 22'h0000c1; 
        10'b0000000001: data <= 22'h000104; 
        10'b0000000010: data <= 22'h000797; 
        10'b0000000011: data <= 22'h0002ed; 
        10'b0000000100: data <= 22'h000c60; 
        10'b0000000101: data <= 22'h3ffa80; 
        10'b0000000110: data <= 22'h3ffc54; 
        10'b0000000111: data <= 22'h000404; 
        10'b0000001000: data <= 22'h000984; 
        10'b0000001001: data <= 22'h000953; 
        10'b0000001010: data <= 22'h3ffabc; 
        10'b0000001011: data <= 22'h00027d; 
        10'b0000001100: data <= 22'h0002b0; 
        10'b0000001101: data <= 22'h3ffe98; 
        10'b0000001110: data <= 22'h0009f6; 
        10'b0000001111: data <= 22'h0002aa; 
        10'b0000010000: data <= 22'h000033; 
        10'b0000010001: data <= 22'h3fffa6; 
        10'b0000010010: data <= 22'h00010d; 
        10'b0000010011: data <= 22'h000373; 
        10'b0000010100: data <= 22'h000667; 
        10'b0000010101: data <= 22'h000c1d; 
        10'b0000010110: data <= 22'h3ffcc1; 
        10'b0000010111: data <= 22'h0008ea; 
        10'b0000011000: data <= 22'h3ffec3; 
        10'b0000011001: data <= 22'h000664; 
        10'b0000011010: data <= 22'h3fff7b; 
        10'b0000011011: data <= 22'h3ffff7; 
        10'b0000011100: data <= 22'h000b69; 
        10'b0000011101: data <= 22'h3ffd90; 
        10'b0000011110: data <= 22'h000290; 
        10'b0000011111: data <= 22'h000b3f; 
        10'b0000100000: data <= 22'h000452; 
        10'b0000100001: data <= 22'h00006a; 
        10'b0000100010: data <= 22'h000b2b; 
        10'b0000100011: data <= 22'h000384; 
        10'b0000100100: data <= 22'h000113; 
        10'b0000100101: data <= 22'h3ffe19; 
        10'b0000100110: data <= 22'h3ffe82; 
        10'b0000100111: data <= 22'h3ffa21; 
        10'b0000101000: data <= 22'h00099b; 
        10'b0000101001: data <= 22'h3fff4e; 
        10'b0000101010: data <= 22'h000b86; 
        10'b0000101011: data <= 22'h3ffcfe; 
        10'b0000101100: data <= 22'h0004fe; 
        10'b0000101101: data <= 22'h0008aa; 
        10'b0000101110: data <= 22'h0009bf; 
        10'b0000101111: data <= 22'h0007c7; 
        10'b0000110000: data <= 22'h000041; 
        10'b0000110001: data <= 22'h0007a9; 
        10'b0000110010: data <= 22'h3fffc6; 
        10'b0000110011: data <= 22'h000c27; 
        10'b0000110100: data <= 22'h00095f; 
        10'b0000110101: data <= 22'h3ffca0; 
        10'b0000110110: data <= 22'h3ffcb3; 
        10'b0000110111: data <= 22'h0004f6; 
        10'b0000111000: data <= 22'h000acf; 
        10'b0000111001: data <= 22'h000aa7; 
        10'b0000111010: data <= 22'h000861; 
        10'b0000111011: data <= 22'h3ffe72; 
        10'b0000111100: data <= 22'h0009b6; 
        10'b0000111101: data <= 22'h3ffb60; 
        10'b0000111110: data <= 22'h3ffc36; 
        10'b0000111111: data <= 22'h00079a; 
        10'b0001000000: data <= 22'h000669; 
        10'b0001000001: data <= 22'h3ffc3e; 
        10'b0001000010: data <= 22'h3fff2a; 
        10'b0001000011: data <= 22'h0004bb; 
        10'b0001000100: data <= 22'h3ffeb0; 
        10'b0001000101: data <= 22'h3ffd84; 
        10'b0001000110: data <= 22'h0002f8; 
        10'b0001000111: data <= 22'h0009c7; 
        10'b0001001000: data <= 22'h0007e4; 
        10'b0001001001: data <= 22'h000176; 
        10'b0001001010: data <= 22'h0003de; 
        10'b0001001011: data <= 22'h000b0c; 
        10'b0001001100: data <= 22'h000960; 
        10'b0001001101: data <= 22'h000adb; 
        10'b0001001110: data <= 22'h3ffa8b; 
        10'b0001001111: data <= 22'h000875; 
        10'b0001010000: data <= 22'h000335; 
        10'b0001010001: data <= 22'h000779; 
        10'b0001010010: data <= 22'h00066f; 
        10'b0001010011: data <= 22'h000985; 
        10'b0001010100: data <= 22'h3fff22; 
        10'b0001010101: data <= 22'h0000a4; 
        10'b0001010110: data <= 22'h0009e7; 
        10'b0001010111: data <= 22'h3ffe7f; 
        10'b0001011000: data <= 22'h00011d; 
        10'b0001011001: data <= 22'h3fff54; 
        10'b0001011010: data <= 22'h3ffc5a; 
        10'b0001011011: data <= 22'h00066f; 
        10'b0001011100: data <= 22'h00000d; 
        10'b0001011101: data <= 22'h000670; 
        10'b0001011110: data <= 22'h3ffab5; 
        10'b0001011111: data <= 22'h00014f; 
        10'b0001100000: data <= 22'h00052e; 
        10'b0001100001: data <= 22'h3ff8dc; 
        10'b0001100010: data <= 22'h0005e1; 
        10'b0001100011: data <= 22'h3ffb28; 
        10'b0001100100: data <= 22'h3ff582; 
        10'b0001100101: data <= 22'h3ff769; 
        10'b0001100110: data <= 22'h3ff8a1; 
        10'b0001100111: data <= 22'h3ffb0b; 
        10'b0001101000: data <= 22'h3ffec3; 
        10'b0001101001: data <= 22'h3ffb73; 
        10'b0001101010: data <= 22'h0003fa; 
        10'b0001101011: data <= 22'h3fff7e; 
        10'b0001101100: data <= 22'h0004cd; 
        10'b0001101101: data <= 22'h000c32; 
        10'b0001101110: data <= 22'h3ffbff; 
        10'b0001101111: data <= 22'h000509; 
        10'b0001110000: data <= 22'h000bd2; 
        10'b0001110001: data <= 22'h3ffbb3; 
        10'b0001110010: data <= 22'h000698; 
        10'b0001110011: data <= 22'h3ffafb; 
        10'b0001110100: data <= 22'h0002c3; 
        10'b0001110101: data <= 22'h3ffdba; 
        10'b0001110110: data <= 22'h000086; 
        10'b0001110111: data <= 22'h3ffb26; 
        10'b0001111000: data <= 22'h0003ae; 
        10'b0001111001: data <= 22'h3ffe45; 
        10'b0001111010: data <= 22'h3ff46c; 
        10'b0001111011: data <= 22'h3fe9ae; 
        10'b0001111100: data <= 22'h3fe88e; 
        10'b0001111101: data <= 22'h3fe99f; 
        10'b0001111110: data <= 22'h3fe554; 
        10'b0001111111: data <= 22'h3fd414; 
        10'b0010000000: data <= 22'h3fe614; 
        10'b0010000001: data <= 22'h3fec7b; 
        10'b0010000010: data <= 22'h3fef09; 
        10'b0010000011: data <= 22'h3ffb6a; 
        10'b0010000100: data <= 22'h3ff357; 
        10'b0010000101: data <= 22'h0005e8; 
        10'b0010000110: data <= 22'h0000e7; 
        10'b0010000111: data <= 22'h3ff9da; 
        10'b0010001000: data <= 22'h000b33; 
        10'b0010001001: data <= 22'h3fff9a; 
        10'b0010001010: data <= 22'h000afa; 
        10'b0010001011: data <= 22'h000aa3; 
        10'b0010001100: data <= 22'h000a14; 
        10'b0010001101: data <= 22'h000067; 
        10'b0010001110: data <= 22'h0009b7; 
        10'b0010001111: data <= 22'h3ffd59; 
        10'b0010010000: data <= 22'h3ff865; 
        10'b0010010001: data <= 22'h3ffeb2; 
        10'b0010010010: data <= 22'h3ffa2c; 
        10'b0010010011: data <= 22'h3ffddf; 
        10'b0010010100: data <= 22'h3ff91a; 
        10'b0010010101: data <= 22'h3feff9; 
        10'b0010010110: data <= 22'h3fd8a5; 
        10'b0010010111: data <= 22'h3fcfb3; 
        10'b0010011000: data <= 22'h3fc335; 
        10'b0010011001: data <= 22'h3fb8c8; 
        10'b0010011010: data <= 22'h3fa724; 
        10'b0010011011: data <= 22'h3fa7ce; 
        10'b0010011100: data <= 22'h3fa384; 
        10'b0010011101: data <= 22'h3fae68; 
        10'b0010011110: data <= 22'h3fbadc; 
        10'b0010011111: data <= 22'h3fcb65; 
        10'b0010100000: data <= 22'h3fdaa0; 
        10'b0010100001: data <= 22'h3ff2ab; 
        10'b0010100010: data <= 22'h3feb63; 
        10'b0010100011: data <= 22'h3ffd6c; 
        10'b0010100100: data <= 22'h000905; 
        10'b0010100101: data <= 22'h000732; 
        10'b0010100110: data <= 22'h3ffe27; 
        10'b0010100111: data <= 22'h000068; 
        10'b0010101000: data <= 22'h000861; 
        10'b0010101001: data <= 22'h000b79; 
        10'b0010101010: data <= 22'h0000ce; 
        10'b0010101011: data <= 22'h0001dd; 
        10'b0010101100: data <= 22'h000c6a; 
        10'b0010101101: data <= 22'h000ec8; 
        10'b0010101110: data <= 22'h00114d; 
        10'b0010101111: data <= 22'h001a0b; 
        10'b0010110000: data <= 22'h0026a2; 
        10'b0010110001: data <= 22'h001ef1; 
        10'b0010110010: data <= 22'h0020ee; 
        10'b0010110011: data <= 22'h0005eb; 
        10'b0010110100: data <= 22'h3fe596; 
        10'b0010110101: data <= 22'h3fc892; 
        10'b0010110110: data <= 22'h3fc627; 
        10'b0010110111: data <= 22'h3fe1f4; 
        10'b0010111000: data <= 22'h3fedc2; 
        10'b0010111001: data <= 22'h3fea58; 
        10'b0010111010: data <= 22'h3fe5bf; 
        10'b0010111011: data <= 22'h3fe1a0; 
        10'b0010111100: data <= 22'h3fd204; 
        10'b0010111101: data <= 22'h3feebf; 
        10'b0010111110: data <= 22'h3fdfc5; 
        10'b0010111111: data <= 22'h3fe88b; 
        10'b0011000000: data <= 22'h3ff04c; 
        10'b0011000001: data <= 22'h3ffabc; 
        10'b0011000010: data <= 22'h3ffa8e; 
        10'b0011000011: data <= 22'h000144; 
        10'b0011000100: data <= 22'h0007a2; 
        10'b0011000101: data <= 22'h000b91; 
        10'b0011000110: data <= 22'h000985; 
        10'b0011000111: data <= 22'h001682; 
        10'b0011001000: data <= 22'h001b4a; 
        10'b0011001001: data <= 22'h00188a; 
        10'b0011001010: data <= 22'h00238b; 
        10'b0011001011: data <= 22'h003654; 
        10'b0011001100: data <= 22'h004a6a; 
        10'b0011001101: data <= 22'h003af5; 
        10'b0011001110: data <= 22'h0028ad; 
        10'b0011001111: data <= 22'h002ccd; 
        10'b0011010000: data <= 22'h002fb9; 
        10'b0011010001: data <= 22'h00092c; 
        10'b0011010010: data <= 22'h0006c6; 
        10'b0011010011: data <= 22'h001115; 
        10'b0011010100: data <= 22'h00325e; 
        10'b0011010101: data <= 22'h0037ff; 
        10'b0011010110: data <= 22'h0025f2; 
        10'b0011010111: data <= 22'h001e6c; 
        10'b0011011000: data <= 22'h00076c; 
        10'b0011011001: data <= 22'h3ff795; 
        10'b0011011010: data <= 22'h0003f4; 
        10'b0011011011: data <= 22'h3ff6ed; 
        10'b0011011100: data <= 22'h3ff784; 
        10'b0011011101: data <= 22'h3fff8d; 
        10'b0011011110: data <= 22'h000601; 
        10'b0011011111: data <= 22'h3ffdbf; 
        10'b0011100000: data <= 22'h3ffa29; 
        10'b0011100001: data <= 22'h000c1f; 
        10'b0011100010: data <= 22'h0004ae; 
        10'b0011100011: data <= 22'h001302; 
        10'b0011100100: data <= 22'h00267d; 
        10'b0011100101: data <= 22'h0022b6; 
        10'b0011100110: data <= 22'h002e79; 
        10'b0011100111: data <= 22'h00536e; 
        10'b0011101000: data <= 22'h003829; 
        10'b0011101001: data <= 22'h0026af; 
        10'b0011101010: data <= 22'h003138; 
        10'b0011101011: data <= 22'h0041ec; 
        10'b0011101100: data <= 22'h003ea8; 
        10'b0011101101: data <= 22'h001f86; 
        10'b0011101110: data <= 22'h00126c; 
        10'b0011101111: data <= 22'h001993; 
        10'b0011110000: data <= 22'h002c6d; 
        10'b0011110001: data <= 22'h00444c; 
        10'b0011110010: data <= 22'h002ece; 
        10'b0011110011: data <= 22'h002818; 
        10'b0011110100: data <= 22'h002001; 
        10'b0011110101: data <= 22'h0000bf; 
        10'b0011110110: data <= 22'h001365; 
        10'b0011110111: data <= 22'h001076; 
        10'b0011111000: data <= 22'h3ff442; 
        10'b0011111001: data <= 22'h3ffa65; 
        10'b0011111010: data <= 22'h00067e; 
        10'b0011111011: data <= 22'h0009fb; 
        10'b0011111100: data <= 22'h000527; 
        10'b0011111101: data <= 22'h0009a7; 
        10'b0011111110: data <= 22'h000cf6; 
        10'b0011111111: data <= 22'h001b68; 
        10'b0100000000: data <= 22'h0025b7; 
        10'b0100000001: data <= 22'h002ad5; 
        10'b0100000010: data <= 22'h000fb7; 
        10'b0100000011: data <= 22'h0014e6; 
        10'b0100000100: data <= 22'h0017b1; 
        10'b0100000101: data <= 22'h000faa; 
        10'b0100000110: data <= 22'h002665; 
        10'b0100000111: data <= 22'h002f0b; 
        10'b0100001000: data <= 22'h003bfb; 
        10'b0100001001: data <= 22'h0030cc; 
        10'b0100001010: data <= 22'h0045e9; 
        10'b0100001011: data <= 22'h00560d; 
        10'b0100001100: data <= 22'h004f46; 
        10'b0100001101: data <= 22'h005878; 
        10'b0100001110: data <= 22'h0039c2; 
        10'b0100001111: data <= 22'h003ad2; 
        10'b0100010000: data <= 22'h003176; 
        10'b0100010001: data <= 22'h002942; 
        10'b0100010010: data <= 22'h001388; 
        10'b0100010011: data <= 22'h3ff8e5; 
        10'b0100010100: data <= 22'h3ff3fd; 
        10'b0100010101: data <= 22'h3ffa1d; 
        10'b0100010110: data <= 22'h000538; 
        10'b0100010111: data <= 22'h3ffd53; 
        10'b0100011000: data <= 22'h0001ff; 
        10'b0100011001: data <= 22'h000a86; 
        10'b0100011010: data <= 22'h000bac; 
        10'b0100011011: data <= 22'h002213; 
        10'b0100011100: data <= 22'h002709; 
        10'b0100011101: data <= 22'h002073; 
        10'b0100011110: data <= 22'h0005fb; 
        10'b0100011111: data <= 22'h0009c2; 
        10'b0100100000: data <= 22'h3ff2e0; 
        10'b0100100001: data <= 22'h3fff81; 
        10'b0100100010: data <= 22'h0017d0; 
        10'b0100100011: data <= 22'h0029ee; 
        10'b0100100100: data <= 22'h001d2c; 
        10'b0100100101: data <= 22'h0043e3; 
        10'b0100100110: data <= 22'h00575a; 
        10'b0100100111: data <= 22'h006b49; 
        10'b0100101000: data <= 22'h007a28; 
        10'b0100101001: data <= 22'h005a88; 
        10'b0100101010: data <= 22'h00474d; 
        10'b0100101011: data <= 22'h004a29; 
        10'b0100101100: data <= 22'h00411c; 
        10'b0100101101: data <= 22'h00375b; 
        10'b0100101110: data <= 22'h001879; 
        10'b0100101111: data <= 22'h3ff603; 
        10'b0100110000: data <= 22'h3fef79; 
        10'b0100110001: data <= 22'h3ff94d; 
        10'b0100110010: data <= 22'h000141; 
        10'b0100110011: data <= 22'h3ffd7f; 
        10'b0100110100: data <= 22'h000943; 
        10'b0100110101: data <= 22'h000681; 
        10'b0100110110: data <= 22'h000bcf; 
        10'b0100110111: data <= 22'h0022e7; 
        10'b0100111000: data <= 22'h002a0f; 
        10'b0100111001: data <= 22'h0014da; 
        10'b0100111010: data <= 22'h000793; 
        10'b0100111011: data <= 22'h0006cc; 
        10'b0100111100: data <= 22'h0001f3; 
        10'b0100111101: data <= 22'h001940; 
        10'b0100111110: data <= 22'h000d06; 
        10'b0100111111: data <= 22'h00106d; 
        10'b0101000000: data <= 22'h001b25; 
        10'b0101000001: data <= 22'h001ae6; 
        10'b0101000010: data <= 22'h001bf8; 
        10'b0101000011: data <= 22'h00521b; 
        10'b0101000100: data <= 22'h006a9e; 
        10'b0101000101: data <= 22'h00470d; 
        10'b0101000110: data <= 22'h0047c1; 
        10'b0101000111: data <= 22'h00372c; 
        10'b0101001000: data <= 22'h00359a; 
        10'b0101001001: data <= 22'h0021b8; 
        10'b0101001010: data <= 22'h001859; 
        10'b0101001011: data <= 22'h3ff78a; 
        10'b0101001100: data <= 22'h3fe75f; 
        10'b0101001101: data <= 22'h3fff50; 
        10'b0101001110: data <= 22'h00025a; 
        10'b0101001111: data <= 22'h000ac9; 
        10'b0101010000: data <= 22'h000840; 
        10'b0101010001: data <= 22'h3fff67; 
        10'b0101010010: data <= 22'h0005df; 
        10'b0101010011: data <= 22'h0015fb; 
        10'b0101010100: data <= 22'h0018ae; 
        10'b0101010101: data <= 22'h000410; 
        10'b0101010110: data <= 22'h000584; 
        10'b0101010111: data <= 22'h00177c; 
        10'b0101011000: data <= 22'h001019; 
        10'b0101011001: data <= 22'h3fff10; 
        10'b0101011010: data <= 22'h3feccc; 
        10'b0101011011: data <= 22'h3fcce1; 
        10'b0101011100: data <= 22'h3f93ef; 
        10'b0101011101: data <= 22'h3f58bc; 
        10'b0101011110: data <= 22'h3f82ce; 
        10'b0101011111: data <= 22'h0002b9; 
        10'b0101100000: data <= 22'h0046b6; 
        10'b0101100001: data <= 22'h00402e; 
        10'b0101100010: data <= 22'h00193f; 
        10'b0101100011: data <= 22'h000912; 
        10'b0101100100: data <= 22'h0001b2; 
        10'b0101100101: data <= 22'h3ff6c0; 
        10'b0101100110: data <= 22'h3ff79c; 
        10'b0101100111: data <= 22'h3ff0e0; 
        10'b0101101000: data <= 22'h3ff51a; 
        10'b0101101001: data <= 22'h000a33; 
        10'b0101101010: data <= 22'h00072b; 
        10'b0101101011: data <= 22'h000017; 
        10'b0101101100: data <= 22'h0008ef; 
        10'b0101101101: data <= 22'h000542; 
        10'b0101101110: data <= 22'h0009a2; 
        10'b0101101111: data <= 22'h0013f2; 
        10'b0101110000: data <= 22'h00076e; 
        10'b0101110001: data <= 22'h000330; 
        10'b0101110010: data <= 22'h3ff974; 
        10'b0101110011: data <= 22'h00044c; 
        10'b0101110100: data <= 22'h3ffcfc; 
        10'b0101110101: data <= 22'h3fef9f; 
        10'b0101110110: data <= 22'h3fca5d; 
        10'b0101110111: data <= 22'h3f8eea; 
        10'b0101111000: data <= 22'h3f3976; 
        10'b0101111001: data <= 22'h3f223c; 
        10'b0101111010: data <= 22'h3f8956; 
        10'b0101111011: data <= 22'h3ff071; 
        10'b0101111100: data <= 22'h002418; 
        10'b0101111101: data <= 22'h001747; 
        10'b0101111110: data <= 22'h000509; 
        10'b0101111111: data <= 22'h000a96; 
        10'b0110000000: data <= 22'h3fea42; 
        10'b0110000001: data <= 22'h3fe42e; 
        10'b0110000010: data <= 22'h3ff979; 
        10'b0110000011: data <= 22'h00020e; 
        10'b0110000100: data <= 22'h3ffab7; 
        10'b0110000101: data <= 22'h3ffbc7; 
        10'b0110000110: data <= 22'h0005a7; 
        10'b0110000111: data <= 22'h3ffa83; 
        10'b0110001000: data <= 22'h3ffd9a; 
        10'b0110001001: data <= 22'h0004c4; 
        10'b0110001010: data <= 22'h0011da; 
        10'b0110001011: data <= 22'h00163d; 
        10'b0110001100: data <= 22'h000e19; 
        10'b0110001101: data <= 22'h00105f; 
        10'b0110001110: data <= 22'h3ffa93; 
        10'b0110001111: data <= 22'h3ff498; 
        10'b0110010000: data <= 22'h3fe6d5; 
        10'b0110010001: data <= 22'h3fc50b; 
        10'b0110010010: data <= 22'h3fa958; 
        10'b0110010011: data <= 22'h3f79f2; 
        10'b0110010100: data <= 22'h3f542b; 
        10'b0110010101: data <= 22'h3f6f0d; 
        10'b0110010110: data <= 22'h3fcadc; 
        10'b0110010111: data <= 22'h00013c; 
        10'b0110011000: data <= 22'h000b0b; 
        10'b0110011001: data <= 22'h0016e3; 
        10'b0110011010: data <= 22'h0041ae; 
        10'b0110011011: data <= 22'h004698; 
        10'b0110011100: data <= 22'h002a79; 
        10'b0110011101: data <= 22'h001b21; 
        10'b0110011110: data <= 22'h001b49; 
        10'b0110011111: data <= 22'h0017a9; 
        10'b0110100000: data <= 22'h000801; 
        10'b0110100001: data <= 22'h000260; 
        10'b0110100010: data <= 22'h3ffc38; 
        10'b0110100011: data <= 22'h3ffc92; 
        10'b0110100100: data <= 22'h0005c2; 
        10'b0110100101: data <= 22'h00087e; 
        10'b0110100110: data <= 22'h00031d; 
        10'b0110100111: data <= 22'h00086c; 
        10'b0110101000: data <= 22'h000865; 
        10'b0110101001: data <= 22'h3fe837; 
        10'b0110101010: data <= 22'h3ff565; 
        10'b0110101011: data <= 22'h3ff143; 
        10'b0110101100: data <= 22'h3fc0ba; 
        10'b0110101101: data <= 22'h3fb339; 
        10'b0110101110: data <= 22'h3f99f0; 
        10'b0110101111: data <= 22'h3f8b0c; 
        10'b0110110000: data <= 22'h3f809c; 
        10'b0110110001: data <= 22'h3fa21d; 
        10'b0110110010: data <= 22'h3fc92a; 
        10'b0110110011: data <= 22'h0001ad; 
        10'b0110110100: data <= 22'h0005fb; 
        10'b0110110101: data <= 22'h005955; 
        10'b0110110110: data <= 22'h006896; 
        10'b0110110111: data <= 22'h005630; 
        10'b0110111000: data <= 22'h004c8a; 
        10'b0110111001: data <= 22'h0041d8; 
        10'b0110111010: data <= 22'h002a8d; 
        10'b0110111011: data <= 22'h001338; 
        10'b0110111100: data <= 22'h3fff34; 
        10'b0110111101: data <= 22'h3ffab1; 
        10'b0110111110: data <= 22'h00016b; 
        10'b0110111111: data <= 22'h000929; 
        10'b0111000000: data <= 22'h0005b4; 
        10'b0111000001: data <= 22'h000b55; 
        10'b0111000010: data <= 22'h3fff10; 
        10'b0111000011: data <= 22'h000be5; 
        10'b0111000100: data <= 22'h00095d; 
        10'b0111000101: data <= 22'h3ff558; 
        10'b0111000110: data <= 22'h3ff0f1; 
        10'b0111000111: data <= 22'h3ffdd6; 
        10'b0111001000: data <= 22'h3fcd10; 
        10'b0111001001: data <= 22'h3fc681; 
        10'b0111001010: data <= 22'h3fa36d; 
        10'b0111001011: data <= 22'h3f91f3; 
        10'b0111001100: data <= 22'h3fbb02; 
        10'b0111001101: data <= 22'h3fd968; 
        10'b0111001110: data <= 22'h3fc80d; 
        10'b0111001111: data <= 22'h001cc8; 
        10'b0111010000: data <= 22'h0022d1; 
        10'b0111010001: data <= 22'h004b95; 
        10'b0111010010: data <= 22'h0040c1; 
        10'b0111010011: data <= 22'h0043d9; 
        10'b0111010100: data <= 22'h0035fc; 
        10'b0111010101: data <= 22'h00291c; 
        10'b0111010110: data <= 22'h00081c; 
        10'b0111010111: data <= 22'h3fef15; 
        10'b0111011000: data <= 22'h3ff581; 
        10'b0111011001: data <= 22'h3ffa08; 
        10'b0111011010: data <= 22'h00066c; 
        10'b0111011011: data <= 22'h000b2e; 
        10'b0111011100: data <= 22'h00005b; 
        10'b0111011101: data <= 22'h000170; 
        10'b0111011110: data <= 22'h0006df; 
        10'b0111011111: data <= 22'h3fff88; 
        10'b0111100000: data <= 22'h000243; 
        10'b0111100001: data <= 22'h3ff933; 
        10'b0111100010: data <= 22'h3fddac; 
        10'b0111100011: data <= 22'h3fd2c4; 
        10'b0111100100: data <= 22'h3fc73b; 
        10'b0111100101: data <= 22'h3fd123; 
        10'b0111100110: data <= 22'h3fc1e1; 
        10'b0111100111: data <= 22'h3fd1e8; 
        10'b0111101000: data <= 22'h3ff146; 
        10'b0111101001: data <= 22'h000b7f; 
        10'b0111101010: data <= 22'h000686; 
        10'b0111101011: data <= 22'h000b74; 
        10'b0111101100: data <= 22'h3ff937; 
        10'b0111101101: data <= 22'h001229; 
        10'b0111101110: data <= 22'h001031; 
        10'b0111101111: data <= 22'h000b82; 
        10'b0111110000: data <= 22'h00061a; 
        10'b0111110001: data <= 22'h3ff697; 
        10'b0111110010: data <= 22'h3feb1d; 
        10'b0111110011: data <= 22'h3ff699; 
        10'b0111110100: data <= 22'h3ff7d5; 
        10'b0111110101: data <= 22'h3ff996; 
        10'b0111110110: data <= 22'h3ffc8d; 
        10'b0111110111: data <= 22'h3ffce6; 
        10'b0111111000: data <= 22'h3ffcd9; 
        10'b0111111001: data <= 22'h3ffefb; 
        10'b0111111010: data <= 22'h0007c7; 
        10'b0111111011: data <= 22'h000267; 
        10'b0111111100: data <= 22'h3ff219; 
        10'b0111111101: data <= 22'h3fdeef; 
        10'b0111111110: data <= 22'h3fc95e; 
        10'b0111111111: data <= 22'h3fbbf9; 
        10'b1000000000: data <= 22'h3fc0d9; 
        10'b1000000001: data <= 22'h3fc4e2; 
        10'b1000000010: data <= 22'h3fb40e; 
        10'b1000000011: data <= 22'h3fe5e0; 
        10'b1000000100: data <= 22'h3ff81c; 
        10'b1000000101: data <= 22'h0000ed; 
        10'b1000000110: data <= 22'h00155d; 
        10'b1000000111: data <= 22'h3fe972; 
        10'b1000001000: data <= 22'h3fe44d; 
        10'b1000001001: data <= 22'h3ff0b1; 
        10'b1000001010: data <= 22'h3fdd1e; 
        10'b1000001011: data <= 22'h3fea99; 
        10'b1000001100: data <= 22'h3fdc13; 
        10'b1000001101: data <= 22'h3fc8cd; 
        10'b1000001110: data <= 22'h3fd79f; 
        10'b1000001111: data <= 22'h3fe680; 
        10'b1000010000: data <= 22'h3febf2; 
        10'b1000010001: data <= 22'h000214; 
        10'b1000010010: data <= 22'h3ffdcb; 
        10'b1000010011: data <= 22'h000079; 
        10'b1000010100: data <= 22'h000ad2; 
        10'b1000010101: data <= 22'h000b97; 
        10'b1000010110: data <= 22'h000a9c; 
        10'b1000010111: data <= 22'h00054a; 
        10'b1000011000: data <= 22'h3ff69d; 
        10'b1000011001: data <= 22'h3fd502; 
        10'b1000011010: data <= 22'h3fbb2c; 
        10'b1000011011: data <= 22'h3fb627; 
        10'b1000011100: data <= 22'h3fb42e; 
        10'b1000011101: data <= 22'h3fb3b5; 
        10'b1000011110: data <= 22'h3fcc56; 
        10'b1000011111: data <= 22'h3fdacf; 
        10'b1000100000: data <= 22'h3fe9c1; 
        10'b1000100001: data <= 22'h0009a5; 
        10'b1000100010: data <= 22'h001e38; 
        10'b1000100011: data <= 22'h3fe072; 
        10'b1000100100: data <= 22'h3fe138; 
        10'b1000100101: data <= 22'h3fd922; 
        10'b1000100110: data <= 22'h3fc237; 
        10'b1000100111: data <= 22'h3fc578; 
        10'b1000101000: data <= 22'h3fb7e8; 
        10'b1000101001: data <= 22'h3fbd70; 
        10'b1000101010: data <= 22'h3fcd55; 
        10'b1000101011: data <= 22'h3fdd18; 
        10'b1000101100: data <= 22'h3fee4d; 
        10'b1000101101: data <= 22'h3ff970; 
        10'b1000101110: data <= 22'h000b19; 
        10'b1000101111: data <= 22'h3ffaf8; 
        10'b1000110000: data <= 22'h3ffa3a; 
        10'b1000110001: data <= 22'h3ffd62; 
        10'b1000110010: data <= 22'h00048f; 
        10'b1000110011: data <= 22'h3ffe24; 
        10'b1000110100: data <= 22'h3ff521; 
        10'b1000110101: data <= 22'h3fded1; 
        10'b1000110110: data <= 22'h3fbaa7; 
        10'b1000110111: data <= 22'h3fb7ab; 
        10'b1000111000: data <= 22'h3fbbc4; 
        10'b1000111001: data <= 22'h3fbd5c; 
        10'b1000111010: data <= 22'h3fd189; 
        10'b1000111011: data <= 22'h3fd010; 
        10'b1000111100: data <= 22'h000378; 
        10'b1000111101: data <= 22'h0004c3; 
        10'b1000111110: data <= 22'h00100a; 
        10'b1000111111: data <= 22'h3fd5b7; 
        10'b1001000000: data <= 22'h3fcb27; 
        10'b1001000001: data <= 22'h3fbaf5; 
        10'b1001000010: data <= 22'h3fa0b4; 
        10'b1001000011: data <= 22'h3fc359; 
        10'b1001000100: data <= 22'h3fac78; 
        10'b1001000101: data <= 22'h3fc04c; 
        10'b1001000110: data <= 22'h3fd1eb; 
        10'b1001000111: data <= 22'h3fec68; 
        10'b1001001000: data <= 22'h3ff2ea; 
        10'b1001001001: data <= 22'h0009e3; 
        10'b1001001010: data <= 22'h000964; 
        10'b1001001011: data <= 22'h000660; 
        10'b1001001100: data <= 22'h0008e8; 
        10'b1001001101: data <= 22'h000955; 
        10'b1001001110: data <= 22'h000218; 
        10'b1001001111: data <= 22'h3ff3ce; 
        10'b1001010000: data <= 22'h3ff9d1; 
        10'b1001010001: data <= 22'h3fe26f; 
        10'b1001010010: data <= 22'h3fdd57; 
        10'b1001010011: data <= 22'h3fce0b; 
        10'b1001010100: data <= 22'h3fd2fd; 
        10'b1001010101: data <= 22'h3fe53c; 
        10'b1001010110: data <= 22'h3fd9e8; 
        10'b1001010111: data <= 22'h3fe0f2; 
        10'b1001011000: data <= 22'h3ff21d; 
        10'b1001011001: data <= 22'h0001e2; 
        10'b1001011010: data <= 22'h3ff7aa; 
        10'b1001011011: data <= 22'h3fe380; 
        10'b1001011100: data <= 22'h3fdf36; 
        10'b1001011101: data <= 22'h3fbbe5; 
        10'b1001011110: data <= 22'h3fbc2a; 
        10'b1001011111: data <= 22'h3fbc06; 
        10'b1001100000: data <= 22'h3fb867; 
        10'b1001100001: data <= 22'h3fc364; 
        10'b1001100010: data <= 22'h3fdc64; 
        10'b1001100011: data <= 22'h3fe511; 
        10'b1001100100: data <= 22'h3ffed1; 
        10'b1001100101: data <= 22'h000427; 
        10'b1001100110: data <= 22'h0008fd; 
        10'b1001100111: data <= 22'h3ffe10; 
        10'b1001101000: data <= 22'h000308; 
        10'b1001101001: data <= 22'h0000b4; 
        10'b1001101010: data <= 22'h000262; 
        10'b1001101011: data <= 22'h3ff87e; 
        10'b1001101100: data <= 22'h3ffc98; 
        10'b1001101101: data <= 22'h000466; 
        10'b1001101110: data <= 22'h3ff52a; 
        10'b1001101111: data <= 22'h000561; 
        10'b1001110000: data <= 22'h000890; 
        10'b1001110001: data <= 22'h3ff250; 
        10'b1001110010: data <= 22'h3fe5f2; 
        10'b1001110011: data <= 22'h3fd38c; 
        10'b1001110100: data <= 22'h3fd673; 
        10'b1001110101: data <= 22'h3fef3e; 
        10'b1001110110: data <= 22'h0004fa; 
        10'b1001110111: data <= 22'h0004e7; 
        10'b1001111000: data <= 22'h3fe62a; 
        10'b1001111001: data <= 22'h3fe001; 
        10'b1001111010: data <= 22'h3fc97d; 
        10'b1001111011: data <= 22'h3fc982; 
        10'b1001111100: data <= 22'h3fc296; 
        10'b1001111101: data <= 22'h3fca3e; 
        10'b1001111110: data <= 22'h3fe4b3; 
        10'b1001111111: data <= 22'h3ff6c5; 
        10'b1010000000: data <= 22'h0005f2; 
        10'b1010000001: data <= 22'h3ffa32; 
        10'b1010000010: data <= 22'h0002d7; 
        10'b1010000011: data <= 22'h00002e; 
        10'b1010000100: data <= 22'h000433; 
        10'b1010000101: data <= 22'h00087d; 
        10'b1010000110: data <= 22'h3ff972; 
        10'b1010000111: data <= 22'h3ffa09; 
        10'b1010001000: data <= 22'h000b43; 
        10'b1010001001: data <= 22'h000f12; 
        10'b1010001010: data <= 22'h0020ca; 
        10'b1010001011: data <= 22'h002bba; 
        10'b1010001100: data <= 22'h0014e2; 
        10'b1010001101: data <= 22'h000429; 
        10'b1010001110: data <= 22'h3ff322; 
        10'b1010001111: data <= 22'h3fe245; 
        10'b1010010000: data <= 22'h3fe7b0; 
        10'b1010010001: data <= 22'h0001af; 
        10'b1010010010: data <= 22'h001109; 
        10'b1010010011: data <= 22'h000fb2; 
        10'b1010010100: data <= 22'h3ff974; 
        10'b1010010101: data <= 22'h3ff64c; 
        10'b1010010110: data <= 22'h3fdd1f; 
        10'b1010010111: data <= 22'h3fcf54; 
        10'b1010011000: data <= 22'h3fce34; 
        10'b1010011001: data <= 22'h3fd920; 
        10'b1010011010: data <= 22'h3fdfee; 
        10'b1010011011: data <= 22'h3feb17; 
        10'b1010011100: data <= 22'h3ff6c4; 
        10'b1010011101: data <= 22'h0000b1; 
        10'b1010011110: data <= 22'h00009b; 
        10'b1010011111: data <= 22'h3ffc8f; 
        10'b1010100000: data <= 22'h3fffeb; 
        10'b1010100001: data <= 22'h3ffedb; 
        10'b1010100010: data <= 22'h00031e; 
        10'b1010100011: data <= 22'h00074e; 
        10'b1010100100: data <= 22'h000fa6; 
        10'b1010100101: data <= 22'h0023fc; 
        10'b1010100110: data <= 22'h003677; 
        10'b1010100111: data <= 22'h003d60; 
        10'b1010101000: data <= 22'h003421; 
        10'b1010101001: data <= 22'h001ae2; 
        10'b1010101010: data <= 22'h0039eb; 
        10'b1010101011: data <= 22'h002233; 
        10'b1010101100: data <= 22'h001dab; 
        10'b1010101101: data <= 22'h0029c9; 
        10'b1010101110: data <= 22'h0019b9; 
        10'b1010101111: data <= 22'h00251e; 
        10'b1010110000: data <= 22'h0015fb; 
        10'b1010110001: data <= 22'h001127; 
        10'b1010110010: data <= 22'h3ffee7; 
        10'b1010110011: data <= 22'h3ff001; 
        10'b1010110100: data <= 22'h3fef00; 
        10'b1010110101: data <= 22'h3feb5c; 
        10'b1010110110: data <= 22'h3fe8b2; 
        10'b1010110111: data <= 22'h3feac9; 
        10'b1010111000: data <= 22'h00033e; 
        10'b1010111001: data <= 22'h3ffe54; 
        10'b1010111010: data <= 22'h3ffa74; 
        10'b1010111011: data <= 22'h00065b; 
        10'b1010111100: data <= 22'h3ffa55; 
        10'b1010111101: data <= 22'h00052f; 
        10'b1010111110: data <= 22'h000963; 
        10'b1010111111: data <= 22'h0008cb; 
        10'b1011000000: data <= 22'h000519; 
        10'b1011000001: data <= 22'h0011f0; 
        10'b1011000010: data <= 22'h001a8e; 
        10'b1011000011: data <= 22'h00290c; 
        10'b1011000100: data <= 22'h003f74; 
        10'b1011000101: data <= 22'h003df0; 
        10'b1011000110: data <= 22'h004953; 
        10'b1011000111: data <= 22'h00443c; 
        10'b1011001000: data <= 22'h003cce; 
        10'b1011001001: data <= 22'h00302a; 
        10'b1011001010: data <= 22'h003132; 
        10'b1011001011: data <= 22'h003422; 
        10'b1011001100: data <= 22'h002bb1; 
        10'b1011001101: data <= 22'h0028d4; 
        10'b1011001110: data <= 22'h0020e9; 
        10'b1011001111: data <= 22'h000b4b; 
        10'b1011010000: data <= 22'h3ff222; 
        10'b1011010001: data <= 22'h0001df; 
        10'b1011010010: data <= 22'h3ff926; 
        10'b1011010011: data <= 22'h3ffaf8; 
        10'b1011010100: data <= 22'h3ffe66; 
        10'b1011010101: data <= 22'h000323; 
        10'b1011010110: data <= 22'h000c6e; 
        10'b1011010111: data <= 22'h000811; 
        10'b1011011000: data <= 22'h3ffb97; 
        10'b1011011001: data <= 22'h000263; 
        10'b1011011010: data <= 22'h000bbf; 
        10'b1011011011: data <= 22'h3ffe00; 
        10'b1011011100: data <= 22'h3ffc03; 
        10'b1011011101: data <= 22'h000afb; 
        10'b1011011110: data <= 22'h0000cb; 
        10'b1011011111: data <= 22'h000a08; 
        10'b1011100000: data <= 22'h000992; 
        10'b1011100001: data <= 22'h000157; 
        10'b1011100010: data <= 22'h000dcd; 
        10'b1011100011: data <= 22'h001457; 
        10'b1011100100: data <= 22'h0005dd; 
        10'b1011100101: data <= 22'h001175; 
        10'b1011100110: data <= 22'h002570; 
        10'b1011100111: data <= 22'h002e3a; 
        10'b1011101000: data <= 22'h002477; 
        10'b1011101001: data <= 22'h002eb8; 
        10'b1011101010: data <= 22'h001aa1; 
        10'b1011101011: data <= 22'h000c93; 
        10'b1011101100: data <= 22'h00006a; 
        10'b1011101101: data <= 22'h0004d5; 
        10'b1011101110: data <= 22'h3ffeb4; 
        10'b1011101111: data <= 22'h0002b2; 
        10'b1011110000: data <= 22'h00008a; 
        10'b1011110001: data <= 22'h3ffcdd; 
        10'b1011110010: data <= 22'h3fff42; 
        10'b1011110011: data <= 22'h3ffe6e; 
        10'b1011110100: data <= 22'h3ffa33; 
        10'b1011110101: data <= 22'h0004bd; 
        10'b1011110110: data <= 22'h000337; 
        10'b1011110111: data <= 22'h0005e6; 
        10'b1011111000: data <= 22'h000804; 
        10'b1011111001: data <= 22'h0004ca; 
        10'b1011111010: data <= 22'h000213; 
        10'b1011111011: data <= 22'h0000dc; 
        10'b1011111100: data <= 22'h000d24; 
        10'b1011111101: data <= 22'h000810; 
        10'b1011111110: data <= 22'h000261; 
        10'b1011111111: data <= 22'h000824; 
        10'b1100000000: data <= 22'h0003f1; 
        10'b1100000001: data <= 22'h000f31; 
        10'b1100000010: data <= 22'h000910; 
        10'b1100000011: data <= 22'h0006eb; 
        10'b1100000100: data <= 22'h00151f; 
        10'b1100000101: data <= 22'h000727; 
        10'b1100000110: data <= 22'h000655; 
        10'b1100000111: data <= 22'h000ea8; 
        10'b1100001000: data <= 22'h0001be; 
        10'b1100001001: data <= 22'h3ffd87; 
        10'b1100001010: data <= 22'h000bf6; 
        10'b1100001011: data <= 22'h00068e; 
        10'b1100001100: data <= 22'h00030b; 
        10'b1100001101: data <= 22'h3ffdd1; 
        10'b1100001110: data <= 22'h3ffb1b; 
        10'b1100001111: data <= 22'h0007f6; 
      endcase 
    end 
  end 
endgenerate 
assign dout = data; 
endmodule
