`timescale 1ns / 1ps

module tb_full_connected_layer();

parameter int BITS = 24;
parameter int WIDTH = 784;
parameter int HEIGHT = 10;

logic clk;
logic reset_nn;
logic [31:0] reset_reg, MAC0_out;
logic [9:0] pixel_counter;
logic [BITS - 1 : 0] input_pixel, MEM0_out;
logic [BITS - 1 : 0] predict_num;
logic new_data;

// Internal signal
(* ASYNC_REG = "TRUE"*) reg [2:0] sync;
wire nn_en;

// Enable for NN (toggle synchronizer)
always @(posedge clk) begin
    sync[2] <= sync[1];
    sync[1] <= sync[0];
    sync[0] <= new_data;
end

assign nn_en = ((~sync[2]) & sync[1]);
               
assign reset_nn = reset_reg[0];               
nn #( 
    .BITS(BITS), 
    .WIDTH(WIDTH), 
    .HEIGHT(HEIGHT)
) dut (
    .clk(clk),
    .reset(reset_nn),
    .en(nn_en),
    .nn_in(input_pixel),
    .CNT_out(pixel_counter),
    .nn_out(predict_num),
    .*
);

logic [BITS - 1 : 0] arr_6 [0 : WIDTH-1]= '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1140, 3067, 1959, 1124, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2361, 4063, 4079, 3067, 176, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1188, 3887, 4063, 4079, 4063, 417, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 562, 3838, 4063, 4063, 4079, 2602, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2345, 4063, 4063, 4063, 3003, 594, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2232, 3742, 4063, 4063, 4063, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3003, 4063, 4063, 4031, 2280, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 690, 3678, 4063, 4063, 2489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2329, 4063, 4063, 4063, 1718, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3228, 4063, 4063, 4063, 1718, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 626, 3646, 4079, 4079, 4079, 2827, 1943, 1959, 96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1301, 4063, 4063, 4063, 4063, 4063, 4063, 4079, 3887, 3067, 273, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1301, 4063, 4063, 4063, 4063, 4063, 4063, 4079, 4063, 4063, 1911, 321, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 883, 3806, 4063, 4063, 4063, 3308, 2778, 4079, 4063, 4063, 4063, 3003, 337, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3228, 4063, 4063, 4063, 2329, 514, 851, 3341, 4063, 4063, 4063, 1638, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 963, 3855, 4063, 4063, 4063, 4063, 3501, 867, 3357, 4063, 4063, 4063, 3196, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 417, 3148, 4063, 4063, 4063, 4063, 4063, 4096, 4063, 4063, 4063, 3903, 1574, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 401, 3164, 4063, 4063, 4063, 4063, 4096, 4063, 4063, 4063, 2762, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 369, 2056, 3871, 4063, 4063, 4096, 4063, 4063, 3196, 353, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 208, 1927, 3051, 2939, 3148, 1927, 305, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}; // 6
//logic [BITS - 1 : 0] arr_6 [0 : WIDTH-1]= '{1, 2, 3, 4, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1140, 3067, 1959, 1124, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2361, 4063, 4079, 3067, 176, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1188, 3887, 4063, 4079, 4063, 417, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 562, 3838, 4063, 4063, 4079, 2602, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2345, 4063, 4063, 4063, 3003, 594, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2232, 3742, 4063, 4063, 4063, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3003, 4063, 4063, 4031, 2280, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 690, 3678, 4063, 4063, 2489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2329, 4063, 4063, 4063, 1718, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3228, 4063, 4063, 4063, 1718, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 626, 3646, 4079, 4079, 4079, 2827, 1943, 1959, 96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1301, 4063, 4063, 4063, 4063, 4063, 4063, 4079, 3887, 3067, 273, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1301, 4063, 4063, 4063, 4063, 4063, 4063, 4079, 4063, 4063, 1911, 321, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 883, 3806, 4063, 4063, 4063, 3308, 2778, 4079, 4063, 4063, 4063, 3003, 337, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3228, 4063, 4063, 4063, 2329, 514, 851, 3341, 4063, 4063, 4063, 1638, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 963, 3855, 4063, 4063, 4063, 4063, 3501, 867, 3357, 4063, 4063, 4063, 3196, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 417, 3148, 4063, 4063, 4063, 4063, 4063, 4096, 4063, 4063, 4063, 3903, 1574, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 401, 3164, 4063, 4063, 4063, 4063, 4096, 4063, 4063, 4063, 2762, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 369, 2056, 3871, 4063, 4063, 4096, 4063, 4063, 3196, 353, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 208, 1927, 3051, 2939, 3148, 1927, 305, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}; // 6
logic [BITS - 1 : 0] arr_0 [0 : WIDTH-1]= '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4096, 4016, 4096, 4016, 2256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2224, 3952, 4016, 3952, 4016, 3952, 4016, 3952, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2224, 4096, 4016, 4048, 4016, 4048, 4016, 4048, 4016, 4048, 4016, 4048, 368, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2224, 3952, 4016, 3952, 4016, 3952, 4016, 3952, 4016, 3952, 4016, 3952, 4016, 3952, 3120, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4096, 4016, 4096, 4016, 2256, 0, 1328, 1296, 4048, 4016, 4048, 4016, 4048, 4016, 4048, 4016, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1296, 4016, 3952, 4016, 3952, 4016, 0, 0, 0, 0, 0, 4016, 3952, 4016, 3952, 4016, 3952, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 432, 4016, 4096, 4016, 4096, 4016, 4048, 0, 0, 0, 0, 0, 4048, 4016, 4048, 4016, 4048, 4016, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4016, 3952, 4016, 3952, 4016, 3952, 2192, 0, 0, 0, 0, 0, 4016, 3952, 4016, 3952, 4016, 3952, 0, 0, 0, 0, 0, 0, 0, 0, 432, 4016, 4048, 4016, 4048, 4016, 4048, 4016, 0, 0, 0, 0, 0, 0, 4048, 4016, 4048, 4016, 4048, 2192, 0, 0, 0, 0, 0, 0, 0, 0, 4016, 3952, 4016, 3952, 4016, 3952, 2192, 0, 0, 0, 0, 0, 2224, 3952, 4016, 3952, 4016, 3952, 4016, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4096, 4016, 4048, 4016, 4048, 4016, 0, 0, 0, 0, 432, 4016, 4048, 4016, 4048, 4016, 4048, 4016, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4016, 3952, 4016, 3952, 4016, 3952, 0, 0, 0, 1296, 4016, 3952, 4016, 3952, 4016, 3952, 4016, 336, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4096, 4016, 4048, 4016, 4048, 4016, 0, 2224, 4048, 4016, 4048, 4016, 4048, 4016, 4048, 4016, 3152, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4016, 3952, 4016, 3952, 4016, 3952, 4016, 3952, 4016, 3952, 4016, 3952, 4016, 3952, 4016, 3952, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4096, 4016, 4048, 4016, 4048, 4016, 4048, 4016, 4048, 4016, 4048, 4016, 4048, 4016, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 368, 3952, 4016, 3952, 4016, 3952, 4016, 3952, 4016, 3952, 4016, 3952, 4016, 336, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3120, 4048, 4016, 4048, 4016, 4048, 4016, 4048, 4016, 3152, 1296, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4016, 3952, 4016, 3952, 4016, 3952, 4016, 3952, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1296, 1328, 3120, 1328, 1296, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0};
logic [BITS - 1 : 0] arr_2 [0 : WIDTH-1]= '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1872, 4048, 4096, 2544, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2192, 3952, 3120, 3120, 3856, 4048, 1360, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3952, 48, 0, 0, 0, 4048, 4048, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2256, 0, 0, 0, 0, 0, 3664, 2512, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3440, 3856, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3440, 3824, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3440, 3088, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3440, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3856, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1296, 3248, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2576, 1296, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 976, 1456, 3952, 4048, 3216, 848, 0, 4048, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3472, 3888, 1488, 1488, 2640, 3088, 4048, 3600, 4048, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2160, 3952, 0, 0, 0, 0, 0, 1136, 4048, 3088, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4048, 144, 0, 0, 0, 0, 0, 368, 4048, 4048, 3568, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2704, 4048, 0, 0, 0, 0, 0, 0, 3824, 0, 0, 3952, 4016, 368, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2992, 4048, 0, 0, 0, 0, 0, 1872, 2768, 0, 0, 0, 1456, 3984, 2384, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2160, 4048, 0, 0, 0, 0, 2448, 3344, 0, 0, 0, 0, 0, 0, 432, 1872, 1872, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3760, 3504, 1968, 3152, 4016, 3312, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2768, 4048, 4048, 1584, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0};

initial begin
    clk = 0;
    forever #5 clk = ~clk;  
end

initial begin
    reset_reg = 0;
    new_data = 0;
    #50;
    reset_reg = 1;
    #100;
    reset_reg = 0;
    #10;

    for (int j = 0; j < WIDTH; j++) begin
        #10;
        input_pixel = arr_2[j];
        new_data = 1;
        #12;
        new_data = 0;
        #20;   
    end

end
endmodule






// Good code
//(* ASYNC_REG = "TRUE"*) reg [6:0] sync;
//wire nn_en;

//// Enable for NN (toggle synchronizer)
//always @(posedge clk) begin
//    sync[6] <= sync[5];
//    sync[5] <= sync[4];
//    sync[4] <= sync[3];
//    sync[3] <= sync[2];
//    sync[2] <= sync[1];
//    sync[1] <= sync[0];
//    sync[0] <= new_data;
//end

//assign nn_en = ((~sync[2]) & sync[1]) | ((~sync[3]) & sync[2]) | ((~sync[4]) & sync[3]) | 
//               ((~sync[5]) & sync[4]) | ((~sync[6]) & sync[5]);
