`timescale 1ns / 1ps 
 
////////////////////////////////////////////////////////////////////////////////// 
// WEIGHT MEMORY (ROM) 
////////////////////////////////////////////////////////////////////////////////// 
module ROM_weights_0 #( 
    parameter int WGHT_INT = 6, // integer part 
    parameter int WGHT_FRC = 16 // fractional part 
)( 
    input logic clk, // clock 
    input logic [9:0] address,
    output [WGHT_INT + WGHT_FRC-1:0] dout 
); 

(* rom_style = "block" *) reg [WGHT_INT + WGHT_FRC-1:0] data;
generate 
  if (WGHT_FRC == 1) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 7'h00; 
        10'b0000000001: data <= 7'h00; 
        10'b0000000010: data <= 7'h00; 
        10'b0000000011: data <= 7'h00; 
        10'b0000000100: data <= 7'h00; 
        10'b0000000101: data <= 7'h00; 
        10'b0000000110: data <= 7'h00; 
        10'b0000000111: data <= 7'h00; 
        10'b0000001000: data <= 7'h00; 
        10'b0000001001: data <= 7'h00; 
        10'b0000001010: data <= 7'h00; 
        10'b0000001011: data <= 7'h00; 
        10'b0000001100: data <= 7'h00; 
        10'b0000001101: data <= 7'h00; 
        10'b0000001110: data <= 7'h00; 
        10'b0000001111: data <= 7'h00; 
        10'b0000010000: data <= 7'h00; 
        10'b0000010001: data <= 7'h00; 
        10'b0000010010: data <= 7'h00; 
        10'b0000010011: data <= 7'h00; 
        10'b0000010100: data <= 7'h00; 
        10'b0000010101: data <= 7'h00; 
        10'b0000010110: data <= 7'h00; 
        10'b0000010111: data <= 7'h00; 
        10'b0000011000: data <= 7'h00; 
        10'b0000011001: data <= 7'h00; 
        10'b0000011010: data <= 7'h00; 
        10'b0000011011: data <= 7'h00; 
        10'b0000011100: data <= 7'h00; 
        10'b0000011101: data <= 7'h00; 
        10'b0000011110: data <= 7'h00; 
        10'b0000011111: data <= 7'h00; 
        10'b0000100000: data <= 7'h00; 
        10'b0000100001: data <= 7'h00; 
        10'b0000100010: data <= 7'h00; 
        10'b0000100011: data <= 7'h00; 
        10'b0000100100: data <= 7'h00; 
        10'b0000100101: data <= 7'h00; 
        10'b0000100110: data <= 7'h00; 
        10'b0000100111: data <= 7'h00; 
        10'b0000101000: data <= 7'h00; 
        10'b0000101001: data <= 7'h00; 
        10'b0000101010: data <= 7'h00; 
        10'b0000101011: data <= 7'h00; 
        10'b0000101100: data <= 7'h00; 
        10'b0000101101: data <= 7'h00; 
        10'b0000101110: data <= 7'h00; 
        10'b0000101111: data <= 7'h00; 
        10'b0000110000: data <= 7'h00; 
        10'b0000110001: data <= 7'h00; 
        10'b0000110010: data <= 7'h00; 
        10'b0000110011: data <= 7'h00; 
        10'b0000110100: data <= 7'h00; 
        10'b0000110101: data <= 7'h00; 
        10'b0000110110: data <= 7'h00; 
        10'b0000110111: data <= 7'h00; 
        10'b0000111000: data <= 7'h00; 
        10'b0000111001: data <= 7'h00; 
        10'b0000111010: data <= 7'h00; 
        10'b0000111011: data <= 7'h00; 
        10'b0000111100: data <= 7'h00; 
        10'b0000111101: data <= 7'h00; 
        10'b0000111110: data <= 7'h00; 
        10'b0000111111: data <= 7'h00; 
        10'b0001000000: data <= 7'h00; 
        10'b0001000001: data <= 7'h00; 
        10'b0001000010: data <= 7'h00; 
        10'b0001000011: data <= 7'h00; 
        10'b0001000100: data <= 7'h00; 
        10'b0001000101: data <= 7'h00; 
        10'b0001000110: data <= 7'h00; 
        10'b0001000111: data <= 7'h00; 
        10'b0001001000: data <= 7'h00; 
        10'b0001001001: data <= 7'h00; 
        10'b0001001010: data <= 7'h00; 
        10'b0001001011: data <= 7'h00; 
        10'b0001001100: data <= 7'h00; 
        10'b0001001101: data <= 7'h00; 
        10'b0001001110: data <= 7'h00; 
        10'b0001001111: data <= 7'h00; 
        10'b0001010000: data <= 7'h00; 
        10'b0001010001: data <= 7'h00; 
        10'b0001010010: data <= 7'h00; 
        10'b0001010011: data <= 7'h00; 
        10'b0001010100: data <= 7'h00; 
        10'b0001010101: data <= 7'h00; 
        10'b0001010110: data <= 7'h00; 
        10'b0001010111: data <= 7'h00; 
        10'b0001011000: data <= 7'h00; 
        10'b0001011001: data <= 7'h00; 
        10'b0001011010: data <= 7'h00; 
        10'b0001011011: data <= 7'h00; 
        10'b0001011100: data <= 7'h00; 
        10'b0001011101: data <= 7'h00; 
        10'b0001011110: data <= 7'h00; 
        10'b0001011111: data <= 7'h00; 
        10'b0001100000: data <= 7'h00; 
        10'b0001100001: data <= 7'h00; 
        10'b0001100010: data <= 7'h00; 
        10'b0001100011: data <= 7'h00; 
        10'b0001100100: data <= 7'h00; 
        10'b0001100101: data <= 7'h00; 
        10'b0001100110: data <= 7'h00; 
        10'b0001100111: data <= 7'h00; 
        10'b0001101000: data <= 7'h00; 
        10'b0001101001: data <= 7'h00; 
        10'b0001101010: data <= 7'h00; 
        10'b0001101011: data <= 7'h00; 
        10'b0001101100: data <= 7'h00; 
        10'b0001101101: data <= 7'h00; 
        10'b0001101110: data <= 7'h00; 
        10'b0001101111: data <= 7'h00; 
        10'b0001110000: data <= 7'h00; 
        10'b0001110001: data <= 7'h00; 
        10'b0001110010: data <= 7'h00; 
        10'b0001110011: data <= 7'h00; 
        10'b0001110100: data <= 7'h00; 
        10'b0001110101: data <= 7'h00; 
        10'b0001110110: data <= 7'h00; 
        10'b0001110111: data <= 7'h00; 
        10'b0001111000: data <= 7'h00; 
        10'b0001111001: data <= 7'h00; 
        10'b0001111010: data <= 7'h00; 
        10'b0001111011: data <= 7'h00; 
        10'b0001111100: data <= 7'h00; 
        10'b0001111101: data <= 7'h00; 
        10'b0001111110: data <= 7'h00; 
        10'b0001111111: data <= 7'h00; 
        10'b0010000000: data <= 7'h00; 
        10'b0010000001: data <= 7'h00; 
        10'b0010000010: data <= 7'h00; 
        10'b0010000011: data <= 7'h00; 
        10'b0010000100: data <= 7'h00; 
        10'b0010000101: data <= 7'h00; 
        10'b0010000110: data <= 7'h00; 
        10'b0010000111: data <= 7'h00; 
        10'b0010001000: data <= 7'h00; 
        10'b0010001001: data <= 7'h00; 
        10'b0010001010: data <= 7'h00; 
        10'b0010001011: data <= 7'h00; 
        10'b0010001100: data <= 7'h00; 
        10'b0010001101: data <= 7'h00; 
        10'b0010001110: data <= 7'h00; 
        10'b0010001111: data <= 7'h00; 
        10'b0010010000: data <= 7'h00; 
        10'b0010010001: data <= 7'h00; 
        10'b0010010010: data <= 7'h00; 
        10'b0010010011: data <= 7'h00; 
        10'b0010010100: data <= 7'h00; 
        10'b0010010101: data <= 7'h00; 
        10'b0010010110: data <= 7'h00; 
        10'b0010010111: data <= 7'h00; 
        10'b0010011000: data <= 7'h00; 
        10'b0010011001: data <= 7'h00; 
        10'b0010011010: data <= 7'h00; 
        10'b0010011011: data <= 7'h00; 
        10'b0010011100: data <= 7'h00; 
        10'b0010011101: data <= 7'h00; 
        10'b0010011110: data <= 7'h00; 
        10'b0010011111: data <= 7'h00; 
        10'b0010100000: data <= 7'h00; 
        10'b0010100001: data <= 7'h00; 
        10'b0010100010: data <= 7'h00; 
        10'b0010100011: data <= 7'h00; 
        10'b0010100100: data <= 7'h00; 
        10'b0010100101: data <= 7'h00; 
        10'b0010100110: data <= 7'h00; 
        10'b0010100111: data <= 7'h00; 
        10'b0010101000: data <= 7'h00; 
        10'b0010101001: data <= 7'h00; 
        10'b0010101010: data <= 7'h00; 
        10'b0010101011: data <= 7'h00; 
        10'b0010101100: data <= 7'h00; 
        10'b0010101101: data <= 7'h00; 
        10'b0010101110: data <= 7'h00; 
        10'b0010101111: data <= 7'h00; 
        10'b0010110000: data <= 7'h00; 
        10'b0010110001: data <= 7'h00; 
        10'b0010110010: data <= 7'h00; 
        10'b0010110011: data <= 7'h00; 
        10'b0010110100: data <= 7'h00; 
        10'b0010110101: data <= 7'h00; 
        10'b0010110110: data <= 7'h00; 
        10'b0010110111: data <= 7'h00; 
        10'b0010111000: data <= 7'h00; 
        10'b0010111001: data <= 7'h00; 
        10'b0010111010: data <= 7'h00; 
        10'b0010111011: data <= 7'h00; 
        10'b0010111100: data <= 7'h00; 
        10'b0010111101: data <= 7'h00; 
        10'b0010111110: data <= 7'h00; 
        10'b0010111111: data <= 7'h00; 
        10'b0011000000: data <= 7'h00; 
        10'b0011000001: data <= 7'h00; 
        10'b0011000010: data <= 7'h00; 
        10'b0011000011: data <= 7'h00; 
        10'b0011000100: data <= 7'h00; 
        10'b0011000101: data <= 7'h00; 
        10'b0011000110: data <= 7'h00; 
        10'b0011000111: data <= 7'h00; 
        10'b0011001000: data <= 7'h00; 
        10'b0011001001: data <= 7'h00; 
        10'b0011001010: data <= 7'h00; 
        10'b0011001011: data <= 7'h00; 
        10'b0011001100: data <= 7'h00; 
        10'b0011001101: data <= 7'h00; 
        10'b0011001110: data <= 7'h00; 
        10'b0011001111: data <= 7'h00; 
        10'b0011010000: data <= 7'h00; 
        10'b0011010001: data <= 7'h00; 
        10'b0011010010: data <= 7'h00; 
        10'b0011010011: data <= 7'h00; 
        10'b0011010100: data <= 7'h00; 
        10'b0011010101: data <= 7'h00; 
        10'b0011010110: data <= 7'h00; 
        10'b0011010111: data <= 7'h00; 
        10'b0011011000: data <= 7'h00; 
        10'b0011011001: data <= 7'h00; 
        10'b0011011010: data <= 7'h00; 
        10'b0011011011: data <= 7'h00; 
        10'b0011011100: data <= 7'h00; 
        10'b0011011101: data <= 7'h00; 
        10'b0011011110: data <= 7'h00; 
        10'b0011011111: data <= 7'h00; 
        10'b0011100000: data <= 7'h00; 
        10'b0011100001: data <= 7'h00; 
        10'b0011100010: data <= 7'h00; 
        10'b0011100011: data <= 7'h00; 
        10'b0011100100: data <= 7'h00; 
        10'b0011100101: data <= 7'h00; 
        10'b0011100110: data <= 7'h00; 
        10'b0011100111: data <= 7'h00; 
        10'b0011101000: data <= 7'h00; 
        10'b0011101001: data <= 7'h00; 
        10'b0011101010: data <= 7'h00; 
        10'b0011101011: data <= 7'h00; 
        10'b0011101100: data <= 7'h00; 
        10'b0011101101: data <= 7'h00; 
        10'b0011101110: data <= 7'h00; 
        10'b0011101111: data <= 7'h00; 
        10'b0011110000: data <= 7'h01; 
        10'b0011110001: data <= 7'h01; 
        10'b0011110010: data <= 7'h00; 
        10'b0011110011: data <= 7'h00; 
        10'b0011110100: data <= 7'h00; 
        10'b0011110101: data <= 7'h00; 
        10'b0011110110: data <= 7'h00; 
        10'b0011110111: data <= 7'h00; 
        10'b0011111000: data <= 7'h00; 
        10'b0011111001: data <= 7'h00; 
        10'b0011111010: data <= 7'h00; 
        10'b0011111011: data <= 7'h00; 
        10'b0011111100: data <= 7'h00; 
        10'b0011111101: data <= 7'h00; 
        10'b0011111110: data <= 7'h00; 
        10'b0011111111: data <= 7'h00; 
        10'b0100000000: data <= 7'h00; 
        10'b0100000001: data <= 7'h00; 
        10'b0100000010: data <= 7'h00; 
        10'b0100000011: data <= 7'h00; 
        10'b0100000100: data <= 7'h00; 
        10'b0100000101: data <= 7'h00; 
        10'b0100000110: data <= 7'h00; 
        10'b0100000111: data <= 7'h00; 
        10'b0100001000: data <= 7'h00; 
        10'b0100001001: data <= 7'h00; 
        10'b0100001010: data <= 7'h00; 
        10'b0100001011: data <= 7'h00; 
        10'b0100001100: data <= 7'h00; 
        10'b0100001101: data <= 7'h00; 
        10'b0100001110: data <= 7'h01; 
        10'b0100001111: data <= 7'h00; 
        10'b0100010000: data <= 7'h00; 
        10'b0100010001: data <= 7'h00; 
        10'b0100010010: data <= 7'h00; 
        10'b0100010011: data <= 7'h01; 
        10'b0100010100: data <= 7'h00; 
        10'b0100010101: data <= 7'h00; 
        10'b0100010110: data <= 7'h00; 
        10'b0100010111: data <= 7'h00; 
        10'b0100011000: data <= 7'h00; 
        10'b0100011001: data <= 7'h00; 
        10'b0100011010: data <= 7'h00; 
        10'b0100011011: data <= 7'h00; 
        10'b0100011100: data <= 7'h00; 
        10'b0100011101: data <= 7'h00; 
        10'b0100011110: data <= 7'h00; 
        10'b0100011111: data <= 7'h00; 
        10'b0100100000: data <= 7'h00; 
        10'b0100100001: data <= 7'h00; 
        10'b0100100010: data <= 7'h00; 
        10'b0100100011: data <= 7'h00; 
        10'b0100100100: data <= 7'h00; 
        10'b0100100101: data <= 7'h00; 
        10'b0100100110: data <= 7'h00; 
        10'b0100100111: data <= 7'h00; 
        10'b0100101000: data <= 7'h00; 
        10'b0100101001: data <= 7'h00; 
        10'b0100101010: data <= 7'h00; 
        10'b0100101011: data <= 7'h00; 
        10'b0100101100: data <= 7'h00; 
        10'b0100101101: data <= 7'h00; 
        10'b0100101110: data <= 7'h00; 
        10'b0100101111: data <= 7'h01; 
        10'b0100110000: data <= 7'h00; 
        10'b0100110001: data <= 7'h00; 
        10'b0100110010: data <= 7'h00; 
        10'b0100110011: data <= 7'h00; 
        10'b0100110100: data <= 7'h00; 
        10'b0100110101: data <= 7'h00; 
        10'b0100110110: data <= 7'h00; 
        10'b0100110111: data <= 7'h00; 
        10'b0100111000: data <= 7'h00; 
        10'b0100111001: data <= 7'h00; 
        10'b0100111010: data <= 7'h00; 
        10'b0100111011: data <= 7'h00; 
        10'b0100111100: data <= 7'h00; 
        10'b0100111101: data <= 7'h00; 
        10'b0100111110: data <= 7'h00; 
        10'b0100111111: data <= 7'h00; 
        10'b0101000000: data <= 7'h00; 
        10'b0101000001: data <= 7'h00; 
        10'b0101000010: data <= 7'h00; 
        10'b0101000011: data <= 7'h7f; 
        10'b0101000100: data <= 7'h7f; 
        10'b0101000101: data <= 7'h00; 
        10'b0101000110: data <= 7'h00; 
        10'b0101000111: data <= 7'h00; 
        10'b0101001000: data <= 7'h00; 
        10'b0101001001: data <= 7'h00; 
        10'b0101001010: data <= 7'h00; 
        10'b0101001011: data <= 7'h01; 
        10'b0101001100: data <= 7'h00; 
        10'b0101001101: data <= 7'h00; 
        10'b0101001110: data <= 7'h00; 
        10'b0101001111: data <= 7'h00; 
        10'b0101010000: data <= 7'h00; 
        10'b0101010001: data <= 7'h00; 
        10'b0101010010: data <= 7'h00; 
        10'b0101010011: data <= 7'h00; 
        10'b0101010100: data <= 7'h00; 
        10'b0101010101: data <= 7'h00; 
        10'b0101010110: data <= 7'h00; 
        10'b0101010111: data <= 7'h00; 
        10'b0101011000: data <= 7'h00; 
        10'b0101011001: data <= 7'h00; 
        10'b0101011010: data <= 7'h00; 
        10'b0101011011: data <= 7'h00; 
        10'b0101011100: data <= 7'h00; 
        10'b0101011101: data <= 7'h00; 
        10'b0101011110: data <= 7'h7f; 
        10'b0101011111: data <= 7'h7f; 
        10'b0101100000: data <= 7'h7f; 
        10'b0101100001: data <= 7'h7f; 
        10'b0101100010: data <= 7'h00; 
        10'b0101100011: data <= 7'h00; 
        10'b0101100100: data <= 7'h00; 
        10'b0101100101: data <= 7'h00; 
        10'b0101100110: data <= 7'h01; 
        10'b0101100111: data <= 7'h01; 
        10'b0101101000: data <= 7'h00; 
        10'b0101101001: data <= 7'h00; 
        10'b0101101010: data <= 7'h00; 
        10'b0101101011: data <= 7'h00; 
        10'b0101101100: data <= 7'h00; 
        10'b0101101101: data <= 7'h00; 
        10'b0101101110: data <= 7'h00; 
        10'b0101101111: data <= 7'h00; 
        10'b0101110000: data <= 7'h00; 
        10'b0101110001: data <= 7'h00; 
        10'b0101110010: data <= 7'h00; 
        10'b0101110011: data <= 7'h00; 
        10'b0101110100: data <= 7'h00; 
        10'b0101110101: data <= 7'h00; 
        10'b0101110110: data <= 7'h00; 
        10'b0101110111: data <= 7'h00; 
        10'b0101111000: data <= 7'h00; 
        10'b0101111001: data <= 7'h7f; 
        10'b0101111010: data <= 7'h7f; 
        10'b0101111011: data <= 7'h7f; 
        10'b0101111100: data <= 7'h7f; 
        10'b0101111101: data <= 7'h00; 
        10'b0101111110: data <= 7'h00; 
        10'b0101111111: data <= 7'h00; 
        10'b0110000000: data <= 7'h00; 
        10'b0110000001: data <= 7'h00; 
        10'b0110000010: data <= 7'h00; 
        10'b0110000011: data <= 7'h01; 
        10'b0110000100: data <= 7'h00; 
        10'b0110000101: data <= 7'h00; 
        10'b0110000110: data <= 7'h00; 
        10'b0110000111: data <= 7'h00; 
        10'b0110001000: data <= 7'h00; 
        10'b0110001001: data <= 7'h00; 
        10'b0110001010: data <= 7'h00; 
        10'b0110001011: data <= 7'h00; 
        10'b0110001100: data <= 7'h00; 
        10'b0110001101: data <= 7'h00; 
        10'b0110001110: data <= 7'h00; 
        10'b0110001111: data <= 7'h00; 
        10'b0110010000: data <= 7'h00; 
        10'b0110010001: data <= 7'h00; 
        10'b0110010010: data <= 7'h00; 
        10'b0110010011: data <= 7'h00; 
        10'b0110010100: data <= 7'h00; 
        10'b0110010101: data <= 7'h00; 
        10'b0110010110: data <= 7'h7f; 
        10'b0110010111: data <= 7'h7f; 
        10'b0110011000: data <= 7'h7f; 
        10'b0110011001: data <= 7'h7f; 
        10'b0110011010: data <= 7'h00; 
        10'b0110011011: data <= 7'h00; 
        10'b0110011100: data <= 7'h00; 
        10'b0110011101: data <= 7'h00; 
        10'b0110011110: data <= 7'h00; 
        10'b0110011111: data <= 7'h01; 
        10'b0110100000: data <= 7'h00; 
        10'b0110100001: data <= 7'h00; 
        10'b0110100010: data <= 7'h00; 
        10'b0110100011: data <= 7'h00; 
        10'b0110100100: data <= 7'h00; 
        10'b0110100101: data <= 7'h00; 
        10'b0110100110: data <= 7'h00; 
        10'b0110100111: data <= 7'h00; 
        10'b0110101000: data <= 7'h00; 
        10'b0110101001: data <= 7'h00; 
        10'b0110101010: data <= 7'h00; 
        10'b0110101011: data <= 7'h00; 
        10'b0110101100: data <= 7'h00; 
        10'b0110101101: data <= 7'h00; 
        10'b0110101110: data <= 7'h00; 
        10'b0110101111: data <= 7'h00; 
        10'b0110110000: data <= 7'h00; 
        10'b0110110001: data <= 7'h7f; 
        10'b0110110010: data <= 7'h7f; 
        10'b0110110011: data <= 7'h7f; 
        10'b0110110100: data <= 7'h7f; 
        10'b0110110101: data <= 7'h00; 
        10'b0110110110: data <= 7'h00; 
        10'b0110110111: data <= 7'h00; 
        10'b0110111000: data <= 7'h00; 
        10'b0110111001: data <= 7'h00; 
        10'b0110111010: data <= 7'h00; 
        10'b0110111011: data <= 7'h00; 
        10'b0110111100: data <= 7'h00; 
        10'b0110111101: data <= 7'h00; 
        10'b0110111110: data <= 7'h00; 
        10'b0110111111: data <= 7'h00; 
        10'b0111000000: data <= 7'h00; 
        10'b0111000001: data <= 7'h00; 
        10'b0111000010: data <= 7'h00; 
        10'b0111000011: data <= 7'h00; 
        10'b0111000100: data <= 7'h00; 
        10'b0111000101: data <= 7'h00; 
        10'b0111000110: data <= 7'h00; 
        10'b0111000111: data <= 7'h00; 
        10'b0111001000: data <= 7'h00; 
        10'b0111001001: data <= 7'h00; 
        10'b0111001010: data <= 7'h00; 
        10'b0111001011: data <= 7'h00; 
        10'b0111001100: data <= 7'h7f; 
        10'b0111001101: data <= 7'h7f; 
        10'b0111001110: data <= 7'h7f; 
        10'b0111001111: data <= 7'h7f; 
        10'b0111010000: data <= 7'h00; 
        10'b0111010001: data <= 7'h00; 
        10'b0111010010: data <= 7'h00; 
        10'b0111010011: data <= 7'h00; 
        10'b0111010100: data <= 7'h00; 
        10'b0111010101: data <= 7'h00; 
        10'b0111010110: data <= 7'h00; 
        10'b0111010111: data <= 7'h00; 
        10'b0111011000: data <= 7'h00; 
        10'b0111011001: data <= 7'h00; 
        10'b0111011010: data <= 7'h00; 
        10'b0111011011: data <= 7'h00; 
        10'b0111011100: data <= 7'h00; 
        10'b0111011101: data <= 7'h00; 
        10'b0111011110: data <= 7'h00; 
        10'b0111011111: data <= 7'h00; 
        10'b0111100000: data <= 7'h00; 
        10'b0111100001: data <= 7'h00; 
        10'b0111100010: data <= 7'h00; 
        10'b0111100011: data <= 7'h00; 
        10'b0111100100: data <= 7'h00; 
        10'b0111100101: data <= 7'h00; 
        10'b0111100110: data <= 7'h00; 
        10'b0111100111: data <= 7'h00; 
        10'b0111101000: data <= 7'h7f; 
        10'b0111101001: data <= 7'h7f; 
        10'b0111101010: data <= 7'h7f; 
        10'b0111101011: data <= 7'h7f; 
        10'b0111101100: data <= 7'h00; 
        10'b0111101101: data <= 7'h00; 
        10'b0111101110: data <= 7'h00; 
        10'b0111101111: data <= 7'h00; 
        10'b0111110000: data <= 7'h00; 
        10'b0111110001: data <= 7'h00; 
        10'b0111110010: data <= 7'h00; 
        10'b0111110011: data <= 7'h00; 
        10'b0111110100: data <= 7'h00; 
        10'b0111110101: data <= 7'h00; 
        10'b0111110110: data <= 7'h00; 
        10'b0111110111: data <= 7'h00; 
        10'b0111111000: data <= 7'h00; 
        10'b0111111001: data <= 7'h00; 
        10'b0111111010: data <= 7'h00; 
        10'b0111111011: data <= 7'h00; 
        10'b0111111100: data <= 7'h00; 
        10'b0111111101: data <= 7'h00; 
        10'b0111111110: data <= 7'h00; 
        10'b0111111111: data <= 7'h00; 
        10'b1000000000: data <= 7'h00; 
        10'b1000000001: data <= 7'h00; 
        10'b1000000010: data <= 7'h01; 
        10'b1000000011: data <= 7'h00; 
        10'b1000000100: data <= 7'h7f; 
        10'b1000000101: data <= 7'h7f; 
        10'b1000000110: data <= 7'h7f; 
        10'b1000000111: data <= 7'h00; 
        10'b1000001000: data <= 7'h00; 
        10'b1000001001: data <= 7'h00; 
        10'b1000001010: data <= 7'h00; 
        10'b1000001011: data <= 7'h00; 
        10'b1000001100: data <= 7'h00; 
        10'b1000001101: data <= 7'h00; 
        10'b1000001110: data <= 7'h00; 
        10'b1000001111: data <= 7'h00; 
        10'b1000010000: data <= 7'h00; 
        10'b1000010001: data <= 7'h00; 
        10'b1000010010: data <= 7'h00; 
        10'b1000010011: data <= 7'h00; 
        10'b1000010100: data <= 7'h00; 
        10'b1000010101: data <= 7'h00; 
        10'b1000010110: data <= 7'h00; 
        10'b1000010111: data <= 7'h00; 
        10'b1000011000: data <= 7'h00; 
        10'b1000011001: data <= 7'h00; 
        10'b1000011010: data <= 7'h00; 
        10'b1000011011: data <= 7'h00; 
        10'b1000011100: data <= 7'h00; 
        10'b1000011101: data <= 7'h00; 
        10'b1000011110: data <= 7'h01; 
        10'b1000011111: data <= 7'h00; 
        10'b1000100000: data <= 7'h00; 
        10'b1000100001: data <= 7'h00; 
        10'b1000100010: data <= 7'h00; 
        10'b1000100011: data <= 7'h00; 
        10'b1000100100: data <= 7'h00; 
        10'b1000100101: data <= 7'h00; 
        10'b1000100110: data <= 7'h00; 
        10'b1000100111: data <= 7'h00; 
        10'b1000101000: data <= 7'h00; 
        10'b1000101001: data <= 7'h00; 
        10'b1000101010: data <= 7'h00; 
        10'b1000101011: data <= 7'h00; 
        10'b1000101100: data <= 7'h00; 
        10'b1000101101: data <= 7'h00; 
        10'b1000101110: data <= 7'h00; 
        10'b1000101111: data <= 7'h00; 
        10'b1000110000: data <= 7'h00; 
        10'b1000110001: data <= 7'h00; 
        10'b1000110010: data <= 7'h00; 
        10'b1000110011: data <= 7'h00; 
        10'b1000110100: data <= 7'h00; 
        10'b1000110101: data <= 7'h00; 
        10'b1000110110: data <= 7'h00; 
        10'b1000110111: data <= 7'h00; 
        10'b1000111000: data <= 7'h00; 
        10'b1000111001: data <= 7'h00; 
        10'b1000111010: data <= 7'h01; 
        10'b1000111011: data <= 7'h01; 
        10'b1000111100: data <= 7'h00; 
        10'b1000111101: data <= 7'h00; 
        10'b1000111110: data <= 7'h00; 
        10'b1000111111: data <= 7'h00; 
        10'b1001000000: data <= 7'h00; 
        10'b1001000001: data <= 7'h00; 
        10'b1001000010: data <= 7'h00; 
        10'b1001000011: data <= 7'h00; 
        10'b1001000100: data <= 7'h00; 
        10'b1001000101: data <= 7'h00; 
        10'b1001000110: data <= 7'h00; 
        10'b1001000111: data <= 7'h00; 
        10'b1001001000: data <= 7'h00; 
        10'b1001001001: data <= 7'h00; 
        10'b1001001010: data <= 7'h00; 
        10'b1001001011: data <= 7'h00; 
        10'b1001001100: data <= 7'h00; 
        10'b1001001101: data <= 7'h00; 
        10'b1001001110: data <= 7'h00; 
        10'b1001001111: data <= 7'h00; 
        10'b1001010000: data <= 7'h00; 
        10'b1001010001: data <= 7'h00; 
        10'b1001010010: data <= 7'h00; 
        10'b1001010011: data <= 7'h00; 
        10'b1001010100: data <= 7'h00; 
        10'b1001010101: data <= 7'h00; 
        10'b1001010110: data <= 7'h01; 
        10'b1001010111: data <= 7'h01; 
        10'b1001011000: data <= 7'h00; 
        10'b1001011001: data <= 7'h00; 
        10'b1001011010: data <= 7'h00; 
        10'b1001011011: data <= 7'h00; 
        10'b1001011100: data <= 7'h00; 
        10'b1001011101: data <= 7'h00; 
        10'b1001011110: data <= 7'h00; 
        10'b1001011111: data <= 7'h00; 
        10'b1001100000: data <= 7'h00; 
        10'b1001100001: data <= 7'h00; 
        10'b1001100010: data <= 7'h00; 
        10'b1001100011: data <= 7'h00; 
        10'b1001100100: data <= 7'h00; 
        10'b1001100101: data <= 7'h00; 
        10'b1001100110: data <= 7'h00; 
        10'b1001100111: data <= 7'h00; 
        10'b1001101000: data <= 7'h00; 
        10'b1001101001: data <= 7'h00; 
        10'b1001101010: data <= 7'h00; 
        10'b1001101011: data <= 7'h00; 
        10'b1001101100: data <= 7'h00; 
        10'b1001101101: data <= 7'h00; 
        10'b1001101110: data <= 7'h00; 
        10'b1001101111: data <= 7'h00; 
        10'b1001110000: data <= 7'h00; 
        10'b1001110001: data <= 7'h00; 
        10'b1001110010: data <= 7'h00; 
        10'b1001110011: data <= 7'h00; 
        10'b1001110100: data <= 7'h00; 
        10'b1001110101: data <= 7'h00; 
        10'b1001110110: data <= 7'h00; 
        10'b1001110111: data <= 7'h00; 
        10'b1001111000: data <= 7'h00; 
        10'b1001111001: data <= 7'h00; 
        10'b1001111010: data <= 7'h00; 
        10'b1001111011: data <= 7'h00; 
        10'b1001111100: data <= 7'h00; 
        10'b1001111101: data <= 7'h00; 
        10'b1001111110: data <= 7'h00; 
        10'b1001111111: data <= 7'h00; 
        10'b1010000000: data <= 7'h00; 
        10'b1010000001: data <= 7'h00; 
        10'b1010000010: data <= 7'h00; 
        10'b1010000011: data <= 7'h00; 
        10'b1010000100: data <= 7'h00; 
        10'b1010000101: data <= 7'h00; 
        10'b1010000110: data <= 7'h00; 
        10'b1010000111: data <= 7'h00; 
        10'b1010001000: data <= 7'h00; 
        10'b1010001001: data <= 7'h00; 
        10'b1010001010: data <= 7'h00; 
        10'b1010001011: data <= 7'h00; 
        10'b1010001100: data <= 7'h00; 
        10'b1010001101: data <= 7'h00; 
        10'b1010001110: data <= 7'h00; 
        10'b1010001111: data <= 7'h01; 
        10'b1010010000: data <= 7'h01; 
        10'b1010010001: data <= 7'h00; 
        10'b1010010010: data <= 7'h00; 
        10'b1010010011: data <= 7'h00; 
        10'b1010010100: data <= 7'h00; 
        10'b1010010101: data <= 7'h00; 
        10'b1010010110: data <= 7'h00; 
        10'b1010010111: data <= 7'h00; 
        10'b1010011000: data <= 7'h00; 
        10'b1010011001: data <= 7'h00; 
        10'b1010011010: data <= 7'h00; 
        10'b1010011011: data <= 7'h00; 
        10'b1010011100: data <= 7'h00; 
        10'b1010011101: data <= 7'h00; 
        10'b1010011110: data <= 7'h00; 
        10'b1010011111: data <= 7'h00; 
        10'b1010100000: data <= 7'h00; 
        10'b1010100001: data <= 7'h00; 
        10'b1010100010: data <= 7'h00; 
        10'b1010100011: data <= 7'h00; 
        10'b1010100100: data <= 7'h00; 
        10'b1010100101: data <= 7'h00; 
        10'b1010100110: data <= 7'h00; 
        10'b1010100111: data <= 7'h00; 
        10'b1010101000: data <= 7'h00; 
        10'b1010101001: data <= 7'h00; 
        10'b1010101010: data <= 7'h00; 
        10'b1010101011: data <= 7'h00; 
        10'b1010101100: data <= 7'h00; 
        10'b1010101101: data <= 7'h00; 
        10'b1010101110: data <= 7'h00; 
        10'b1010101111: data <= 7'h00; 
        10'b1010110000: data <= 7'h00; 
        10'b1010110001: data <= 7'h00; 
        10'b1010110010: data <= 7'h00; 
        10'b1010110011: data <= 7'h00; 
        10'b1010110100: data <= 7'h00; 
        10'b1010110101: data <= 7'h00; 
        10'b1010110110: data <= 7'h00; 
        10'b1010110111: data <= 7'h00; 
        10'b1010111000: data <= 7'h00; 
        10'b1010111001: data <= 7'h00; 
        10'b1010111010: data <= 7'h00; 
        10'b1010111011: data <= 7'h00; 
        10'b1010111100: data <= 7'h00; 
        10'b1010111101: data <= 7'h00; 
        10'b1010111110: data <= 7'h00; 
        10'b1010111111: data <= 7'h00; 
        10'b1011000000: data <= 7'h00; 
        10'b1011000001: data <= 7'h00; 
        10'b1011000010: data <= 7'h00; 
        10'b1011000011: data <= 7'h00; 
        10'b1011000100: data <= 7'h00; 
        10'b1011000101: data <= 7'h00; 
        10'b1011000110: data <= 7'h00; 
        10'b1011000111: data <= 7'h00; 
        10'b1011001000: data <= 7'h00; 
        10'b1011001001: data <= 7'h00; 
        10'b1011001010: data <= 7'h00; 
        10'b1011001011: data <= 7'h00; 
        10'b1011001100: data <= 7'h00; 
        10'b1011001101: data <= 7'h00; 
        10'b1011001110: data <= 7'h00; 
        10'b1011001111: data <= 7'h00; 
        10'b1011010000: data <= 7'h00; 
        10'b1011010001: data <= 7'h00; 
        10'b1011010010: data <= 7'h00; 
        10'b1011010011: data <= 7'h00; 
        10'b1011010100: data <= 7'h00; 
        10'b1011010101: data <= 7'h00; 
        10'b1011010110: data <= 7'h00; 
        10'b1011010111: data <= 7'h00; 
        10'b1011011000: data <= 7'h00; 
        10'b1011011001: data <= 7'h00; 
        10'b1011011010: data <= 7'h00; 
        10'b1011011011: data <= 7'h00; 
        10'b1011011100: data <= 7'h00; 
        10'b1011011101: data <= 7'h00; 
        10'b1011011110: data <= 7'h00; 
        10'b1011011111: data <= 7'h00; 
        10'b1011100000: data <= 7'h00; 
        10'b1011100001: data <= 7'h00; 
        10'b1011100010: data <= 7'h00; 
        10'b1011100011: data <= 7'h00; 
        10'b1011100100: data <= 7'h00; 
        10'b1011100101: data <= 7'h00; 
        10'b1011100110: data <= 7'h00; 
        10'b1011100111: data <= 7'h00; 
        10'b1011101000: data <= 7'h00; 
        10'b1011101001: data <= 7'h00; 
        10'b1011101010: data <= 7'h00; 
        10'b1011101011: data <= 7'h00; 
        10'b1011101100: data <= 7'h00; 
        10'b1011101101: data <= 7'h00; 
        10'b1011101110: data <= 7'h00; 
        10'b1011101111: data <= 7'h00; 
        10'b1011110000: data <= 7'h00; 
        10'b1011110001: data <= 7'h00; 
        10'b1011110010: data <= 7'h00; 
        10'b1011110011: data <= 7'h00; 
        10'b1011110100: data <= 7'h00; 
        10'b1011110101: data <= 7'h00; 
        10'b1011110110: data <= 7'h00; 
        10'b1011110111: data <= 7'h00; 
        10'b1011111000: data <= 7'h00; 
        10'b1011111001: data <= 7'h00; 
        10'b1011111010: data <= 7'h00; 
        10'b1011111011: data <= 7'h00; 
        10'b1011111100: data <= 7'h00; 
        10'b1011111101: data <= 7'h00; 
        10'b1011111110: data <= 7'h00; 
        10'b1011111111: data <= 7'h00; 
        10'b1100000000: data <= 7'h00; 
        10'b1100000001: data <= 7'h00; 
        10'b1100000010: data <= 7'h00; 
        10'b1100000011: data <= 7'h00; 
        10'b1100000100: data <= 7'h00; 
        10'b1100000101: data <= 7'h00; 
        10'b1100000110: data <= 7'h00; 
        10'b1100000111: data <= 7'h00; 
        10'b1100001000: data <= 7'h00; 
        10'b1100001001: data <= 7'h00; 
        10'b1100001010: data <= 7'h00; 
        10'b1100001011: data <= 7'h00; 
        10'b1100001100: data <= 7'h00; 
        10'b1100001101: data <= 7'h00; 
        10'b1100001110: data <= 7'h00; 
        10'b1100001111: data <= 7'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 2) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 8'h00; 
        10'b0000000001: data <= 8'h00; 
        10'b0000000010: data <= 8'h00; 
        10'b0000000011: data <= 8'h00; 
        10'b0000000100: data <= 8'h00; 
        10'b0000000101: data <= 8'h00; 
        10'b0000000110: data <= 8'h00; 
        10'b0000000111: data <= 8'h00; 
        10'b0000001000: data <= 8'h00; 
        10'b0000001001: data <= 8'h00; 
        10'b0000001010: data <= 8'h00; 
        10'b0000001011: data <= 8'h00; 
        10'b0000001100: data <= 8'h00; 
        10'b0000001101: data <= 8'h00; 
        10'b0000001110: data <= 8'h00; 
        10'b0000001111: data <= 8'h00; 
        10'b0000010000: data <= 8'h00; 
        10'b0000010001: data <= 8'h00; 
        10'b0000010010: data <= 8'h00; 
        10'b0000010011: data <= 8'h00; 
        10'b0000010100: data <= 8'h00; 
        10'b0000010101: data <= 8'h00; 
        10'b0000010110: data <= 8'h00; 
        10'b0000010111: data <= 8'h00; 
        10'b0000011000: data <= 8'h00; 
        10'b0000011001: data <= 8'h00; 
        10'b0000011010: data <= 8'h00; 
        10'b0000011011: data <= 8'h00; 
        10'b0000011100: data <= 8'h00; 
        10'b0000011101: data <= 8'h00; 
        10'b0000011110: data <= 8'h00; 
        10'b0000011111: data <= 8'h00; 
        10'b0000100000: data <= 8'h00; 
        10'b0000100001: data <= 8'h00; 
        10'b0000100010: data <= 8'h00; 
        10'b0000100011: data <= 8'h00; 
        10'b0000100100: data <= 8'h00; 
        10'b0000100101: data <= 8'h00; 
        10'b0000100110: data <= 8'h00; 
        10'b0000100111: data <= 8'h00; 
        10'b0000101000: data <= 8'h00; 
        10'b0000101001: data <= 8'h00; 
        10'b0000101010: data <= 8'h00; 
        10'b0000101011: data <= 8'h00; 
        10'b0000101100: data <= 8'h00; 
        10'b0000101101: data <= 8'h00; 
        10'b0000101110: data <= 8'h00; 
        10'b0000101111: data <= 8'h00; 
        10'b0000110000: data <= 8'h00; 
        10'b0000110001: data <= 8'h00; 
        10'b0000110010: data <= 8'h00; 
        10'b0000110011: data <= 8'h00; 
        10'b0000110100: data <= 8'h00; 
        10'b0000110101: data <= 8'h00; 
        10'b0000110110: data <= 8'h00; 
        10'b0000110111: data <= 8'h00; 
        10'b0000111000: data <= 8'h00; 
        10'b0000111001: data <= 8'h00; 
        10'b0000111010: data <= 8'h00; 
        10'b0000111011: data <= 8'h00; 
        10'b0000111100: data <= 8'h00; 
        10'b0000111101: data <= 8'h00; 
        10'b0000111110: data <= 8'h00; 
        10'b0000111111: data <= 8'h00; 
        10'b0001000000: data <= 8'h00; 
        10'b0001000001: data <= 8'h00; 
        10'b0001000010: data <= 8'h00; 
        10'b0001000011: data <= 8'h00; 
        10'b0001000100: data <= 8'h00; 
        10'b0001000101: data <= 8'h00; 
        10'b0001000110: data <= 8'h00; 
        10'b0001000111: data <= 8'h00; 
        10'b0001001000: data <= 8'h00; 
        10'b0001001001: data <= 8'h00; 
        10'b0001001010: data <= 8'h00; 
        10'b0001001011: data <= 8'h00; 
        10'b0001001100: data <= 8'h00; 
        10'b0001001101: data <= 8'h00; 
        10'b0001001110: data <= 8'h00; 
        10'b0001001111: data <= 8'h00; 
        10'b0001010000: data <= 8'h00; 
        10'b0001010001: data <= 8'h00; 
        10'b0001010010: data <= 8'h00; 
        10'b0001010011: data <= 8'h00; 
        10'b0001010100: data <= 8'h00; 
        10'b0001010101: data <= 8'h00; 
        10'b0001010110: data <= 8'h00; 
        10'b0001010111: data <= 8'h00; 
        10'b0001011000: data <= 8'h00; 
        10'b0001011001: data <= 8'h00; 
        10'b0001011010: data <= 8'h00; 
        10'b0001011011: data <= 8'h00; 
        10'b0001011100: data <= 8'h00; 
        10'b0001011101: data <= 8'h00; 
        10'b0001011110: data <= 8'h00; 
        10'b0001011111: data <= 8'h00; 
        10'b0001100000: data <= 8'h00; 
        10'b0001100001: data <= 8'h00; 
        10'b0001100010: data <= 8'h00; 
        10'b0001100011: data <= 8'h00; 
        10'b0001100100: data <= 8'h00; 
        10'b0001100101: data <= 8'h00; 
        10'b0001100110: data <= 8'h00; 
        10'b0001100111: data <= 8'h00; 
        10'b0001101000: data <= 8'h00; 
        10'b0001101001: data <= 8'h00; 
        10'b0001101010: data <= 8'h00; 
        10'b0001101011: data <= 8'h00; 
        10'b0001101100: data <= 8'h00; 
        10'b0001101101: data <= 8'h00; 
        10'b0001101110: data <= 8'h00; 
        10'b0001101111: data <= 8'h00; 
        10'b0001110000: data <= 8'h00; 
        10'b0001110001: data <= 8'h00; 
        10'b0001110010: data <= 8'h00; 
        10'b0001110011: data <= 8'h00; 
        10'b0001110100: data <= 8'h00; 
        10'b0001110101: data <= 8'h00; 
        10'b0001110110: data <= 8'h00; 
        10'b0001110111: data <= 8'h00; 
        10'b0001111000: data <= 8'h00; 
        10'b0001111001: data <= 8'h00; 
        10'b0001111010: data <= 8'h00; 
        10'b0001111011: data <= 8'h00; 
        10'b0001111100: data <= 8'h00; 
        10'b0001111101: data <= 8'h00; 
        10'b0001111110: data <= 8'h00; 
        10'b0001111111: data <= 8'h00; 
        10'b0010000000: data <= 8'h00; 
        10'b0010000001: data <= 8'h00; 
        10'b0010000010: data <= 8'h00; 
        10'b0010000011: data <= 8'h00; 
        10'b0010000100: data <= 8'h00; 
        10'b0010000101: data <= 8'h00; 
        10'b0010000110: data <= 8'h00; 
        10'b0010000111: data <= 8'h00; 
        10'b0010001000: data <= 8'h00; 
        10'b0010001001: data <= 8'h00; 
        10'b0010001010: data <= 8'h00; 
        10'b0010001011: data <= 8'h00; 
        10'b0010001100: data <= 8'h00; 
        10'b0010001101: data <= 8'h00; 
        10'b0010001110: data <= 8'h00; 
        10'b0010001111: data <= 8'h00; 
        10'b0010010000: data <= 8'h00; 
        10'b0010010001: data <= 8'h00; 
        10'b0010010010: data <= 8'h00; 
        10'b0010010011: data <= 8'h00; 
        10'b0010010100: data <= 8'h00; 
        10'b0010010101: data <= 8'h00; 
        10'b0010010110: data <= 8'h00; 
        10'b0010010111: data <= 8'h00; 
        10'b0010011000: data <= 8'h00; 
        10'b0010011001: data <= 8'h01; 
        10'b0010011010: data <= 8'h01; 
        10'b0010011011: data <= 8'h01; 
        10'b0010011100: data <= 8'h01; 
        10'b0010011101: data <= 8'h01; 
        10'b0010011110: data <= 8'h01; 
        10'b0010011111: data <= 8'h00; 
        10'b0010100000: data <= 8'h00; 
        10'b0010100001: data <= 8'h00; 
        10'b0010100010: data <= 8'h00; 
        10'b0010100011: data <= 8'h00; 
        10'b0010100100: data <= 8'h00; 
        10'b0010100101: data <= 8'h00; 
        10'b0010100110: data <= 8'h00; 
        10'b0010100111: data <= 8'h00; 
        10'b0010101000: data <= 8'h00; 
        10'b0010101001: data <= 8'h00; 
        10'b0010101010: data <= 8'h00; 
        10'b0010101011: data <= 8'h00; 
        10'b0010101100: data <= 8'h00; 
        10'b0010101101: data <= 8'h00; 
        10'b0010101110: data <= 8'h00; 
        10'b0010101111: data <= 8'h00; 
        10'b0010110000: data <= 8'h00; 
        10'b0010110001: data <= 8'h00; 
        10'b0010110010: data <= 8'h00; 
        10'b0010110011: data <= 8'h00; 
        10'b0010110100: data <= 8'h00; 
        10'b0010110101: data <= 8'h00; 
        10'b0010110110: data <= 8'h00; 
        10'b0010110111: data <= 8'h01; 
        10'b0010111000: data <= 8'h01; 
        10'b0010111001: data <= 8'h01; 
        10'b0010111010: data <= 8'h01; 
        10'b0010111011: data <= 8'h01; 
        10'b0010111100: data <= 8'h01; 
        10'b0010111101: data <= 8'h01; 
        10'b0010111110: data <= 8'h00; 
        10'b0010111111: data <= 8'h00; 
        10'b0011000000: data <= 8'h00; 
        10'b0011000001: data <= 8'h00; 
        10'b0011000010: data <= 8'h00; 
        10'b0011000011: data <= 8'h00; 
        10'b0011000100: data <= 8'h00; 
        10'b0011000101: data <= 8'h00; 
        10'b0011000110: data <= 8'h00; 
        10'b0011000111: data <= 8'h00; 
        10'b0011001000: data <= 8'h00; 
        10'b0011001001: data <= 8'h00; 
        10'b0011001010: data <= 8'h00; 
        10'b0011001011: data <= 8'h00; 
        10'b0011001100: data <= 8'h00; 
        10'b0011001101: data <= 8'h00; 
        10'b0011001110: data <= 8'h00; 
        10'b0011001111: data <= 8'h00; 
        10'b0011010000: data <= 8'h01; 
        10'b0011010001: data <= 8'h01; 
        10'b0011010010: data <= 8'h00; 
        10'b0011010011: data <= 8'h00; 
        10'b0011010100: data <= 8'h01; 
        10'b0011010101: data <= 8'h01; 
        10'b0011010110: data <= 8'h01; 
        10'b0011010111: data <= 8'h01; 
        10'b0011011000: data <= 8'h00; 
        10'b0011011001: data <= 8'h00; 
        10'b0011011010: data <= 8'h01; 
        10'b0011011011: data <= 8'h00; 
        10'b0011011100: data <= 8'h00; 
        10'b0011011101: data <= 8'h00; 
        10'b0011011110: data <= 8'h00; 
        10'b0011011111: data <= 8'h00; 
        10'b0011100000: data <= 8'h00; 
        10'b0011100001: data <= 8'h00; 
        10'b0011100010: data <= 8'h00; 
        10'b0011100011: data <= 8'h00; 
        10'b0011100100: data <= 8'h00; 
        10'b0011100101: data <= 8'h00; 
        10'b0011100110: data <= 8'h00; 
        10'b0011100111: data <= 8'h00; 
        10'b0011101000: data <= 8'h00; 
        10'b0011101001: data <= 8'h00; 
        10'b0011101010: data <= 8'h00; 
        10'b0011101011: data <= 8'h00; 
        10'b0011101100: data <= 8'h00; 
        10'b0011101101: data <= 8'h00; 
        10'b0011101110: data <= 8'h00; 
        10'b0011101111: data <= 8'h00; 
        10'b0011110000: data <= 8'h01; 
        10'b0011110001: data <= 8'h01; 
        10'b0011110010: data <= 8'h01; 
        10'b0011110011: data <= 8'h00; 
        10'b0011110100: data <= 8'h00; 
        10'b0011110101: data <= 8'h00; 
        10'b0011110110: data <= 8'h01; 
        10'b0011110111: data <= 8'h01; 
        10'b0011111000: data <= 8'h00; 
        10'b0011111001: data <= 8'h00; 
        10'b0011111010: data <= 8'h00; 
        10'b0011111011: data <= 8'h00; 
        10'b0011111100: data <= 8'h00; 
        10'b0011111101: data <= 8'h00; 
        10'b0011111110: data <= 8'h00; 
        10'b0011111111: data <= 8'h00; 
        10'b0100000000: data <= 8'h00; 
        10'b0100000001: data <= 8'h00; 
        10'b0100000010: data <= 8'h00; 
        10'b0100000011: data <= 8'h00; 
        10'b0100000100: data <= 8'h00; 
        10'b0100000101: data <= 8'h00; 
        10'b0100000110: data <= 8'h00; 
        10'b0100000111: data <= 8'h00; 
        10'b0100001000: data <= 8'h00; 
        10'b0100001001: data <= 8'h00; 
        10'b0100001010: data <= 8'h00; 
        10'b0100001011: data <= 8'h00; 
        10'b0100001100: data <= 8'h01; 
        10'b0100001101: data <= 8'h01; 
        10'b0100001110: data <= 8'h01; 
        10'b0100001111: data <= 8'h01; 
        10'b0100010000: data <= 8'h00; 
        10'b0100010001: data <= 8'h00; 
        10'b0100010010: data <= 8'h00; 
        10'b0100010011: data <= 8'h01; 
        10'b0100010100: data <= 8'h00; 
        10'b0100010101: data <= 8'h00; 
        10'b0100010110: data <= 8'h00; 
        10'b0100010111: data <= 8'h00; 
        10'b0100011000: data <= 8'h00; 
        10'b0100011001: data <= 8'h00; 
        10'b0100011010: data <= 8'h00; 
        10'b0100011011: data <= 8'h00; 
        10'b0100011100: data <= 8'h00; 
        10'b0100011101: data <= 8'h00; 
        10'b0100011110: data <= 8'h00; 
        10'b0100011111: data <= 8'h00; 
        10'b0100100000: data <= 8'h00; 
        10'b0100100001: data <= 8'h00; 
        10'b0100100010: data <= 8'h00; 
        10'b0100100011: data <= 8'h00; 
        10'b0100100100: data <= 8'h00; 
        10'b0100100101: data <= 8'h00; 
        10'b0100100110: data <= 8'h00; 
        10'b0100100111: data <= 8'hff; 
        10'b0100101000: data <= 8'h00; 
        10'b0100101001: data <= 8'h00; 
        10'b0100101010: data <= 8'h01; 
        10'b0100101011: data <= 8'h01; 
        10'b0100101100: data <= 8'h01; 
        10'b0100101101: data <= 8'h01; 
        10'b0100101110: data <= 8'h01; 
        10'b0100101111: data <= 8'h01; 
        10'b0100110000: data <= 8'h01; 
        10'b0100110001: data <= 8'h00; 
        10'b0100110010: data <= 8'h00; 
        10'b0100110011: data <= 8'h00; 
        10'b0100110100: data <= 8'h00; 
        10'b0100110101: data <= 8'h00; 
        10'b0100110110: data <= 8'h00; 
        10'b0100110111: data <= 8'h00; 
        10'b0100111000: data <= 8'h00; 
        10'b0100111001: data <= 8'h00; 
        10'b0100111010: data <= 8'h00; 
        10'b0100111011: data <= 8'h00; 
        10'b0100111100: data <= 8'h00; 
        10'b0100111101: data <= 8'h00; 
        10'b0100111110: data <= 8'h00; 
        10'b0100111111: data <= 8'h00; 
        10'b0101000000: data <= 8'h00; 
        10'b0101000001: data <= 8'h00; 
        10'b0101000010: data <= 8'hff; 
        10'b0101000011: data <= 8'hfe; 
        10'b0101000100: data <= 8'hfe; 
        10'b0101000101: data <= 8'hff; 
        10'b0101000110: data <= 8'h00; 
        10'b0101000111: data <= 8'h00; 
        10'b0101001000: data <= 8'h01; 
        10'b0101001001: data <= 8'h01; 
        10'b0101001010: data <= 8'h01; 
        10'b0101001011: data <= 8'h01; 
        10'b0101001100: data <= 8'h01; 
        10'b0101001101: data <= 8'h00; 
        10'b0101001110: data <= 8'h00; 
        10'b0101001111: data <= 8'h00; 
        10'b0101010000: data <= 8'h00; 
        10'b0101010001: data <= 8'h00; 
        10'b0101010010: data <= 8'h00; 
        10'b0101010011: data <= 8'h00; 
        10'b0101010100: data <= 8'h00; 
        10'b0101010101: data <= 8'h00; 
        10'b0101010110: data <= 8'h00; 
        10'b0101010111: data <= 8'h00; 
        10'b0101011000: data <= 8'h00; 
        10'b0101011001: data <= 8'h00; 
        10'b0101011010: data <= 8'h00; 
        10'b0101011011: data <= 8'h00; 
        10'b0101011100: data <= 8'h00; 
        10'b0101011101: data <= 8'h00; 
        10'b0101011110: data <= 8'hfe; 
        10'b0101011111: data <= 8'hfe; 
        10'b0101100000: data <= 8'hfe; 
        10'b0101100001: data <= 8'hff; 
        10'b0101100010: data <= 8'h00; 
        10'b0101100011: data <= 8'h00; 
        10'b0101100100: data <= 8'h00; 
        10'b0101100101: data <= 8'h00; 
        10'b0101100110: data <= 8'h01; 
        10'b0101100111: data <= 8'h01; 
        10'b0101101000: data <= 8'h01; 
        10'b0101101001: data <= 8'h00; 
        10'b0101101010: data <= 8'h00; 
        10'b0101101011: data <= 8'h00; 
        10'b0101101100: data <= 8'h00; 
        10'b0101101101: data <= 8'h00; 
        10'b0101101110: data <= 8'h00; 
        10'b0101101111: data <= 8'h00; 
        10'b0101110000: data <= 8'h00; 
        10'b0101110001: data <= 8'h00; 
        10'b0101110010: data <= 8'h00; 
        10'b0101110011: data <= 8'h01; 
        10'b0101110100: data <= 8'h00; 
        10'b0101110101: data <= 8'h00; 
        10'b0101110110: data <= 8'h00; 
        10'b0101110111: data <= 8'h00; 
        10'b0101111000: data <= 8'h00; 
        10'b0101111001: data <= 8'hff; 
        10'b0101111010: data <= 8'hfe; 
        10'b0101111011: data <= 8'hfe; 
        10'b0101111100: data <= 8'hfe; 
        10'b0101111101: data <= 8'hff; 
        10'b0101111110: data <= 8'h00; 
        10'b0101111111: data <= 8'hff; 
        10'b0110000000: data <= 8'h00; 
        10'b0110000001: data <= 8'h00; 
        10'b0110000010: data <= 8'h01; 
        10'b0110000011: data <= 8'h01; 
        10'b0110000100: data <= 8'h01; 
        10'b0110000101: data <= 8'h00; 
        10'b0110000110: data <= 8'h00; 
        10'b0110000111: data <= 8'h00; 
        10'b0110001000: data <= 8'h00; 
        10'b0110001001: data <= 8'h00; 
        10'b0110001010: data <= 8'h00; 
        10'b0110001011: data <= 8'h00; 
        10'b0110001100: data <= 8'h00; 
        10'b0110001101: data <= 8'h01; 
        10'b0110001110: data <= 8'h01; 
        10'b0110001111: data <= 8'h01; 
        10'b0110010000: data <= 8'h00; 
        10'b0110010001: data <= 8'h01; 
        10'b0110010010: data <= 8'h01; 
        10'b0110010011: data <= 8'h00; 
        10'b0110010100: data <= 8'h00; 
        10'b0110010101: data <= 8'hff; 
        10'b0110010110: data <= 8'hfe; 
        10'b0110010111: data <= 8'hfe; 
        10'b0110011000: data <= 8'hfe; 
        10'b0110011001: data <= 8'hff; 
        10'b0110011010: data <= 8'h00; 
        10'b0110011011: data <= 8'hff; 
        10'b0110011100: data <= 8'h00; 
        10'b0110011101: data <= 8'h00; 
        10'b0110011110: data <= 8'h01; 
        10'b0110011111: data <= 8'h01; 
        10'b0110100000: data <= 8'h01; 
        10'b0110100001: data <= 8'h00; 
        10'b0110100010: data <= 8'h00; 
        10'b0110100011: data <= 8'h00; 
        10'b0110100100: data <= 8'h00; 
        10'b0110100101: data <= 8'h00; 
        10'b0110100110: data <= 8'h00; 
        10'b0110100111: data <= 8'h00; 
        10'b0110101000: data <= 8'h00; 
        10'b0110101001: data <= 8'h01; 
        10'b0110101010: data <= 8'h01; 
        10'b0110101011: data <= 8'h01; 
        10'b0110101100: data <= 8'h01; 
        10'b0110101101: data <= 8'h01; 
        10'b0110101110: data <= 8'h01; 
        10'b0110101111: data <= 8'h00; 
        10'b0110110000: data <= 8'hff; 
        10'b0110110001: data <= 8'hfe; 
        10'b0110110010: data <= 8'hfe; 
        10'b0110110011: data <= 8'hfe; 
        10'b0110110100: data <= 8'hfe; 
        10'b0110110101: data <= 8'hff; 
        10'b0110110110: data <= 8'h00; 
        10'b0110110111: data <= 8'h00; 
        10'b0110111000: data <= 8'h00; 
        10'b0110111001: data <= 8'h00; 
        10'b0110111010: data <= 8'h01; 
        10'b0110111011: data <= 8'h01; 
        10'b0110111100: data <= 8'h00; 
        10'b0110111101: data <= 8'h00; 
        10'b0110111110: data <= 8'h00; 
        10'b0110111111: data <= 8'h00; 
        10'b0111000000: data <= 8'h00; 
        10'b0111000001: data <= 8'h00; 
        10'b0111000010: data <= 8'h00; 
        10'b0111000011: data <= 8'h00; 
        10'b0111000100: data <= 8'h00; 
        10'b0111000101: data <= 8'h01; 
        10'b0111000110: data <= 8'h01; 
        10'b0111000111: data <= 8'h01; 
        10'b0111001000: data <= 8'h00; 
        10'b0111001001: data <= 8'h00; 
        10'b0111001010: data <= 8'h01; 
        10'b0111001011: data <= 8'h00; 
        10'b0111001100: data <= 8'hff; 
        10'b0111001101: data <= 8'hfe; 
        10'b0111001110: data <= 8'hfe; 
        10'b0111001111: data <= 8'hfe; 
        10'b0111010000: data <= 8'hff; 
        10'b0111010001: data <= 8'h00; 
        10'b0111010010: data <= 8'h00; 
        10'b0111010011: data <= 8'h00; 
        10'b0111010100: data <= 8'h00; 
        10'b0111010101: data <= 8'h01; 
        10'b0111010110: data <= 8'h01; 
        10'b0111010111: data <= 8'h01; 
        10'b0111011000: data <= 8'h00; 
        10'b0111011001: data <= 8'h00; 
        10'b0111011010: data <= 8'h00; 
        10'b0111011011: data <= 8'h00; 
        10'b0111011100: data <= 8'h00; 
        10'b0111011101: data <= 8'h00; 
        10'b0111011110: data <= 8'h00; 
        10'b0111011111: data <= 8'h00; 
        10'b0111100000: data <= 8'h00; 
        10'b0111100001: data <= 8'h01; 
        10'b0111100010: data <= 8'h01; 
        10'b0111100011: data <= 8'h01; 
        10'b0111100100: data <= 8'h00; 
        10'b0111100101: data <= 8'h01; 
        10'b0111100110: data <= 8'h01; 
        10'b0111100111: data <= 8'h00; 
        10'b0111101000: data <= 8'hfe; 
        10'b0111101001: data <= 8'hfe; 
        10'b0111101010: data <= 8'hfe; 
        10'b0111101011: data <= 8'hff; 
        10'b0111101100: data <= 8'h00; 
        10'b0111101101: data <= 8'h00; 
        10'b0111101110: data <= 8'h00; 
        10'b0111101111: data <= 8'h00; 
        10'b0111110000: data <= 8'h01; 
        10'b0111110001: data <= 8'h00; 
        10'b0111110010: data <= 8'h00; 
        10'b0111110011: data <= 8'h00; 
        10'b0111110100: data <= 8'h00; 
        10'b0111110101: data <= 8'h00; 
        10'b0111110110: data <= 8'h00; 
        10'b0111110111: data <= 8'h00; 
        10'b0111111000: data <= 8'h00; 
        10'b0111111001: data <= 8'h00; 
        10'b0111111010: data <= 8'h00; 
        10'b0111111011: data <= 8'h00; 
        10'b0111111100: data <= 8'h00; 
        10'b0111111101: data <= 8'h00; 
        10'b0111111110: data <= 8'h01; 
        10'b0111111111: data <= 8'h00; 
        10'b1000000000: data <= 8'h00; 
        10'b1000000001: data <= 8'h01; 
        10'b1000000010: data <= 8'h01; 
        10'b1000000011: data <= 8'h00; 
        10'b1000000100: data <= 8'hff; 
        10'b1000000101: data <= 8'hfe; 
        10'b1000000110: data <= 8'hff; 
        10'b1000000111: data <= 8'h00; 
        10'b1000001000: data <= 8'h00; 
        10'b1000001001: data <= 8'h00; 
        10'b1000001010: data <= 8'h00; 
        10'b1000001011: data <= 8'h00; 
        10'b1000001100: data <= 8'h00; 
        10'b1000001101: data <= 8'h00; 
        10'b1000001110: data <= 8'h00; 
        10'b1000001111: data <= 8'h00; 
        10'b1000010000: data <= 8'h00; 
        10'b1000010001: data <= 8'h00; 
        10'b1000010010: data <= 8'h00; 
        10'b1000010011: data <= 8'h00; 
        10'b1000010100: data <= 8'h00; 
        10'b1000010101: data <= 8'h00; 
        10'b1000010110: data <= 8'h00; 
        10'b1000010111: data <= 8'h00; 
        10'b1000011000: data <= 8'h00; 
        10'b1000011001: data <= 8'h00; 
        10'b1000011010: data <= 8'h01; 
        10'b1000011011: data <= 8'h01; 
        10'b1000011100: data <= 8'h01; 
        10'b1000011101: data <= 8'h01; 
        10'b1000011110: data <= 8'h01; 
        10'b1000011111: data <= 8'h01; 
        10'b1000100000: data <= 8'h00; 
        10'b1000100001: data <= 8'h00; 
        10'b1000100010: data <= 8'h00; 
        10'b1000100011: data <= 8'h00; 
        10'b1000100100: data <= 8'h00; 
        10'b1000100101: data <= 8'h00; 
        10'b1000100110: data <= 8'h00; 
        10'b1000100111: data <= 8'h00; 
        10'b1000101000: data <= 8'h00; 
        10'b1000101001: data <= 8'h00; 
        10'b1000101010: data <= 8'h00; 
        10'b1000101011: data <= 8'h00; 
        10'b1000101100: data <= 8'h00; 
        10'b1000101101: data <= 8'h00; 
        10'b1000101110: data <= 8'h00; 
        10'b1000101111: data <= 8'h00; 
        10'b1000110000: data <= 8'h00; 
        10'b1000110001: data <= 8'h00; 
        10'b1000110010: data <= 8'h00; 
        10'b1000110011: data <= 8'h00; 
        10'b1000110100: data <= 8'h00; 
        10'b1000110101: data <= 8'h00; 
        10'b1000110110: data <= 8'h01; 
        10'b1000110111: data <= 8'h01; 
        10'b1000111000: data <= 8'h01; 
        10'b1000111001: data <= 8'h01; 
        10'b1000111010: data <= 8'h01; 
        10'b1000111011: data <= 8'h01; 
        10'b1000111100: data <= 8'h01; 
        10'b1000111101: data <= 8'h00; 
        10'b1000111110: data <= 8'h00; 
        10'b1000111111: data <= 8'h00; 
        10'b1001000000: data <= 8'h00; 
        10'b1001000001: data <= 8'h00; 
        10'b1001000010: data <= 8'h00; 
        10'b1001000011: data <= 8'h00; 
        10'b1001000100: data <= 8'h00; 
        10'b1001000101: data <= 8'h00; 
        10'b1001000110: data <= 8'h00; 
        10'b1001000111: data <= 8'h00; 
        10'b1001001000: data <= 8'h00; 
        10'b1001001001: data <= 8'h00; 
        10'b1001001010: data <= 8'h00; 
        10'b1001001011: data <= 8'h00; 
        10'b1001001100: data <= 8'h00; 
        10'b1001001101: data <= 8'h00; 
        10'b1001001110: data <= 8'h00; 
        10'b1001001111: data <= 8'h00; 
        10'b1001010000: data <= 8'h00; 
        10'b1001010001: data <= 8'h00; 
        10'b1001010010: data <= 8'h00; 
        10'b1001010011: data <= 8'h01; 
        10'b1001010100: data <= 8'h00; 
        10'b1001010101: data <= 8'h01; 
        10'b1001010110: data <= 8'h01; 
        10'b1001010111: data <= 8'h01; 
        10'b1001011000: data <= 8'h01; 
        10'b1001011001: data <= 8'h00; 
        10'b1001011010: data <= 8'h00; 
        10'b1001011011: data <= 8'h00; 
        10'b1001011100: data <= 8'h00; 
        10'b1001011101: data <= 8'h00; 
        10'b1001011110: data <= 8'h00; 
        10'b1001011111: data <= 8'h00; 
        10'b1001100000: data <= 8'h00; 
        10'b1001100001: data <= 8'h00; 
        10'b1001100010: data <= 8'h00; 
        10'b1001100011: data <= 8'h00; 
        10'b1001100100: data <= 8'h00; 
        10'b1001100101: data <= 8'h00; 
        10'b1001100110: data <= 8'h00; 
        10'b1001100111: data <= 8'h00; 
        10'b1001101000: data <= 8'h00; 
        10'b1001101001: data <= 8'h00; 
        10'b1001101010: data <= 8'h00; 
        10'b1001101011: data <= 8'h00; 
        10'b1001101100: data <= 8'h00; 
        10'b1001101101: data <= 8'h00; 
        10'b1001101110: data <= 8'h00; 
        10'b1001101111: data <= 8'h00; 
        10'b1001110000: data <= 8'h01; 
        10'b1001110001: data <= 8'h01; 
        10'b1001110010: data <= 8'h01; 
        10'b1001110011: data <= 8'h01; 
        10'b1001110100: data <= 8'h01; 
        10'b1001110101: data <= 8'h01; 
        10'b1001110110: data <= 8'h00; 
        10'b1001110111: data <= 8'h00; 
        10'b1001111000: data <= 8'h00; 
        10'b1001111001: data <= 8'h00; 
        10'b1001111010: data <= 8'h00; 
        10'b1001111011: data <= 8'h00; 
        10'b1001111100: data <= 8'h00; 
        10'b1001111101: data <= 8'h00; 
        10'b1001111110: data <= 8'h00; 
        10'b1001111111: data <= 8'h00; 
        10'b1010000000: data <= 8'h00; 
        10'b1010000001: data <= 8'h00; 
        10'b1010000010: data <= 8'h00; 
        10'b1010000011: data <= 8'h00; 
        10'b1010000100: data <= 8'h00; 
        10'b1010000101: data <= 8'h00; 
        10'b1010000110: data <= 8'h00; 
        10'b1010000111: data <= 8'h00; 
        10'b1010001000: data <= 8'h00; 
        10'b1010001001: data <= 8'h00; 
        10'b1010001010: data <= 8'h00; 
        10'b1010001011: data <= 8'h00; 
        10'b1010001100: data <= 8'h00; 
        10'b1010001101: data <= 8'h01; 
        10'b1010001110: data <= 8'h01; 
        10'b1010001111: data <= 8'h01; 
        10'b1010010000: data <= 8'h01; 
        10'b1010010001: data <= 8'h01; 
        10'b1010010010: data <= 8'h01; 
        10'b1010010011: data <= 8'h00; 
        10'b1010010100: data <= 8'h00; 
        10'b1010010101: data <= 8'h00; 
        10'b1010010110: data <= 8'h00; 
        10'b1010010111: data <= 8'hff; 
        10'b1010011000: data <= 8'h00; 
        10'b1010011001: data <= 8'h00; 
        10'b1010011010: data <= 8'h00; 
        10'b1010011011: data <= 8'h00; 
        10'b1010011100: data <= 8'h00; 
        10'b1010011101: data <= 8'h00; 
        10'b1010011110: data <= 8'h00; 
        10'b1010011111: data <= 8'h00; 
        10'b1010100000: data <= 8'h00; 
        10'b1010100001: data <= 8'h00; 
        10'b1010100010: data <= 8'h00; 
        10'b1010100011: data <= 8'h00; 
        10'b1010100100: data <= 8'h00; 
        10'b1010100101: data <= 8'h00; 
        10'b1010100110: data <= 8'h00; 
        10'b1010100111: data <= 8'h00; 
        10'b1010101000: data <= 8'h00; 
        10'b1010101001: data <= 8'h00; 
        10'b1010101010: data <= 8'h00; 
        10'b1010101011: data <= 8'h00; 
        10'b1010101100: data <= 8'h00; 
        10'b1010101101: data <= 8'h00; 
        10'b1010101110: data <= 8'h00; 
        10'b1010101111: data <= 8'h00; 
        10'b1010110000: data <= 8'h00; 
        10'b1010110001: data <= 8'h00; 
        10'b1010110010: data <= 8'h00; 
        10'b1010110011: data <= 8'h00; 
        10'b1010110100: data <= 8'h00; 
        10'b1010110101: data <= 8'h00; 
        10'b1010110110: data <= 8'h00; 
        10'b1010110111: data <= 8'h00; 
        10'b1010111000: data <= 8'h00; 
        10'b1010111001: data <= 8'h00; 
        10'b1010111010: data <= 8'h00; 
        10'b1010111011: data <= 8'h00; 
        10'b1010111100: data <= 8'h00; 
        10'b1010111101: data <= 8'h00; 
        10'b1010111110: data <= 8'h00; 
        10'b1010111111: data <= 8'h00; 
        10'b1011000000: data <= 8'h00; 
        10'b1011000001: data <= 8'h00; 
        10'b1011000010: data <= 8'h00; 
        10'b1011000011: data <= 8'h00; 
        10'b1011000100: data <= 8'h00; 
        10'b1011000101: data <= 8'h00; 
        10'b1011000110: data <= 8'h00; 
        10'b1011000111: data <= 8'hff; 
        10'b1011001000: data <= 8'hff; 
        10'b1011001001: data <= 8'hff; 
        10'b1011001010: data <= 8'hff; 
        10'b1011001011: data <= 8'hff; 
        10'b1011001100: data <= 8'hff; 
        10'b1011001101: data <= 8'h00; 
        10'b1011001110: data <= 8'h00; 
        10'b1011001111: data <= 8'h00; 
        10'b1011010000: data <= 8'h00; 
        10'b1011010001: data <= 8'h00; 
        10'b1011010010: data <= 8'h00; 
        10'b1011010011: data <= 8'h00; 
        10'b1011010100: data <= 8'h00; 
        10'b1011010101: data <= 8'h00; 
        10'b1011010110: data <= 8'h00; 
        10'b1011010111: data <= 8'h00; 
        10'b1011011000: data <= 8'h00; 
        10'b1011011001: data <= 8'h00; 
        10'b1011011010: data <= 8'h00; 
        10'b1011011011: data <= 8'h00; 
        10'b1011011100: data <= 8'h00; 
        10'b1011011101: data <= 8'h00; 
        10'b1011011110: data <= 8'h00; 
        10'b1011011111: data <= 8'h00; 
        10'b1011100000: data <= 8'h00; 
        10'b1011100001: data <= 8'h00; 
        10'b1011100010: data <= 8'h00; 
        10'b1011100011: data <= 8'h00; 
        10'b1011100100: data <= 8'h00; 
        10'b1011100101: data <= 8'h00; 
        10'b1011100110: data <= 8'h00; 
        10'b1011100111: data <= 8'h00; 
        10'b1011101000: data <= 8'h00; 
        10'b1011101001: data <= 8'h00; 
        10'b1011101010: data <= 8'h00; 
        10'b1011101011: data <= 8'h00; 
        10'b1011101100: data <= 8'h00; 
        10'b1011101101: data <= 8'h00; 
        10'b1011101110: data <= 8'h00; 
        10'b1011101111: data <= 8'h00; 
        10'b1011110000: data <= 8'h00; 
        10'b1011110001: data <= 8'h00; 
        10'b1011110010: data <= 8'h00; 
        10'b1011110011: data <= 8'h00; 
        10'b1011110100: data <= 8'h00; 
        10'b1011110101: data <= 8'h00; 
        10'b1011110110: data <= 8'h00; 
        10'b1011110111: data <= 8'h00; 
        10'b1011111000: data <= 8'h00; 
        10'b1011111001: data <= 8'h00; 
        10'b1011111010: data <= 8'h00; 
        10'b1011111011: data <= 8'h00; 
        10'b1011111100: data <= 8'h00; 
        10'b1011111101: data <= 8'h00; 
        10'b1011111110: data <= 8'h00; 
        10'b1011111111: data <= 8'h00; 
        10'b1100000000: data <= 8'h00; 
        10'b1100000001: data <= 8'h00; 
        10'b1100000010: data <= 8'h00; 
        10'b1100000011: data <= 8'h00; 
        10'b1100000100: data <= 8'h00; 
        10'b1100000101: data <= 8'h00; 
        10'b1100000110: data <= 8'h00; 
        10'b1100000111: data <= 8'h00; 
        10'b1100001000: data <= 8'h00; 
        10'b1100001001: data <= 8'h00; 
        10'b1100001010: data <= 8'h00; 
        10'b1100001011: data <= 8'h00; 
        10'b1100001100: data <= 8'h00; 
        10'b1100001101: data <= 8'h00; 
        10'b1100001110: data <= 8'h00; 
        10'b1100001111: data <= 8'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 3) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 9'h000; 
        10'b0000000001: data <= 9'h000; 
        10'b0000000010: data <= 9'h000; 
        10'b0000000011: data <= 9'h000; 
        10'b0000000100: data <= 9'h000; 
        10'b0000000101: data <= 9'h000; 
        10'b0000000110: data <= 9'h000; 
        10'b0000000111: data <= 9'h000; 
        10'b0000001000: data <= 9'h000; 
        10'b0000001001: data <= 9'h000; 
        10'b0000001010: data <= 9'h000; 
        10'b0000001011: data <= 9'h000; 
        10'b0000001100: data <= 9'h000; 
        10'b0000001101: data <= 9'h000; 
        10'b0000001110: data <= 9'h000; 
        10'b0000001111: data <= 9'h000; 
        10'b0000010000: data <= 9'h000; 
        10'b0000010001: data <= 9'h000; 
        10'b0000010010: data <= 9'h000; 
        10'b0000010011: data <= 9'h000; 
        10'b0000010100: data <= 9'h000; 
        10'b0000010101: data <= 9'h000; 
        10'b0000010110: data <= 9'h000; 
        10'b0000010111: data <= 9'h000; 
        10'b0000011000: data <= 9'h000; 
        10'b0000011001: data <= 9'h000; 
        10'b0000011010: data <= 9'h000; 
        10'b0000011011: data <= 9'h000; 
        10'b0000011100: data <= 9'h000; 
        10'b0000011101: data <= 9'h000; 
        10'b0000011110: data <= 9'h000; 
        10'b0000011111: data <= 9'h000; 
        10'b0000100000: data <= 9'h000; 
        10'b0000100001: data <= 9'h000; 
        10'b0000100010: data <= 9'h000; 
        10'b0000100011: data <= 9'h000; 
        10'b0000100100: data <= 9'h000; 
        10'b0000100101: data <= 9'h000; 
        10'b0000100110: data <= 9'h000; 
        10'b0000100111: data <= 9'h000; 
        10'b0000101000: data <= 9'h000; 
        10'b0000101001: data <= 9'h000; 
        10'b0000101010: data <= 9'h000; 
        10'b0000101011: data <= 9'h000; 
        10'b0000101100: data <= 9'h000; 
        10'b0000101101: data <= 9'h000; 
        10'b0000101110: data <= 9'h000; 
        10'b0000101111: data <= 9'h000; 
        10'b0000110000: data <= 9'h000; 
        10'b0000110001: data <= 9'h000; 
        10'b0000110010: data <= 9'h000; 
        10'b0000110011: data <= 9'h000; 
        10'b0000110100: data <= 9'h000; 
        10'b0000110101: data <= 9'h000; 
        10'b0000110110: data <= 9'h000; 
        10'b0000110111: data <= 9'h000; 
        10'b0000111000: data <= 9'h000; 
        10'b0000111001: data <= 9'h000; 
        10'b0000111010: data <= 9'h000; 
        10'b0000111011: data <= 9'h000; 
        10'b0000111100: data <= 9'h000; 
        10'b0000111101: data <= 9'h000; 
        10'b0000111110: data <= 9'h000; 
        10'b0000111111: data <= 9'h000; 
        10'b0001000000: data <= 9'h000; 
        10'b0001000001: data <= 9'h000; 
        10'b0001000010: data <= 9'h000; 
        10'b0001000011: data <= 9'h000; 
        10'b0001000100: data <= 9'h000; 
        10'b0001000101: data <= 9'h000; 
        10'b0001000110: data <= 9'h000; 
        10'b0001000111: data <= 9'h1ff; 
        10'b0001001000: data <= 9'h000; 
        10'b0001001001: data <= 9'h000; 
        10'b0001001010: data <= 9'h000; 
        10'b0001001011: data <= 9'h000; 
        10'b0001001100: data <= 9'h000; 
        10'b0001001101: data <= 9'h000; 
        10'b0001001110: data <= 9'h000; 
        10'b0001001111: data <= 9'h000; 
        10'b0001010000: data <= 9'h000; 
        10'b0001010001: data <= 9'h000; 
        10'b0001010010: data <= 9'h000; 
        10'b0001010011: data <= 9'h000; 
        10'b0001010100: data <= 9'h000; 
        10'b0001010101: data <= 9'h000; 
        10'b0001010110: data <= 9'h000; 
        10'b0001010111: data <= 9'h000; 
        10'b0001011000: data <= 9'h000; 
        10'b0001011001: data <= 9'h000; 
        10'b0001011010: data <= 9'h000; 
        10'b0001011011: data <= 9'h000; 
        10'b0001011100: data <= 9'h000; 
        10'b0001011101: data <= 9'h000; 
        10'b0001011110: data <= 9'h000; 
        10'b0001011111: data <= 9'h000; 
        10'b0001100000: data <= 9'h1ff; 
        10'b0001100001: data <= 9'h000; 
        10'b0001100010: data <= 9'h000; 
        10'b0001100011: data <= 9'h1ff; 
        10'b0001100100: data <= 9'h000; 
        10'b0001100101: data <= 9'h000; 
        10'b0001100110: data <= 9'h1ff; 
        10'b0001100111: data <= 9'h1ff; 
        10'b0001101000: data <= 9'h1ff; 
        10'b0001101001: data <= 9'h1ff; 
        10'b0001101010: data <= 9'h1ff; 
        10'b0001101011: data <= 9'h000; 
        10'b0001101100: data <= 9'h000; 
        10'b0001101101: data <= 9'h000; 
        10'b0001101110: data <= 9'h000; 
        10'b0001101111: data <= 9'h000; 
        10'b0001110000: data <= 9'h000; 
        10'b0001110001: data <= 9'h000; 
        10'b0001110010: data <= 9'h000; 
        10'b0001110011: data <= 9'h000; 
        10'b0001110100: data <= 9'h000; 
        10'b0001110101: data <= 9'h000; 
        10'b0001110110: data <= 9'h000; 
        10'b0001110111: data <= 9'h000; 
        10'b0001111000: data <= 9'h000; 
        10'b0001111001: data <= 9'h000; 
        10'b0001111010: data <= 9'h1ff; 
        10'b0001111011: data <= 9'h1ff; 
        10'b0001111100: data <= 9'h1ff; 
        10'b0001111101: data <= 9'h1ff; 
        10'b0001111110: data <= 9'h000; 
        10'b0001111111: data <= 9'h000; 
        10'b0010000000: data <= 9'h000; 
        10'b0010000001: data <= 9'h000; 
        10'b0010000010: data <= 9'h000; 
        10'b0010000011: data <= 9'h1ff; 
        10'b0010000100: data <= 9'h000; 
        10'b0010000101: data <= 9'h1ff; 
        10'b0010000110: data <= 9'h000; 
        10'b0010000111: data <= 9'h000; 
        10'b0010001000: data <= 9'h000; 
        10'b0010001001: data <= 9'h000; 
        10'b0010001010: data <= 9'h000; 
        10'b0010001011: data <= 9'h000; 
        10'b0010001100: data <= 9'h000; 
        10'b0010001101: data <= 9'h000; 
        10'b0010001110: data <= 9'h000; 
        10'b0010001111: data <= 9'h000; 
        10'b0010010000: data <= 9'h000; 
        10'b0010010001: data <= 9'h000; 
        10'b0010010010: data <= 9'h000; 
        10'b0010010011: data <= 9'h000; 
        10'b0010010100: data <= 9'h000; 
        10'b0010010101: data <= 9'h000; 
        10'b0010010110: data <= 9'h000; 
        10'b0010010111: data <= 9'h000; 
        10'b0010011000: data <= 9'h000; 
        10'b0010011001: data <= 9'h001; 
        10'b0010011010: data <= 9'h001; 
        10'b0010011011: data <= 9'h001; 
        10'b0010011100: data <= 9'h001; 
        10'b0010011101: data <= 9'h001; 
        10'b0010011110: data <= 9'h002; 
        10'b0010011111: data <= 9'h001; 
        10'b0010100000: data <= 9'h000; 
        10'b0010100001: data <= 9'h000; 
        10'b0010100010: data <= 9'h000; 
        10'b0010100011: data <= 9'h000; 
        10'b0010100100: data <= 9'h1ff; 
        10'b0010100101: data <= 9'h000; 
        10'b0010100110: data <= 9'h000; 
        10'b0010100111: data <= 9'h000; 
        10'b0010101000: data <= 9'h000; 
        10'b0010101001: data <= 9'h000; 
        10'b0010101010: data <= 9'h000; 
        10'b0010101011: data <= 9'h000; 
        10'b0010101100: data <= 9'h000; 
        10'b0010101101: data <= 9'h000; 
        10'b0010101110: data <= 9'h000; 
        10'b0010101111: data <= 9'h000; 
        10'b0010110000: data <= 9'h000; 
        10'b0010110001: data <= 9'h1ff; 
        10'b0010110010: data <= 9'h000; 
        10'b0010110011: data <= 9'h000; 
        10'b0010110100: data <= 9'h001; 
        10'b0010110101: data <= 9'h001; 
        10'b0010110110: data <= 9'h001; 
        10'b0010110111: data <= 9'h001; 
        10'b0010111000: data <= 9'h001; 
        10'b0010111001: data <= 9'h002; 
        10'b0010111010: data <= 9'h002; 
        10'b0010111011: data <= 9'h001; 
        10'b0010111100: data <= 9'h001; 
        10'b0010111101: data <= 9'h002; 
        10'b0010111110: data <= 9'h001; 
        10'b0010111111: data <= 9'h000; 
        10'b0011000000: data <= 9'h1ff; 
        10'b0011000001: data <= 9'h1ff; 
        10'b0011000010: data <= 9'h000; 
        10'b0011000011: data <= 9'h000; 
        10'b0011000100: data <= 9'h000; 
        10'b0011000101: data <= 9'h000; 
        10'b0011000110: data <= 9'h000; 
        10'b0011000111: data <= 9'h000; 
        10'b0011001000: data <= 9'h1ff; 
        10'b0011001001: data <= 9'h000; 
        10'b0011001010: data <= 9'h000; 
        10'b0011001011: data <= 9'h000; 
        10'b0011001100: data <= 9'h000; 
        10'b0011001101: data <= 9'h000; 
        10'b0011001110: data <= 9'h000; 
        10'b0011001111: data <= 9'h001; 
        10'b0011010000: data <= 9'h001; 
        10'b0011010001: data <= 9'h001; 
        10'b0011010010: data <= 9'h000; 
        10'b0011010011: data <= 9'h001; 
        10'b0011010100: data <= 9'h001; 
        10'b0011010101: data <= 9'h002; 
        10'b0011010110: data <= 9'h001; 
        10'b0011010111: data <= 9'h001; 
        10'b0011011000: data <= 9'h001; 
        10'b0011011001: data <= 9'h001; 
        10'b0011011010: data <= 9'h001; 
        10'b0011011011: data <= 9'h001; 
        10'b0011011100: data <= 9'h000; 
        10'b0011011101: data <= 9'h1ff; 
        10'b0011011110: data <= 9'h1ff; 
        10'b0011011111: data <= 9'h000; 
        10'b0011100000: data <= 9'h000; 
        10'b0011100001: data <= 9'h000; 
        10'b0011100010: data <= 9'h000; 
        10'b0011100011: data <= 9'h000; 
        10'b0011100100: data <= 9'h000; 
        10'b0011100101: data <= 9'h000; 
        10'b0011100110: data <= 9'h000; 
        10'b0011100111: data <= 9'h000; 
        10'b0011101000: data <= 9'h000; 
        10'b0011101001: data <= 9'h000; 
        10'b0011101010: data <= 9'h001; 
        10'b0011101011: data <= 9'h001; 
        10'b0011101100: data <= 9'h000; 
        10'b0011101101: data <= 9'h000; 
        10'b0011101110: data <= 9'h000; 
        10'b0011101111: data <= 9'h001; 
        10'b0011110000: data <= 9'h003; 
        10'b0011110001: data <= 9'h002; 
        10'b0011110010: data <= 9'h002; 
        10'b0011110011: data <= 9'h001; 
        10'b0011110100: data <= 9'h001; 
        10'b0011110101: data <= 9'h000; 
        10'b0011110110: data <= 9'h001; 
        10'b0011110111: data <= 9'h002; 
        10'b0011111000: data <= 9'h000; 
        10'b0011111001: data <= 9'h1ff; 
        10'b0011111010: data <= 9'h000; 
        10'b0011111011: data <= 9'h000; 
        10'b0011111100: data <= 9'h000; 
        10'b0011111101: data <= 9'h000; 
        10'b0011111110: data <= 9'h000; 
        10'b0011111111: data <= 9'h000; 
        10'b0100000000: data <= 9'h1ff; 
        10'b0100000001: data <= 9'h000; 
        10'b0100000010: data <= 9'h1ff; 
        10'b0100000011: data <= 9'h000; 
        10'b0100000100: data <= 9'h000; 
        10'b0100000101: data <= 9'h000; 
        10'b0100000110: data <= 9'h000; 
        10'b0100000111: data <= 9'h000; 
        10'b0100001000: data <= 9'h000; 
        10'b0100001001: data <= 9'h001; 
        10'b0100001010: data <= 9'h001; 
        10'b0100001011: data <= 9'h000; 
        10'b0100001100: data <= 9'h001; 
        10'b0100001101: data <= 9'h002; 
        10'b0100001110: data <= 9'h002; 
        10'b0100001111: data <= 9'h001; 
        10'b0100010000: data <= 9'h000; 
        10'b0100010001: data <= 9'h000; 
        10'b0100010010: data <= 9'h001; 
        10'b0100010011: data <= 9'h002; 
        10'b0100010100: data <= 9'h001; 
        10'b0100010101: data <= 9'h000; 
        10'b0100010110: data <= 9'h000; 
        10'b0100010111: data <= 9'h000; 
        10'b0100011000: data <= 9'h000; 
        10'b0100011001: data <= 9'h000; 
        10'b0100011010: data <= 9'h000; 
        10'b0100011011: data <= 9'h000; 
        10'b0100011100: data <= 9'h000; 
        10'b0100011101: data <= 9'h000; 
        10'b0100011110: data <= 9'h000; 
        10'b0100011111: data <= 9'h000; 
        10'b0100100000: data <= 9'h000; 
        10'b0100100001: data <= 9'h000; 
        10'b0100100010: data <= 9'h000; 
        10'b0100100011: data <= 9'h000; 
        10'b0100100100: data <= 9'h000; 
        10'b0100100101: data <= 9'h000; 
        10'b0100100110: data <= 9'h1ff; 
        10'b0100100111: data <= 9'h1ff; 
        10'b0100101000: data <= 9'h1ff; 
        10'b0100101001: data <= 9'h001; 
        10'b0100101010: data <= 9'h002; 
        10'b0100101011: data <= 9'h002; 
        10'b0100101100: data <= 9'h002; 
        10'b0100101101: data <= 9'h001; 
        10'b0100101110: data <= 9'h002; 
        10'b0100101111: data <= 9'h002; 
        10'b0100110000: data <= 9'h001; 
        10'b0100110001: data <= 9'h000; 
        10'b0100110010: data <= 9'h000; 
        10'b0100110011: data <= 9'h000; 
        10'b0100110100: data <= 9'h000; 
        10'b0100110101: data <= 9'h000; 
        10'b0100110110: data <= 9'h000; 
        10'b0100110111: data <= 9'h000; 
        10'b0100111000: data <= 9'h1ff; 
        10'b0100111001: data <= 9'h000; 
        10'b0100111010: data <= 9'h000; 
        10'b0100111011: data <= 9'h001; 
        10'b0100111100: data <= 9'h000; 
        10'b0100111101: data <= 9'h000; 
        10'b0100111110: data <= 9'h000; 
        10'b0100111111: data <= 9'h000; 
        10'b0101000000: data <= 9'h000; 
        10'b0101000001: data <= 9'h000; 
        10'b0101000010: data <= 9'h1fe; 
        10'b0101000011: data <= 9'h1fd; 
        10'b0101000100: data <= 9'h1fd; 
        10'b0101000101: data <= 9'h1ff; 
        10'b0101000110: data <= 9'h000; 
        10'b0101000111: data <= 9'h001; 
        10'b0101001000: data <= 9'h001; 
        10'b0101001001: data <= 9'h001; 
        10'b0101001010: data <= 9'h002; 
        10'b0101001011: data <= 9'h002; 
        10'b0101001100: data <= 9'h001; 
        10'b0101001101: data <= 9'h000; 
        10'b0101001110: data <= 9'h000; 
        10'b0101001111: data <= 9'h000; 
        10'b0101010000: data <= 9'h000; 
        10'b0101010001: data <= 9'h000; 
        10'b0101010010: data <= 9'h000; 
        10'b0101010011: data <= 9'h000; 
        10'b0101010100: data <= 9'h000; 
        10'b0101010101: data <= 9'h000; 
        10'b0101010110: data <= 9'h001; 
        10'b0101010111: data <= 9'h001; 
        10'b0101011000: data <= 9'h000; 
        10'b0101011001: data <= 9'h000; 
        10'b0101011010: data <= 9'h001; 
        10'b0101011011: data <= 9'h000; 
        10'b0101011100: data <= 9'h001; 
        10'b0101011101: data <= 9'h1ff; 
        10'b0101011110: data <= 9'h1fc; 
        10'b0101011111: data <= 9'h1fc; 
        10'b0101100000: data <= 9'h1fc; 
        10'b0101100001: data <= 9'h1fe; 
        10'b0101100010: data <= 9'h000; 
        10'b0101100011: data <= 9'h000; 
        10'b0101100100: data <= 9'h000; 
        10'b0101100101: data <= 9'h001; 
        10'b0101100110: data <= 9'h002; 
        10'b0101100111: data <= 9'h002; 
        10'b0101101000: data <= 9'h002; 
        10'b0101101001: data <= 9'h000; 
        10'b0101101010: data <= 9'h000; 
        10'b0101101011: data <= 9'h000; 
        10'b0101101100: data <= 9'h000; 
        10'b0101101101: data <= 9'h000; 
        10'b0101101110: data <= 9'h000; 
        10'b0101101111: data <= 9'h000; 
        10'b0101110000: data <= 9'h000; 
        10'b0101110001: data <= 9'h000; 
        10'b0101110010: data <= 9'h001; 
        10'b0101110011: data <= 9'h001; 
        10'b0101110100: data <= 9'h001; 
        10'b0101110101: data <= 9'h001; 
        10'b0101110110: data <= 9'h001; 
        10'b0101110111: data <= 9'h001; 
        10'b0101111000: data <= 9'h000; 
        10'b0101111001: data <= 9'h1fe; 
        10'b0101111010: data <= 9'h1fc; 
        10'b0101111011: data <= 9'h1fb; 
        10'b0101111100: data <= 9'h1fc; 
        10'b0101111101: data <= 9'h1fe; 
        10'b0101111110: data <= 9'h1ff; 
        10'b0101111111: data <= 9'h1ff; 
        10'b0110000000: data <= 9'h1ff; 
        10'b0110000001: data <= 9'h000; 
        10'b0110000010: data <= 9'h002; 
        10'b0110000011: data <= 9'h002; 
        10'b0110000100: data <= 9'h001; 
        10'b0110000101: data <= 9'h000; 
        10'b0110000110: data <= 9'h000; 
        10'b0110000111: data <= 9'h000; 
        10'b0110001000: data <= 9'h000; 
        10'b0110001001: data <= 9'h000; 
        10'b0110001010: data <= 9'h000; 
        10'b0110001011: data <= 9'h000; 
        10'b0110001100: data <= 9'h000; 
        10'b0110001101: data <= 9'h001; 
        10'b0110001110: data <= 9'h001; 
        10'b0110001111: data <= 9'h002; 
        10'b0110010000: data <= 9'h001; 
        10'b0110010001: data <= 9'h001; 
        10'b0110010010: data <= 9'h002; 
        10'b0110010011: data <= 9'h001; 
        10'b0110010100: data <= 9'h000; 
        10'b0110010101: data <= 9'h1fe; 
        10'b0110010110: data <= 9'h1fc; 
        10'b0110010111: data <= 9'h1fb; 
        10'b0110011000: data <= 9'h1fc; 
        10'b0110011001: data <= 9'h1fe; 
        10'b0110011010: data <= 9'h1ff; 
        10'b0110011011: data <= 9'h1ff; 
        10'b0110011100: data <= 9'h000; 
        10'b0110011101: data <= 9'h001; 
        10'b0110011110: data <= 9'h001; 
        10'b0110011111: data <= 9'h002; 
        10'b0110100000: data <= 9'h001; 
        10'b0110100001: data <= 9'h000; 
        10'b0110100010: data <= 9'h000; 
        10'b0110100011: data <= 9'h000; 
        10'b0110100100: data <= 9'h000; 
        10'b0110100101: data <= 9'h000; 
        10'b0110100110: data <= 9'h000; 
        10'b0110100111: data <= 9'h000; 
        10'b0110101000: data <= 9'h000; 
        10'b0110101001: data <= 9'h002; 
        10'b0110101010: data <= 9'h001; 
        10'b0110101011: data <= 9'h002; 
        10'b0110101100: data <= 9'h001; 
        10'b0110101101: data <= 9'h001; 
        10'b0110101110: data <= 9'h002; 
        10'b0110101111: data <= 9'h001; 
        10'b0110110000: data <= 9'h1ff; 
        10'b0110110001: data <= 9'h1fc; 
        10'b0110110010: data <= 9'h1fb; 
        10'b0110110011: data <= 9'h1fb; 
        10'b0110110100: data <= 9'h1fd; 
        10'b0110110101: data <= 9'h1fe; 
        10'b0110110110: data <= 9'h1ff; 
        10'b0110110111: data <= 9'h1ff; 
        10'b0110111000: data <= 9'h000; 
        10'b0110111001: data <= 9'h000; 
        10'b0110111010: data <= 9'h002; 
        10'b0110111011: data <= 9'h002; 
        10'b0110111100: data <= 9'h001; 
        10'b0110111101: data <= 9'h000; 
        10'b0110111110: data <= 9'h000; 
        10'b0110111111: data <= 9'h000; 
        10'b0111000000: data <= 9'h000; 
        10'b0111000001: data <= 9'h000; 
        10'b0111000010: data <= 9'h000; 
        10'b0111000011: data <= 9'h000; 
        10'b0111000100: data <= 9'h000; 
        10'b0111000101: data <= 9'h001; 
        10'b0111000110: data <= 9'h002; 
        10'b0111000111: data <= 9'h001; 
        10'b0111001000: data <= 9'h001; 
        10'b0111001001: data <= 9'h001; 
        10'b0111001010: data <= 9'h002; 
        10'b0111001011: data <= 9'h000; 
        10'b0111001100: data <= 9'h1fd; 
        10'b0111001101: data <= 9'h1fb; 
        10'b0111001110: data <= 9'h1fb; 
        10'b0111001111: data <= 9'h1fc; 
        10'b0111010000: data <= 9'h1fe; 
        10'b0111010001: data <= 9'h1ff; 
        10'b0111010010: data <= 9'h000; 
        10'b0111010011: data <= 9'h000; 
        10'b0111010100: data <= 9'h001; 
        10'b0111010101: data <= 9'h001; 
        10'b0111010110: data <= 9'h001; 
        10'b0111010111: data <= 9'h001; 
        10'b0111011000: data <= 9'h001; 
        10'b0111011001: data <= 9'h000; 
        10'b0111011010: data <= 9'h000; 
        10'b0111011011: data <= 9'h000; 
        10'b0111011100: data <= 9'h000; 
        10'b0111011101: data <= 9'h000; 
        10'b0111011110: data <= 9'h000; 
        10'b0111011111: data <= 9'h1ff; 
        10'b0111100000: data <= 9'h000; 
        10'b0111100001: data <= 9'h001; 
        10'b0111100010: data <= 9'h001; 
        10'b0111100011: data <= 9'h001; 
        10'b0111100100: data <= 9'h000; 
        10'b0111100101: data <= 9'h001; 
        10'b0111100110: data <= 9'h002; 
        10'b0111100111: data <= 9'h000; 
        10'b0111101000: data <= 9'h1fd; 
        10'b0111101001: data <= 9'h1fb; 
        10'b0111101010: data <= 9'h1fc; 
        10'b0111101011: data <= 9'h1fe; 
        10'b0111101100: data <= 9'h000; 
        10'b0111101101: data <= 9'h001; 
        10'b0111101110: data <= 9'h001; 
        10'b0111101111: data <= 9'h001; 
        10'b0111110000: data <= 9'h001; 
        10'b0111110001: data <= 9'h001; 
        10'b0111110010: data <= 9'h001; 
        10'b0111110011: data <= 9'h001; 
        10'b0111110100: data <= 9'h000; 
        10'b0111110101: data <= 9'h000; 
        10'b0111110110: data <= 9'h000; 
        10'b0111110111: data <= 9'h000; 
        10'b0111111000: data <= 9'h000; 
        10'b0111111001: data <= 9'h000; 
        10'b0111111010: data <= 9'h000; 
        10'b0111111011: data <= 9'h000; 
        10'b0111111100: data <= 9'h000; 
        10'b0111111101: data <= 9'h001; 
        10'b0111111110: data <= 9'h001; 
        10'b0111111111: data <= 9'h001; 
        10'b1000000000: data <= 9'h000; 
        10'b1000000001: data <= 9'h001; 
        10'b1000000010: data <= 9'h003; 
        10'b1000000011: data <= 9'h000; 
        10'b1000000100: data <= 9'h1fe; 
        10'b1000000101: data <= 9'h1fd; 
        10'b1000000110: data <= 9'h1fe; 
        10'b1000000111: data <= 9'h1ff; 
        10'b1000001000: data <= 9'h001; 
        10'b1000001001: data <= 9'h001; 
        10'b1000001010: data <= 9'h001; 
        10'b1000001011: data <= 9'h000; 
        10'b1000001100: data <= 9'h000; 
        10'b1000001101: data <= 9'h000; 
        10'b1000001110: data <= 9'h001; 
        10'b1000001111: data <= 9'h000; 
        10'b1000010000: data <= 9'h000; 
        10'b1000010001: data <= 9'h000; 
        10'b1000010010: data <= 9'h000; 
        10'b1000010011: data <= 9'h000; 
        10'b1000010100: data <= 9'h000; 
        10'b1000010101: data <= 9'h000; 
        10'b1000010110: data <= 9'h000; 
        10'b1000010111: data <= 9'h1ff; 
        10'b1000011000: data <= 9'h000; 
        10'b1000011001: data <= 9'h001; 
        10'b1000011010: data <= 9'h002; 
        10'b1000011011: data <= 9'h002; 
        10'b1000011100: data <= 9'h001; 
        10'b1000011101: data <= 9'h002; 
        10'b1000011110: data <= 9'h003; 
        10'b1000011111: data <= 9'h002; 
        10'b1000100000: data <= 9'h000; 
        10'b1000100001: data <= 9'h1ff; 
        10'b1000100010: data <= 9'h000; 
        10'b1000100011: data <= 9'h000; 
        10'b1000100100: data <= 9'h000; 
        10'b1000100101: data <= 9'h000; 
        10'b1000100110: data <= 9'h000; 
        10'b1000100111: data <= 9'h000; 
        10'b1000101000: data <= 9'h000; 
        10'b1000101001: data <= 9'h000; 
        10'b1000101010: data <= 9'h001; 
        10'b1000101011: data <= 9'h000; 
        10'b1000101100: data <= 9'h000; 
        10'b1000101101: data <= 9'h000; 
        10'b1000101110: data <= 9'h000; 
        10'b1000101111: data <= 9'h000; 
        10'b1000110000: data <= 9'h000; 
        10'b1000110001: data <= 9'h000; 
        10'b1000110010: data <= 9'h000; 
        10'b1000110011: data <= 9'h000; 
        10'b1000110100: data <= 9'h000; 
        10'b1000110101: data <= 9'h001; 
        10'b1000110110: data <= 9'h001; 
        10'b1000110111: data <= 9'h001; 
        10'b1000111000: data <= 9'h001; 
        10'b1000111001: data <= 9'h002; 
        10'b1000111010: data <= 9'h002; 
        10'b1000111011: data <= 9'h002; 
        10'b1000111100: data <= 9'h001; 
        10'b1000111101: data <= 9'h000; 
        10'b1000111110: data <= 9'h000; 
        10'b1000111111: data <= 9'h000; 
        10'b1001000000: data <= 9'h000; 
        10'b1001000001: data <= 9'h000; 
        10'b1001000010: data <= 9'h000; 
        10'b1001000011: data <= 9'h000; 
        10'b1001000100: data <= 9'h000; 
        10'b1001000101: data <= 9'h000; 
        10'b1001000110: data <= 9'h000; 
        10'b1001000111: data <= 9'h000; 
        10'b1001001000: data <= 9'h000; 
        10'b1001001001: data <= 9'h000; 
        10'b1001001010: data <= 9'h000; 
        10'b1001001011: data <= 9'h000; 
        10'b1001001100: data <= 9'h000; 
        10'b1001001101: data <= 9'h000; 
        10'b1001001110: data <= 9'h000; 
        10'b1001001111: data <= 9'h000; 
        10'b1001010000: data <= 9'h000; 
        10'b1001010001: data <= 9'h000; 
        10'b1001010010: data <= 9'h001; 
        10'b1001010011: data <= 9'h001; 
        10'b1001010100: data <= 9'h001; 
        10'b1001010101: data <= 9'h001; 
        10'b1001010110: data <= 9'h002; 
        10'b1001010111: data <= 9'h002; 
        10'b1001011000: data <= 9'h002; 
        10'b1001011001: data <= 9'h001; 
        10'b1001011010: data <= 9'h000; 
        10'b1001011011: data <= 9'h000; 
        10'b1001011100: data <= 9'h000; 
        10'b1001011101: data <= 9'h1ff; 
        10'b1001011110: data <= 9'h000; 
        10'b1001011111: data <= 9'h000; 
        10'b1001100000: data <= 9'h000; 
        10'b1001100001: data <= 9'h000; 
        10'b1001100010: data <= 9'h000; 
        10'b1001100011: data <= 9'h000; 
        10'b1001100100: data <= 9'h000; 
        10'b1001100101: data <= 9'h000; 
        10'b1001100110: data <= 9'h000; 
        10'b1001100111: data <= 9'h000; 
        10'b1001101000: data <= 9'h000; 
        10'b1001101001: data <= 9'h000; 
        10'b1001101010: data <= 9'h000; 
        10'b1001101011: data <= 9'h000; 
        10'b1001101100: data <= 9'h000; 
        10'b1001101101: data <= 9'h000; 
        10'b1001101110: data <= 9'h001; 
        10'b1001101111: data <= 9'h001; 
        10'b1001110000: data <= 9'h002; 
        10'b1001110001: data <= 9'h001; 
        10'b1001110010: data <= 9'h001; 
        10'b1001110011: data <= 9'h002; 
        10'b1001110100: data <= 9'h001; 
        10'b1001110101: data <= 9'h002; 
        10'b1001110110: data <= 9'h001; 
        10'b1001110111: data <= 9'h001; 
        10'b1001111000: data <= 9'h000; 
        10'b1001111001: data <= 9'h000; 
        10'b1001111010: data <= 9'h000; 
        10'b1001111011: data <= 9'h000; 
        10'b1001111100: data <= 9'h000; 
        10'b1001111101: data <= 9'h000; 
        10'b1001111110: data <= 9'h000; 
        10'b1001111111: data <= 9'h000; 
        10'b1010000000: data <= 9'h000; 
        10'b1010000001: data <= 9'h000; 
        10'b1010000010: data <= 9'h000; 
        10'b1010000011: data <= 9'h000; 
        10'b1010000100: data <= 9'h000; 
        10'b1010000101: data <= 9'h000; 
        10'b1010000110: data <= 9'h000; 
        10'b1010000111: data <= 9'h000; 
        10'b1010001000: data <= 9'h000; 
        10'b1010001001: data <= 9'h000; 
        10'b1010001010: data <= 9'h000; 
        10'b1010001011: data <= 9'h000; 
        10'b1010001100: data <= 9'h001; 
        10'b1010001101: data <= 9'h001; 
        10'b1010001110: data <= 9'h002; 
        10'b1010001111: data <= 9'h002; 
        10'b1010010000: data <= 9'h002; 
        10'b1010010001: data <= 9'h001; 
        10'b1010010010: data <= 9'h001; 
        10'b1010010011: data <= 9'h001; 
        10'b1010010100: data <= 9'h000; 
        10'b1010010101: data <= 9'h000; 
        10'b1010010110: data <= 9'h1ff; 
        10'b1010010111: data <= 9'h1ff; 
        10'b1010011000: data <= 9'h1ff; 
        10'b1010011001: data <= 9'h000; 
        10'b1010011010: data <= 9'h000; 
        10'b1010011011: data <= 9'h000; 
        10'b1010011100: data <= 9'h000; 
        10'b1010011101: data <= 9'h000; 
        10'b1010011110: data <= 9'h000; 
        10'b1010011111: data <= 9'h000; 
        10'b1010100000: data <= 9'h000; 
        10'b1010100001: data <= 9'h000; 
        10'b1010100010: data <= 9'h000; 
        10'b1010100011: data <= 9'h000; 
        10'b1010100100: data <= 9'h000; 
        10'b1010100101: data <= 9'h000; 
        10'b1010100110: data <= 9'h000; 
        10'b1010100111: data <= 9'h1ff; 
        10'b1010101000: data <= 9'h000; 
        10'b1010101001: data <= 9'h000; 
        10'b1010101010: data <= 9'h000; 
        10'b1010101011: data <= 9'h000; 
        10'b1010101100: data <= 9'h001; 
        10'b1010101101: data <= 9'h001; 
        10'b1010101110: data <= 9'h000; 
        10'b1010101111: data <= 9'h000; 
        10'b1010110000: data <= 9'h1ff; 
        10'b1010110001: data <= 9'h1ff; 
        10'b1010110010: data <= 9'h1ff; 
        10'b1010110011: data <= 9'h1ff; 
        10'b1010110100: data <= 9'h1ff; 
        10'b1010110101: data <= 9'h1ff; 
        10'b1010110110: data <= 9'h000; 
        10'b1010110111: data <= 9'h000; 
        10'b1010111000: data <= 9'h000; 
        10'b1010111001: data <= 9'h000; 
        10'b1010111010: data <= 9'h000; 
        10'b1010111011: data <= 9'h000; 
        10'b1010111100: data <= 9'h000; 
        10'b1010111101: data <= 9'h000; 
        10'b1010111110: data <= 9'h000; 
        10'b1010111111: data <= 9'h000; 
        10'b1011000000: data <= 9'h000; 
        10'b1011000001: data <= 9'h000; 
        10'b1011000010: data <= 9'h000; 
        10'b1011000011: data <= 9'h000; 
        10'b1011000100: data <= 9'h1ff; 
        10'b1011000101: data <= 9'h1ff; 
        10'b1011000110: data <= 9'h1ff; 
        10'b1011000111: data <= 9'h1ff; 
        10'b1011001000: data <= 9'h1ff; 
        10'b1011001001: data <= 9'h1ff; 
        10'b1011001010: data <= 9'h1ff; 
        10'b1011001011: data <= 9'h1ff; 
        10'b1011001100: data <= 9'h1ff; 
        10'b1011001101: data <= 9'h1ff; 
        10'b1011001110: data <= 9'h1ff; 
        10'b1011001111: data <= 9'h000; 
        10'b1011010000: data <= 9'h1ff; 
        10'b1011010001: data <= 9'h000; 
        10'b1011010010: data <= 9'h000; 
        10'b1011010011: data <= 9'h000; 
        10'b1011010100: data <= 9'h000; 
        10'b1011010101: data <= 9'h000; 
        10'b1011010110: data <= 9'h000; 
        10'b1011010111: data <= 9'h000; 
        10'b1011011000: data <= 9'h000; 
        10'b1011011001: data <= 9'h000; 
        10'b1011011010: data <= 9'h000; 
        10'b1011011011: data <= 9'h000; 
        10'b1011011100: data <= 9'h000; 
        10'b1011011101: data <= 9'h000; 
        10'b1011011110: data <= 9'h000; 
        10'b1011011111: data <= 9'h000; 
        10'b1011100000: data <= 9'h000; 
        10'b1011100001: data <= 9'h1ff; 
        10'b1011100010: data <= 9'h1ff; 
        10'b1011100011: data <= 9'h1ff; 
        10'b1011100100: data <= 9'h000; 
        10'b1011100101: data <= 9'h1ff; 
        10'b1011100110: data <= 9'h1ff; 
        10'b1011100111: data <= 9'h000; 
        10'b1011101000: data <= 9'h1ff; 
        10'b1011101001: data <= 9'h000; 
        10'b1011101010: data <= 9'h000; 
        10'b1011101011: data <= 9'h000; 
        10'b1011101100: data <= 9'h000; 
        10'b1011101101: data <= 9'h1ff; 
        10'b1011101110: data <= 9'h000; 
        10'b1011101111: data <= 9'h000; 
        10'b1011110000: data <= 9'h000; 
        10'b1011110001: data <= 9'h000; 
        10'b1011110010: data <= 9'h000; 
        10'b1011110011: data <= 9'h000; 
        10'b1011110100: data <= 9'h000; 
        10'b1011110101: data <= 9'h000; 
        10'b1011110110: data <= 9'h000; 
        10'b1011110111: data <= 9'h000; 
        10'b1011111000: data <= 9'h000; 
        10'b1011111001: data <= 9'h000; 
        10'b1011111010: data <= 9'h000; 
        10'b1011111011: data <= 9'h000; 
        10'b1011111100: data <= 9'h000; 
        10'b1011111101: data <= 9'h000; 
        10'b1011111110: data <= 9'h000; 
        10'b1011111111: data <= 9'h000; 
        10'b1100000000: data <= 9'h000; 
        10'b1100000001: data <= 9'h000; 
        10'b1100000010: data <= 9'h000; 
        10'b1100000011: data <= 9'h000; 
        10'b1100000100: data <= 9'h000; 
        10'b1100000101: data <= 9'h000; 
        10'b1100000110: data <= 9'h000; 
        10'b1100000111: data <= 9'h000; 
        10'b1100001000: data <= 9'h000; 
        10'b1100001001: data <= 9'h000; 
        10'b1100001010: data <= 9'h000; 
        10'b1100001011: data <= 9'h000; 
        10'b1100001100: data <= 9'h000; 
        10'b1100001101: data <= 9'h000; 
        10'b1100001110: data <= 9'h000; 
        10'b1100001111: data <= 9'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 4) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 10'h3ff; 
        10'b0000000001: data <= 10'h000; 
        10'b0000000010: data <= 10'h000; 
        10'b0000000011: data <= 10'h000; 
        10'b0000000100: data <= 10'h000; 
        10'b0000000101: data <= 10'h000; 
        10'b0000000110: data <= 10'h000; 
        10'b0000000111: data <= 10'h000; 
        10'b0000001000: data <= 10'h000; 
        10'b0000001001: data <= 10'h000; 
        10'b0000001010: data <= 10'h000; 
        10'b0000001011: data <= 10'h000; 
        10'b0000001100: data <= 10'h000; 
        10'b0000001101: data <= 10'h3ff; 
        10'b0000001110: data <= 10'h000; 
        10'b0000001111: data <= 10'h3ff; 
        10'b0000010000: data <= 10'h3ff; 
        10'b0000010001: data <= 10'h000; 
        10'b0000010010: data <= 10'h3ff; 
        10'b0000010011: data <= 10'h000; 
        10'b0000010100: data <= 10'h3ff; 
        10'b0000010101: data <= 10'h000; 
        10'b0000010110: data <= 10'h3ff; 
        10'b0000010111: data <= 10'h000; 
        10'b0000011000: data <= 10'h000; 
        10'b0000011001: data <= 10'h000; 
        10'b0000011010: data <= 10'h000; 
        10'b0000011011: data <= 10'h000; 
        10'b0000011100: data <= 10'h000; 
        10'b0000011101: data <= 10'h000; 
        10'b0000011110: data <= 10'h000; 
        10'b0000011111: data <= 10'h3ff; 
        10'b0000100000: data <= 10'h3ff; 
        10'b0000100001: data <= 10'h000; 
        10'b0000100010: data <= 10'h3ff; 
        10'b0000100011: data <= 10'h000; 
        10'b0000100100: data <= 10'h000; 
        10'b0000100101: data <= 10'h3ff; 
        10'b0000100110: data <= 10'h000; 
        10'b0000100111: data <= 10'h000; 
        10'b0000101000: data <= 10'h000; 
        10'b0000101001: data <= 10'h3ff; 
        10'b0000101010: data <= 10'h000; 
        10'b0000101011: data <= 10'h000; 
        10'b0000101100: data <= 10'h000; 
        10'b0000101101: data <= 10'h3ff; 
        10'b0000101110: data <= 10'h000; 
        10'b0000101111: data <= 10'h000; 
        10'b0000110000: data <= 10'h3ff; 
        10'b0000110001: data <= 10'h000; 
        10'b0000110010: data <= 10'h000; 
        10'b0000110011: data <= 10'h3ff; 
        10'b0000110100: data <= 10'h000; 
        10'b0000110101: data <= 10'h000; 
        10'b0000110110: data <= 10'h000; 
        10'b0000110111: data <= 10'h000; 
        10'b0000111000: data <= 10'h3ff; 
        10'b0000111001: data <= 10'h000; 
        10'b0000111010: data <= 10'h000; 
        10'b0000111011: data <= 10'h000; 
        10'b0000111100: data <= 10'h000; 
        10'b0000111101: data <= 10'h3ff; 
        10'b0000111110: data <= 10'h000; 
        10'b0000111111: data <= 10'h000; 
        10'b0001000000: data <= 10'h000; 
        10'b0001000001: data <= 10'h000; 
        10'b0001000010: data <= 10'h000; 
        10'b0001000011: data <= 10'h3ff; 
        10'b0001000100: data <= 10'h3ff; 
        10'b0001000101: data <= 10'h000; 
        10'b0001000110: data <= 10'h3ff; 
        10'b0001000111: data <= 10'h3ff; 
        10'b0001001000: data <= 10'h3ff; 
        10'b0001001001: data <= 10'h000; 
        10'b0001001010: data <= 10'h3ff; 
        10'b0001001011: data <= 10'h3ff; 
        10'b0001001100: data <= 10'h000; 
        10'b0001001101: data <= 10'h000; 
        10'b0001001110: data <= 10'h000; 
        10'b0001001111: data <= 10'h000; 
        10'b0001010000: data <= 10'h000; 
        10'b0001010001: data <= 10'h3ff; 
        10'b0001010010: data <= 10'h000; 
        10'b0001010011: data <= 10'h000; 
        10'b0001010100: data <= 10'h3ff; 
        10'b0001010101: data <= 10'h000; 
        10'b0001010110: data <= 10'h000; 
        10'b0001010111: data <= 10'h3ff; 
        10'b0001011000: data <= 10'h000; 
        10'b0001011001: data <= 10'h000; 
        10'b0001011010: data <= 10'h000; 
        10'b0001011011: data <= 10'h000; 
        10'b0001011100: data <= 10'h000; 
        10'b0001011101: data <= 10'h000; 
        10'b0001011110: data <= 10'h000; 
        10'b0001011111: data <= 10'h3ff; 
        10'b0001100000: data <= 10'h3ff; 
        10'b0001100001: data <= 10'h3ff; 
        10'b0001100010: data <= 10'h3ff; 
        10'b0001100011: data <= 10'h3ff; 
        10'b0001100100: data <= 10'h000; 
        10'b0001100101: data <= 10'h000; 
        10'b0001100110: data <= 10'h3ff; 
        10'b0001100111: data <= 10'h3ff; 
        10'b0001101000: data <= 10'h3ff; 
        10'b0001101001: data <= 10'h3ff; 
        10'b0001101010: data <= 10'h3ff; 
        10'b0001101011: data <= 10'h3ff; 
        10'b0001101100: data <= 10'h3ff; 
        10'b0001101101: data <= 10'h000; 
        10'b0001101110: data <= 10'h000; 
        10'b0001101111: data <= 10'h000; 
        10'b0001110000: data <= 10'h000; 
        10'b0001110001: data <= 10'h3ff; 
        10'b0001110010: data <= 10'h000; 
        10'b0001110011: data <= 10'h3ff; 
        10'b0001110100: data <= 10'h3ff; 
        10'b0001110101: data <= 10'h000; 
        10'b0001110110: data <= 10'h000; 
        10'b0001110111: data <= 10'h3ff; 
        10'b0001111000: data <= 10'h000; 
        10'b0001111001: data <= 10'h000; 
        10'b0001111010: data <= 10'h3ff; 
        10'b0001111011: data <= 10'h3ff; 
        10'b0001111100: data <= 10'h3ff; 
        10'b0001111101: data <= 10'h3ff; 
        10'b0001111110: data <= 10'h000; 
        10'b0001111111: data <= 10'h000; 
        10'b0010000000: data <= 10'h3ff; 
        10'b0010000001: data <= 10'h3ff; 
        10'b0010000010: data <= 10'h3ff; 
        10'b0010000011: data <= 10'h3ff; 
        10'b0010000100: data <= 10'h000; 
        10'b0010000101: data <= 10'h3ff; 
        10'b0010000110: data <= 10'h3ff; 
        10'b0010000111: data <= 10'h000; 
        10'b0010001000: data <= 10'h3ff; 
        10'b0010001001: data <= 10'h000; 
        10'b0010001010: data <= 10'h000; 
        10'b0010001011: data <= 10'h000; 
        10'b0010001100: data <= 10'h000; 
        10'b0010001101: data <= 10'h000; 
        10'b0010001110: data <= 10'h000; 
        10'b0010001111: data <= 10'h3ff; 
        10'b0010010000: data <= 10'h000; 
        10'b0010010001: data <= 10'h000; 
        10'b0010010010: data <= 10'h000; 
        10'b0010010011: data <= 10'h000; 
        10'b0010010100: data <= 10'h000; 
        10'b0010010101: data <= 10'h3ff; 
        10'b0010010110: data <= 10'h000; 
        10'b0010010111: data <= 10'h000; 
        10'b0010011000: data <= 10'h001; 
        10'b0010011001: data <= 10'h002; 
        10'b0010011010: data <= 10'h002; 
        10'b0010011011: data <= 10'h002; 
        10'b0010011100: data <= 10'h003; 
        10'b0010011101: data <= 10'h003; 
        10'b0010011110: data <= 10'h003; 
        10'b0010011111: data <= 10'h001; 
        10'b0010100000: data <= 10'h000; 
        10'b0010100001: data <= 10'h001; 
        10'b0010100010: data <= 10'h000; 
        10'b0010100011: data <= 10'h000; 
        10'b0010100100: data <= 10'h3ff; 
        10'b0010100101: data <= 10'h3ff; 
        10'b0010100110: data <= 10'h000; 
        10'b0010100111: data <= 10'h3ff; 
        10'b0010101000: data <= 10'h000; 
        10'b0010101001: data <= 10'h000; 
        10'b0010101010: data <= 10'h000; 
        10'b0010101011: data <= 10'h000; 
        10'b0010101100: data <= 10'h000; 
        10'b0010101101: data <= 10'h000; 
        10'b0010101110: data <= 10'h000; 
        10'b0010101111: data <= 10'h000; 
        10'b0010110000: data <= 10'h3ff; 
        10'b0010110001: data <= 10'h3ff; 
        10'b0010110010: data <= 10'h001; 
        10'b0010110011: data <= 10'h000; 
        10'b0010110100: data <= 10'h002; 
        10'b0010110101: data <= 10'h001; 
        10'b0010110110: data <= 10'h001; 
        10'b0010110111: data <= 10'h002; 
        10'b0010111000: data <= 10'h003; 
        10'b0010111001: data <= 10'h004; 
        10'b0010111010: data <= 10'h003; 
        10'b0010111011: data <= 10'h003; 
        10'b0010111100: data <= 10'h003; 
        10'b0010111101: data <= 10'h003; 
        10'b0010111110: data <= 10'h002; 
        10'b0010111111: data <= 10'h001; 
        10'b0011000000: data <= 10'h3ff; 
        10'b0011000001: data <= 10'h3ff; 
        10'b0011000010: data <= 10'h3ff; 
        10'b0011000011: data <= 10'h000; 
        10'b0011000100: data <= 10'h000; 
        10'b0011000101: data <= 10'h000; 
        10'b0011000110: data <= 10'h000; 
        10'b0011000111: data <= 10'h3ff; 
        10'b0011001000: data <= 10'h3ff; 
        10'b0011001001: data <= 10'h000; 
        10'b0011001010: data <= 10'h3ff; 
        10'b0011001011: data <= 10'h000; 
        10'b0011001100: data <= 10'h3ff; 
        10'b0011001101: data <= 10'h000; 
        10'b0011001110: data <= 10'h000; 
        10'b0011001111: data <= 10'h001; 
        10'b0011010000: data <= 10'h003; 
        10'b0011010001: data <= 10'h002; 
        10'b0011010010: data <= 10'h001; 
        10'b0011010011: data <= 10'h001; 
        10'b0011010100: data <= 10'h002; 
        10'b0011010101: data <= 10'h004; 
        10'b0011010110: data <= 10'h003; 
        10'b0011010111: data <= 10'h003; 
        10'b0011011000: data <= 10'h001; 
        10'b0011011001: data <= 10'h002; 
        10'b0011011010: data <= 10'h002; 
        10'b0011011011: data <= 10'h001; 
        10'b0011011100: data <= 10'h3ff; 
        10'b0011011101: data <= 10'h3ff; 
        10'b0011011110: data <= 10'h3ff; 
        10'b0011011111: data <= 10'h000; 
        10'b0011100000: data <= 10'h000; 
        10'b0011100001: data <= 10'h000; 
        10'b0011100010: data <= 10'h000; 
        10'b0011100011: data <= 10'h000; 
        10'b0011100100: data <= 10'h3ff; 
        10'b0011100101: data <= 10'h3ff; 
        10'b0011100110: data <= 10'h3ff; 
        10'b0011100111: data <= 10'h3ff; 
        10'b0011101000: data <= 10'h000; 
        10'b0011101001: data <= 10'h000; 
        10'b0011101010: data <= 10'h001; 
        10'b0011101011: data <= 10'h001; 
        10'b0011101100: data <= 10'h001; 
        10'b0011101101: data <= 10'h000; 
        10'b0011101110: data <= 10'h000; 
        10'b0011101111: data <= 10'h002; 
        10'b0011110000: data <= 10'h005; 
        10'b0011110001: data <= 10'h004; 
        10'b0011110010: data <= 10'h004; 
        10'b0011110011: data <= 10'h001; 
        10'b0011110100: data <= 10'h001; 
        10'b0011110101: data <= 10'h001; 
        10'b0011110110: data <= 10'h002; 
        10'b0011110111: data <= 10'h004; 
        10'b0011111000: data <= 10'h000; 
        10'b0011111001: data <= 10'h3ff; 
        10'b0011111010: data <= 10'h000; 
        10'b0011111011: data <= 10'h3ff; 
        10'b0011111100: data <= 10'h000; 
        10'b0011111101: data <= 10'h000; 
        10'b0011111110: data <= 10'h000; 
        10'b0011111111: data <= 10'h000; 
        10'b0100000000: data <= 10'h3ff; 
        10'b0100000001: data <= 10'h3ff; 
        10'b0100000010: data <= 10'h3ff; 
        10'b0100000011: data <= 10'h3ff; 
        10'b0100000100: data <= 10'h3ff; 
        10'b0100000101: data <= 10'h000; 
        10'b0100000110: data <= 10'h001; 
        10'b0100000111: data <= 10'h3ff; 
        10'b0100001000: data <= 10'h000; 
        10'b0100001001: data <= 10'h001; 
        10'b0100001010: data <= 10'h001; 
        10'b0100001011: data <= 10'h001; 
        10'b0100001100: data <= 10'h003; 
        10'b0100001101: data <= 10'h004; 
        10'b0100001110: data <= 10'h004; 
        10'b0100001111: data <= 10'h003; 
        10'b0100010000: data <= 10'h001; 
        10'b0100010001: data <= 10'h000; 
        10'b0100010010: data <= 10'h002; 
        10'b0100010011: data <= 10'h004; 
        10'b0100010100: data <= 10'h001; 
        10'b0100010101: data <= 10'h3ff; 
        10'b0100010110: data <= 10'h000; 
        10'b0100010111: data <= 10'h000; 
        10'b0100011000: data <= 10'h3ff; 
        10'b0100011001: data <= 10'h000; 
        10'b0100011010: data <= 10'h3ff; 
        10'b0100011011: data <= 10'h3ff; 
        10'b0100011100: data <= 10'h3ff; 
        10'b0100011101: data <= 10'h3ff; 
        10'b0100011110: data <= 10'h3ff; 
        10'b0100011111: data <= 10'h000; 
        10'b0100100000: data <= 10'h000; 
        10'b0100100001: data <= 10'h000; 
        10'b0100100010: data <= 10'h3ff; 
        10'b0100100011: data <= 10'h000; 
        10'b0100100100: data <= 10'h000; 
        10'b0100100101: data <= 10'h000; 
        10'b0100100110: data <= 10'h3ff; 
        10'b0100100111: data <= 10'h3fe; 
        10'b0100101000: data <= 10'h3ff; 
        10'b0100101001: data <= 10'h001; 
        10'b0100101010: data <= 10'h003; 
        10'b0100101011: data <= 10'h004; 
        10'b0100101100: data <= 10'h003; 
        10'b0100101101: data <= 10'h002; 
        10'b0100101110: data <= 10'h003; 
        10'b0100101111: data <= 10'h005; 
        10'b0100110000: data <= 10'h002; 
        10'b0100110001: data <= 10'h3ff; 
        10'b0100110010: data <= 10'h3ff; 
        10'b0100110011: data <= 10'h3ff; 
        10'b0100110100: data <= 10'h000; 
        10'b0100110101: data <= 10'h3ff; 
        10'b0100110110: data <= 10'h000; 
        10'b0100110111: data <= 10'h000; 
        10'b0100111000: data <= 10'h3fe; 
        10'b0100111001: data <= 10'h000; 
        10'b0100111010: data <= 10'h000; 
        10'b0100111011: data <= 10'h001; 
        10'b0100111100: data <= 10'h001; 
        10'b0100111101: data <= 10'h000; 
        10'b0100111110: data <= 10'h000; 
        10'b0100111111: data <= 10'h000; 
        10'b0101000000: data <= 10'h001; 
        10'b0101000001: data <= 10'h000; 
        10'b0101000010: data <= 10'h3fc; 
        10'b0101000011: data <= 10'h3f9; 
        10'b0101000100: data <= 10'h3fa; 
        10'b0101000101: data <= 10'h3fd; 
        10'b0101000110: data <= 10'h000; 
        10'b0101000111: data <= 10'h002; 
        10'b0101001000: data <= 10'h003; 
        10'b0101001001: data <= 10'h003; 
        10'b0101001010: data <= 10'h004; 
        10'b0101001011: data <= 10'h004; 
        10'b0101001100: data <= 10'h003; 
        10'b0101001101: data <= 10'h3ff; 
        10'b0101001110: data <= 10'h000; 
        10'b0101001111: data <= 10'h3ff; 
        10'b0101010000: data <= 10'h000; 
        10'b0101010001: data <= 10'h000; 
        10'b0101010010: data <= 10'h000; 
        10'b0101010011: data <= 10'h000; 
        10'b0101010100: data <= 10'h3ff; 
        10'b0101010101: data <= 10'h000; 
        10'b0101010110: data <= 10'h001; 
        10'b0101010111: data <= 10'h001; 
        10'b0101011000: data <= 10'h001; 
        10'b0101011001: data <= 10'h000; 
        10'b0101011010: data <= 10'h001; 
        10'b0101011011: data <= 10'h001; 
        10'b0101011100: data <= 10'h001; 
        10'b0101011101: data <= 10'h3ff; 
        10'b0101011110: data <= 10'h3f9; 
        10'b0101011111: data <= 10'h3f7; 
        10'b0101100000: data <= 10'h3f7; 
        10'b0101100001: data <= 10'h3fb; 
        10'b0101100010: data <= 10'h3ff; 
        10'b0101100011: data <= 10'h000; 
        10'b0101100100: data <= 10'h000; 
        10'b0101100101: data <= 10'h001; 
        10'b0101100110: data <= 10'h005; 
        10'b0101100111: data <= 10'h004; 
        10'b0101101000: data <= 10'h003; 
        10'b0101101001: data <= 10'h000; 
        10'b0101101010: data <= 10'h000; 
        10'b0101101011: data <= 10'h000; 
        10'b0101101100: data <= 10'h3ff; 
        10'b0101101101: data <= 10'h000; 
        10'b0101101110: data <= 10'h000; 
        10'b0101101111: data <= 10'h3ff; 
        10'b0101110000: data <= 10'h000; 
        10'b0101110001: data <= 10'h001; 
        10'b0101110010: data <= 10'h002; 
        10'b0101110011: data <= 10'h002; 
        10'b0101110100: data <= 10'h002; 
        10'b0101110101: data <= 10'h001; 
        10'b0101110110: data <= 10'h002; 
        10'b0101110111: data <= 10'h001; 
        10'b0101111000: data <= 10'h001; 
        10'b0101111001: data <= 10'h3fc; 
        10'b0101111010: data <= 10'h3f9; 
        10'b0101111011: data <= 10'h3f7; 
        10'b0101111100: data <= 10'h3f8; 
        10'b0101111101: data <= 10'h3fc; 
        10'b0101111110: data <= 10'h3fe; 
        10'b0101111111: data <= 10'h3fe; 
        10'b0110000000: data <= 10'h3fe; 
        10'b0110000001: data <= 10'h001; 
        10'b0110000010: data <= 10'h003; 
        10'b0110000011: data <= 10'h005; 
        10'b0110000100: data <= 10'h003; 
        10'b0110000101: data <= 10'h000; 
        10'b0110000110: data <= 10'h000; 
        10'b0110000111: data <= 10'h000; 
        10'b0110001000: data <= 10'h000; 
        10'b0110001001: data <= 10'h000; 
        10'b0110001010: data <= 10'h3ff; 
        10'b0110001011: data <= 10'h000; 
        10'b0110001100: data <= 10'h3ff; 
        10'b0110001101: data <= 10'h002; 
        10'b0110001110: data <= 10'h003; 
        10'b0110001111: data <= 10'h004; 
        10'b0110010000: data <= 10'h002; 
        10'b0110010001: data <= 10'h002; 
        10'b0110010010: data <= 10'h003; 
        10'b0110010011: data <= 10'h002; 
        10'b0110010100: data <= 10'h000; 
        10'b0110010101: data <= 10'h3fc; 
        10'b0110010110: data <= 10'h3f7; 
        10'b0110010111: data <= 10'h3f7; 
        10'b0110011000: data <= 10'h3f9; 
        10'b0110011001: data <= 10'h3fc; 
        10'b0110011010: data <= 10'h3fe; 
        10'b0110011011: data <= 10'h3fe; 
        10'b0110011100: data <= 10'h000; 
        10'b0110011101: data <= 10'h002; 
        10'b0110011110: data <= 10'h002; 
        10'b0110011111: data <= 10'h005; 
        10'b0110100000: data <= 10'h003; 
        10'b0110100001: data <= 10'h3ff; 
        10'b0110100010: data <= 10'h000; 
        10'b0110100011: data <= 10'h3ff; 
        10'b0110100100: data <= 10'h000; 
        10'b0110100101: data <= 10'h000; 
        10'b0110100110: data <= 10'h000; 
        10'b0110100111: data <= 10'h000; 
        10'b0110101000: data <= 10'h000; 
        10'b0110101001: data <= 10'h003; 
        10'b0110101010: data <= 10'h002; 
        10'b0110101011: data <= 10'h003; 
        10'b0110101100: data <= 10'h002; 
        10'b0110101101: data <= 10'h003; 
        10'b0110101110: data <= 10'h004; 
        10'b0110101111: data <= 10'h001; 
        10'b0110110000: data <= 10'h3fd; 
        10'b0110110001: data <= 10'h3f9; 
        10'b0110110010: data <= 10'h3f6; 
        10'b0110110011: data <= 10'h3f7; 
        10'b0110110100: data <= 10'h3fa; 
        10'b0110110101: data <= 10'h3fd; 
        10'b0110110110: data <= 10'h3ff; 
        10'b0110110111: data <= 10'h3ff; 
        10'b0110111000: data <= 10'h001; 
        10'b0110111001: data <= 10'h001; 
        10'b0110111010: data <= 10'h003; 
        10'b0110111011: data <= 10'h004; 
        10'b0110111100: data <= 10'h002; 
        10'b0110111101: data <= 10'h000; 
        10'b0110111110: data <= 10'h000; 
        10'b0110111111: data <= 10'h3ff; 
        10'b0111000000: data <= 10'h000; 
        10'b0111000001: data <= 10'h000; 
        10'b0111000010: data <= 10'h3ff; 
        10'b0111000011: data <= 10'h000; 
        10'b0111000100: data <= 10'h001; 
        10'b0111000101: data <= 10'h003; 
        10'b0111000110: data <= 10'h004; 
        10'b0111000111: data <= 10'h003; 
        10'b0111001000: data <= 10'h002; 
        10'b0111001001: data <= 10'h002; 
        10'b0111001010: data <= 10'h003; 
        10'b0111001011: data <= 10'h000; 
        10'b0111001100: data <= 10'h3fb; 
        10'b0111001101: data <= 10'h3f6; 
        10'b0111001110: data <= 10'h3f7; 
        10'b0111001111: data <= 10'h3f9; 
        10'b0111010000: data <= 10'h3fc; 
        10'b0111010001: data <= 10'h3fe; 
        10'b0111010010: data <= 10'h000; 
        10'b0111010011: data <= 10'h001; 
        10'b0111010100: data <= 10'h001; 
        10'b0111010101: data <= 10'h002; 
        10'b0111010110: data <= 10'h003; 
        10'b0111010111: data <= 10'h003; 
        10'b0111011000: data <= 10'h001; 
        10'b0111011001: data <= 10'h000; 
        10'b0111011010: data <= 10'h000; 
        10'b0111011011: data <= 10'h000; 
        10'b0111011100: data <= 10'h000; 
        10'b0111011101: data <= 10'h000; 
        10'b0111011110: data <= 10'h3ff; 
        10'b0111011111: data <= 10'h3ff; 
        10'b0111100000: data <= 10'h000; 
        10'b0111100001: data <= 10'h002; 
        10'b0111100010: data <= 10'h003; 
        10'b0111100011: data <= 10'h003; 
        10'b0111100100: data <= 10'h001; 
        10'b0111100101: data <= 10'h002; 
        10'b0111100110: data <= 10'h003; 
        10'b0111100111: data <= 10'h000; 
        10'b0111101000: data <= 10'h3f9; 
        10'b0111101001: data <= 10'h3f7; 
        10'b0111101010: data <= 10'h3f8; 
        10'b0111101011: data <= 10'h3fb; 
        10'b0111101100: data <= 10'h3ff; 
        10'b0111101101: data <= 10'h001; 
        10'b0111101110: data <= 10'h002; 
        10'b0111101111: data <= 10'h002; 
        10'b0111110000: data <= 10'h002; 
        10'b0111110001: data <= 10'h002; 
        10'b0111110010: data <= 10'h001; 
        10'b0111110011: data <= 10'h001; 
        10'b0111110100: data <= 10'h000; 
        10'b0111110101: data <= 10'h000; 
        10'b0111110110: data <= 10'h000; 
        10'b0111110111: data <= 10'h3ff; 
        10'b0111111000: data <= 10'h000; 
        10'b0111111001: data <= 10'h000; 
        10'b0111111010: data <= 10'h000; 
        10'b0111111011: data <= 10'h000; 
        10'b0111111100: data <= 10'h000; 
        10'b0111111101: data <= 10'h001; 
        10'b0111111110: data <= 10'h003; 
        10'b0111111111: data <= 10'h002; 
        10'b1000000000: data <= 10'h001; 
        10'b1000000001: data <= 10'h003; 
        10'b1000000010: data <= 10'h005; 
        10'b1000000011: data <= 10'h000; 
        10'b1000000100: data <= 10'h3fc; 
        10'b1000000101: data <= 10'h3f9; 
        10'b1000000110: data <= 10'h3fb; 
        10'b1000000111: data <= 10'h3ff; 
        10'b1000001000: data <= 10'h002; 
        10'b1000001001: data <= 10'h002; 
        10'b1000001010: data <= 10'h002; 
        10'b1000001011: data <= 10'h001; 
        10'b1000001100: data <= 10'h000; 
        10'b1000001101: data <= 10'h001; 
        10'b1000001110: data <= 10'h001; 
        10'b1000001111: data <= 10'h001; 
        10'b1000010000: data <= 10'h000; 
        10'b1000010001: data <= 10'h000; 
        10'b1000010010: data <= 10'h000; 
        10'b1000010011: data <= 10'h000; 
        10'b1000010100: data <= 10'h000; 
        10'b1000010101: data <= 10'h000; 
        10'b1000010110: data <= 10'h000; 
        10'b1000010111: data <= 10'h3ff; 
        10'b1000011000: data <= 10'h001; 
        10'b1000011001: data <= 10'h001; 
        10'b1000011010: data <= 10'h003; 
        10'b1000011011: data <= 10'h003; 
        10'b1000011100: data <= 10'h002; 
        10'b1000011101: data <= 10'h003; 
        10'b1000011110: data <= 10'h005; 
        10'b1000011111: data <= 10'h004; 
        10'b1000100000: data <= 10'h001; 
        10'b1000100001: data <= 10'h3fe; 
        10'b1000100010: data <= 10'h3ff; 
        10'b1000100011: data <= 10'h000; 
        10'b1000100100: data <= 10'h001; 
        10'b1000100101: data <= 10'h000; 
        10'b1000100110: data <= 10'h3ff; 
        10'b1000100111: data <= 10'h000; 
        10'b1000101000: data <= 10'h001; 
        10'b1000101001: data <= 10'h001; 
        10'b1000101010: data <= 10'h001; 
        10'b1000101011: data <= 10'h000; 
        10'b1000101100: data <= 10'h000; 
        10'b1000101101: data <= 10'h000; 
        10'b1000101110: data <= 10'h3ff; 
        10'b1000101111: data <= 10'h000; 
        10'b1000110000: data <= 10'h000; 
        10'b1000110001: data <= 10'h000; 
        10'b1000110010: data <= 10'h000; 
        10'b1000110011: data <= 10'h3ff; 
        10'b1000110100: data <= 10'h000; 
        10'b1000110101: data <= 10'h001; 
        10'b1000110110: data <= 10'h003; 
        10'b1000110111: data <= 10'h002; 
        10'b1000111000: data <= 10'h003; 
        10'b1000111001: data <= 10'h003; 
        10'b1000111010: data <= 10'h005; 
        10'b1000111011: data <= 10'h005; 
        10'b1000111100: data <= 10'h002; 
        10'b1000111101: data <= 10'h001; 
        10'b1000111110: data <= 10'h3ff; 
        10'b1000111111: data <= 10'h000; 
        10'b1001000000: data <= 10'h000; 
        10'b1001000001: data <= 10'h3ff; 
        10'b1001000010: data <= 10'h3ff; 
        10'b1001000011: data <= 10'h3ff; 
        10'b1001000100: data <= 10'h000; 
        10'b1001000101: data <= 10'h001; 
        10'b1001000110: data <= 10'h001; 
        10'b1001000111: data <= 10'h000; 
        10'b1001001000: data <= 10'h000; 
        10'b1001001001: data <= 10'h000; 
        10'b1001001010: data <= 10'h3ff; 
        10'b1001001011: data <= 10'h000; 
        10'b1001001100: data <= 10'h000; 
        10'b1001001101: data <= 10'h3ff; 
        10'b1001001110: data <= 10'h000; 
        10'b1001001111: data <= 10'h000; 
        10'b1001010000: data <= 10'h000; 
        10'b1001010001: data <= 10'h000; 
        10'b1001010010: data <= 10'h002; 
        10'b1001010011: data <= 10'h003; 
        10'b1001010100: data <= 10'h002; 
        10'b1001010101: data <= 10'h002; 
        10'b1001010110: data <= 10'h004; 
        10'b1001010111: data <= 10'h005; 
        10'b1001011000: data <= 10'h003; 
        10'b1001011001: data <= 10'h001; 
        10'b1001011010: data <= 10'h000; 
        10'b1001011011: data <= 10'h000; 
        10'b1001011100: data <= 10'h000; 
        10'b1001011101: data <= 10'h3ff; 
        10'b1001011110: data <= 10'h3ff; 
        10'b1001011111: data <= 10'h3ff; 
        10'b1001100000: data <= 10'h000; 
        10'b1001100001: data <= 10'h000; 
        10'b1001100010: data <= 10'h3ff; 
        10'b1001100011: data <= 10'h3ff; 
        10'b1001100100: data <= 10'h000; 
        10'b1001100101: data <= 10'h000; 
        10'b1001100110: data <= 10'h000; 
        10'b1001100111: data <= 10'h000; 
        10'b1001101000: data <= 10'h3ff; 
        10'b1001101001: data <= 10'h000; 
        10'b1001101010: data <= 10'h000; 
        10'b1001101011: data <= 10'h000; 
        10'b1001101100: data <= 10'h3ff; 
        10'b1001101101: data <= 10'h000; 
        10'b1001101110: data <= 10'h001; 
        10'b1001101111: data <= 10'h001; 
        10'b1001110000: data <= 10'h003; 
        10'b1001110001: data <= 10'h003; 
        10'b1001110010: data <= 10'h003; 
        10'b1001110011: data <= 10'h003; 
        10'b1001110100: data <= 10'h003; 
        10'b1001110101: data <= 10'h004; 
        10'b1001110110: data <= 10'h002; 
        10'b1001110111: data <= 10'h002; 
        10'b1001111000: data <= 10'h001; 
        10'b1001111001: data <= 10'h3ff; 
        10'b1001111010: data <= 10'h3ff; 
        10'b1001111011: data <= 10'h000; 
        10'b1001111100: data <= 10'h3ff; 
        10'b1001111101: data <= 10'h3ff; 
        10'b1001111110: data <= 10'h000; 
        10'b1001111111: data <= 10'h000; 
        10'b1010000000: data <= 10'h000; 
        10'b1010000001: data <= 10'h000; 
        10'b1010000010: data <= 10'h000; 
        10'b1010000011: data <= 10'h000; 
        10'b1010000100: data <= 10'h3ff; 
        10'b1010000101: data <= 10'h000; 
        10'b1010000110: data <= 10'h000; 
        10'b1010000111: data <= 10'h3ff; 
        10'b1010001000: data <= 10'h3ff; 
        10'b1010001001: data <= 10'h000; 
        10'b1010001010: data <= 10'h000; 
        10'b1010001011: data <= 10'h001; 
        10'b1010001100: data <= 10'h001; 
        10'b1010001101: data <= 10'h003; 
        10'b1010001110: data <= 10'h004; 
        10'b1010001111: data <= 10'h004; 
        10'b1010010000: data <= 10'h004; 
        10'b1010010001: data <= 10'h003; 
        10'b1010010010: data <= 10'h002; 
        10'b1010010011: data <= 10'h001; 
        10'b1010010100: data <= 10'h000; 
        10'b1010010101: data <= 10'h000; 
        10'b1010010110: data <= 10'h3fe; 
        10'b1010010111: data <= 10'h3fe; 
        10'b1010011000: data <= 10'h3fe; 
        10'b1010011001: data <= 10'h3ff; 
        10'b1010011010: data <= 10'h3ff; 
        10'b1010011011: data <= 10'h000; 
        10'b1010011100: data <= 10'h000; 
        10'b1010011101: data <= 10'h000; 
        10'b1010011110: data <= 10'h000; 
        10'b1010011111: data <= 10'h3ff; 
        10'b1010100000: data <= 10'h000; 
        10'b1010100001: data <= 10'h000; 
        10'b1010100010: data <= 10'h3ff; 
        10'b1010100011: data <= 10'h000; 
        10'b1010100100: data <= 10'h000; 
        10'b1010100101: data <= 10'h000; 
        10'b1010100110: data <= 10'h3ff; 
        10'b1010100111: data <= 10'h3ff; 
        10'b1010101000: data <= 10'h3ff; 
        10'b1010101001: data <= 10'h3ff; 
        10'b1010101010: data <= 10'h001; 
        10'b1010101011: data <= 10'h000; 
        10'b1010101100: data <= 10'h001; 
        10'b1010101101: data <= 10'h002; 
        10'b1010101110: data <= 10'h001; 
        10'b1010101111: data <= 10'h3ff; 
        10'b1010110000: data <= 10'h3ff; 
        10'b1010110001: data <= 10'h3ff; 
        10'b1010110010: data <= 10'h3ff; 
        10'b1010110011: data <= 10'h3fe; 
        10'b1010110100: data <= 10'h3ff; 
        10'b1010110101: data <= 10'h3ff; 
        10'b1010110110: data <= 10'h000; 
        10'b1010110111: data <= 10'h000; 
        10'b1010111000: data <= 10'h3ff; 
        10'b1010111001: data <= 10'h000; 
        10'b1010111010: data <= 10'h000; 
        10'b1010111011: data <= 10'h3ff; 
        10'b1010111100: data <= 10'h000; 
        10'b1010111101: data <= 10'h000; 
        10'b1010111110: data <= 10'h000; 
        10'b1010111111: data <= 10'h000; 
        10'b1011000000: data <= 10'h000; 
        10'b1011000001: data <= 10'h000; 
        10'b1011000010: data <= 10'h3ff; 
        10'b1011000011: data <= 10'h000; 
        10'b1011000100: data <= 10'h3ff; 
        10'b1011000101: data <= 10'h3ff; 
        10'b1011000110: data <= 10'h3fe; 
        10'b1011000111: data <= 10'h3fe; 
        10'b1011001000: data <= 10'h3fd; 
        10'b1011001001: data <= 10'h3fe; 
        10'b1011001010: data <= 10'h3fd; 
        10'b1011001011: data <= 10'h3fe; 
        10'b1011001100: data <= 10'h3fe; 
        10'b1011001101: data <= 10'h3ff; 
        10'b1011001110: data <= 10'h3ff; 
        10'b1011001111: data <= 10'h3ff; 
        10'b1011010000: data <= 10'h3ff; 
        10'b1011010001: data <= 10'h3ff; 
        10'b1011010010: data <= 10'h000; 
        10'b1011010011: data <= 10'h000; 
        10'b1011010100: data <= 10'h000; 
        10'b1011010101: data <= 10'h000; 
        10'b1011010110: data <= 10'h000; 
        10'b1011010111: data <= 10'h000; 
        10'b1011011000: data <= 10'h000; 
        10'b1011011001: data <= 10'h000; 
        10'b1011011010: data <= 10'h000; 
        10'b1011011011: data <= 10'h000; 
        10'b1011011100: data <= 10'h000; 
        10'b1011011101: data <= 10'h000; 
        10'b1011011110: data <= 10'h3ff; 
        10'b1011011111: data <= 10'h000; 
        10'b1011100000: data <= 10'h000; 
        10'b1011100001: data <= 10'h3ff; 
        10'b1011100010: data <= 10'h3ff; 
        10'b1011100011: data <= 10'h3ff; 
        10'b1011100100: data <= 10'h000; 
        10'b1011100101: data <= 10'h3ff; 
        10'b1011100110: data <= 10'h3ff; 
        10'b1011100111: data <= 10'h000; 
        10'b1011101000: data <= 10'h3ff; 
        10'b1011101001: data <= 10'h3ff; 
        10'b1011101010: data <= 10'h3ff; 
        10'b1011101011: data <= 10'h3ff; 
        10'b1011101100: data <= 10'h000; 
        10'b1011101101: data <= 10'h3ff; 
        10'b1011101110: data <= 10'h3ff; 
        10'b1011101111: data <= 10'h000; 
        10'b1011110000: data <= 10'h3ff; 
        10'b1011110001: data <= 10'h000; 
        10'b1011110010: data <= 10'h000; 
        10'b1011110011: data <= 10'h000; 
        10'b1011110100: data <= 10'h3ff; 
        10'b1011110101: data <= 10'h000; 
        10'b1011110110: data <= 10'h000; 
        10'b1011110111: data <= 10'h000; 
        10'b1011111000: data <= 10'h000; 
        10'b1011111001: data <= 10'h000; 
        10'b1011111010: data <= 10'h000; 
        10'b1011111011: data <= 10'h3ff; 
        10'b1011111100: data <= 10'h000; 
        10'b1011111101: data <= 10'h000; 
        10'b1011111110: data <= 10'h000; 
        10'b1011111111: data <= 10'h000; 
        10'b1100000000: data <= 10'h000; 
        10'b1100000001: data <= 10'h000; 
        10'b1100000010: data <= 10'h000; 
        10'b1100000011: data <= 10'h3ff; 
        10'b1100000100: data <= 10'h000; 
        10'b1100000101: data <= 10'h000; 
        10'b1100000110: data <= 10'h000; 
        10'b1100000111: data <= 10'h000; 
        10'b1100001000: data <= 10'h3ff; 
        10'b1100001001: data <= 10'h3ff; 
        10'b1100001010: data <= 10'h3ff; 
        10'b1100001011: data <= 10'h000; 
        10'b1100001100: data <= 10'h000; 
        10'b1100001101: data <= 10'h3ff; 
        10'b1100001110: data <= 10'h3ff; 
        10'b1100001111: data <= 10'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 5) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 11'h7ff; 
        10'b0000000001: data <= 11'h001; 
        10'b0000000010: data <= 11'h000; 
        10'b0000000011: data <= 11'h000; 
        10'b0000000100: data <= 11'h001; 
        10'b0000000101: data <= 11'h000; 
        10'b0000000110: data <= 11'h7ff; 
        10'b0000000111: data <= 11'h7ff; 
        10'b0000001000: data <= 11'h000; 
        10'b0000001001: data <= 11'h000; 
        10'b0000001010: data <= 11'h001; 
        10'b0000001011: data <= 11'h000; 
        10'b0000001100: data <= 11'h000; 
        10'b0000001101: data <= 11'h7ff; 
        10'b0000001110: data <= 11'h000; 
        10'b0000001111: data <= 11'h7ff; 
        10'b0000010000: data <= 11'h7ff; 
        10'b0000010001: data <= 11'h000; 
        10'b0000010010: data <= 11'h7ff; 
        10'b0000010011: data <= 11'h001; 
        10'b0000010100: data <= 11'h7ff; 
        10'b0000010101: data <= 11'h000; 
        10'b0000010110: data <= 11'h7ff; 
        10'b0000010111: data <= 11'h000; 
        10'b0000011000: data <= 11'h000; 
        10'b0000011001: data <= 11'h000; 
        10'b0000011010: data <= 11'h000; 
        10'b0000011011: data <= 11'h000; 
        10'b0000011100: data <= 11'h000; 
        10'b0000011101: data <= 11'h001; 
        10'b0000011110: data <= 11'h000; 
        10'b0000011111: data <= 11'h7ff; 
        10'b0000100000: data <= 11'h7ff; 
        10'b0000100001: data <= 11'h000; 
        10'b0000100010: data <= 11'h7ff; 
        10'b0000100011: data <= 11'h000; 
        10'b0000100100: data <= 11'h7ff; 
        10'b0000100101: data <= 11'h7ff; 
        10'b0000100110: data <= 11'h7ff; 
        10'b0000100111: data <= 11'h000; 
        10'b0000101000: data <= 11'h001; 
        10'b0000101001: data <= 11'h7ff; 
        10'b0000101010: data <= 11'h7ff; 
        10'b0000101011: data <= 11'h000; 
        10'b0000101100: data <= 11'h7ff; 
        10'b0000101101: data <= 11'h7ff; 
        10'b0000101110: data <= 11'h000; 
        10'b0000101111: data <= 11'h001; 
        10'b0000110000: data <= 11'h7ff; 
        10'b0000110001: data <= 11'h000; 
        10'b0000110010: data <= 11'h7ff; 
        10'b0000110011: data <= 11'h7ff; 
        10'b0000110100: data <= 11'h000; 
        10'b0000110101: data <= 11'h000; 
        10'b0000110110: data <= 11'h000; 
        10'b0000110111: data <= 11'h001; 
        10'b0000111000: data <= 11'h7ff; 
        10'b0000111001: data <= 11'h7ff; 
        10'b0000111010: data <= 11'h7ff; 
        10'b0000111011: data <= 11'h000; 
        10'b0000111100: data <= 11'h000; 
        10'b0000111101: data <= 11'h7ff; 
        10'b0000111110: data <= 11'h000; 
        10'b0000111111: data <= 11'h001; 
        10'b0001000000: data <= 11'h000; 
        10'b0001000001: data <= 11'h7ff; 
        10'b0001000010: data <= 11'h7ff; 
        10'b0001000011: data <= 11'h7fe; 
        10'b0001000100: data <= 11'h7fe; 
        10'b0001000101: data <= 11'h7ff; 
        10'b0001000110: data <= 11'h7fe; 
        10'b0001000111: data <= 11'h7fe; 
        10'b0001001000: data <= 11'h7fe; 
        10'b0001001001: data <= 11'h000; 
        10'b0001001010: data <= 11'h7ff; 
        10'b0001001011: data <= 11'h7fe; 
        10'b0001001100: data <= 11'h000; 
        10'b0001001101: data <= 11'h001; 
        10'b0001001110: data <= 11'h000; 
        10'b0001001111: data <= 11'h7ff; 
        10'b0001010000: data <= 11'h001; 
        10'b0001010001: data <= 11'h7ff; 
        10'b0001010010: data <= 11'h000; 
        10'b0001010011: data <= 11'h000; 
        10'b0001010100: data <= 11'h7ff; 
        10'b0001010101: data <= 11'h000; 
        10'b0001010110: data <= 11'h001; 
        10'b0001010111: data <= 11'h7ff; 
        10'b0001011000: data <= 11'h7ff; 
        10'b0001011001: data <= 11'h001; 
        10'b0001011010: data <= 11'h000; 
        10'b0001011011: data <= 11'h000; 
        10'b0001011100: data <= 11'h000; 
        10'b0001011101: data <= 11'h000; 
        10'b0001011110: data <= 11'h000; 
        10'b0001011111: data <= 11'h7fe; 
        10'b0001100000: data <= 11'h7fe; 
        10'b0001100001: data <= 11'h7ff; 
        10'b0001100010: data <= 11'h7fe; 
        10'b0001100011: data <= 11'h7fe; 
        10'b0001100100: data <= 11'h000; 
        10'b0001100101: data <= 11'h000; 
        10'b0001100110: data <= 11'h7fe; 
        10'b0001100111: data <= 11'h7fe; 
        10'b0001101000: data <= 11'h7fd; 
        10'b0001101001: data <= 11'h7fe; 
        10'b0001101010: data <= 11'h7fd; 
        10'b0001101011: data <= 11'h7fe; 
        10'b0001101100: data <= 11'h7ff; 
        10'b0001101101: data <= 11'h000; 
        10'b0001101110: data <= 11'h000; 
        10'b0001101111: data <= 11'h7ff; 
        10'b0001110000: data <= 11'h000; 
        10'b0001110001: data <= 11'h7ff; 
        10'b0001110010: data <= 11'h7ff; 
        10'b0001110011: data <= 11'h7ff; 
        10'b0001110100: data <= 11'h7ff; 
        10'b0001110101: data <= 11'h000; 
        10'b0001110110: data <= 11'h000; 
        10'b0001110111: data <= 11'h7ff; 
        10'b0001111000: data <= 11'h000; 
        10'b0001111001: data <= 11'h000; 
        10'b0001111010: data <= 11'h7fe; 
        10'b0001111011: data <= 11'h7fe; 
        10'b0001111100: data <= 11'h7fe; 
        10'b0001111101: data <= 11'h7fe; 
        10'b0001111110: data <= 11'h7ff; 
        10'b0001111111: data <= 11'h000; 
        10'b0010000000: data <= 11'h7fe; 
        10'b0010000001: data <= 11'h7fe; 
        10'b0010000010: data <= 11'h7fe; 
        10'b0010000011: data <= 11'h7fe; 
        10'b0010000100: data <= 11'h7ff; 
        10'b0010000101: data <= 11'h7fd; 
        10'b0010000110: data <= 11'h7ff; 
        10'b0010000111: data <= 11'h000; 
        10'b0010001000: data <= 11'h7ff; 
        10'b0010001001: data <= 11'h7ff; 
        10'b0010001010: data <= 11'h7ff; 
        10'b0010001011: data <= 11'h000; 
        10'b0010001100: data <= 11'h000; 
        10'b0010001101: data <= 11'h7ff; 
        10'b0010001110: data <= 11'h000; 
        10'b0010001111: data <= 11'h7ff; 
        10'b0010010000: data <= 11'h000; 
        10'b0010010001: data <= 11'h7ff; 
        10'b0010010010: data <= 11'h000; 
        10'b0010010011: data <= 11'h7ff; 
        10'b0010010100: data <= 11'h000; 
        10'b0010010101: data <= 11'h7fe; 
        10'b0010010110: data <= 11'h7ff; 
        10'b0010010111: data <= 11'h000; 
        10'b0010011000: data <= 11'h002; 
        10'b0010011001: data <= 11'h004; 
        10'b0010011010: data <= 11'h005; 
        10'b0010011011: data <= 11'h005; 
        10'b0010011100: data <= 11'h005; 
        10'b0010011101: data <= 11'h006; 
        10'b0010011110: data <= 11'h006; 
        10'b0010011111: data <= 11'h002; 
        10'b0010100000: data <= 11'h000; 
        10'b0010100001: data <= 11'h001; 
        10'b0010100010: data <= 11'h7ff; 
        10'b0010100011: data <= 11'h000; 
        10'b0010100100: data <= 11'h7fd; 
        10'b0010100101: data <= 11'h7fe; 
        10'b0010100110: data <= 11'h000; 
        10'b0010100111: data <= 11'h7ff; 
        10'b0010101000: data <= 11'h7ff; 
        10'b0010101001: data <= 11'h000; 
        10'b0010101010: data <= 11'h000; 
        10'b0010101011: data <= 11'h000; 
        10'b0010101100: data <= 11'h000; 
        10'b0010101101: data <= 11'h000; 
        10'b0010101110: data <= 11'h000; 
        10'b0010101111: data <= 11'h000; 
        10'b0010110000: data <= 11'h7ff; 
        10'b0010110001: data <= 11'h7fe; 
        10'b0010110010: data <= 11'h001; 
        10'b0010110011: data <= 11'h000; 
        10'b0010110100: data <= 11'h003; 
        10'b0010110101: data <= 11'h003; 
        10'b0010110110: data <= 11'h003; 
        10'b0010110111: data <= 11'h004; 
        10'b0010111000: data <= 11'h005; 
        10'b0010111001: data <= 11'h007; 
        10'b0010111010: data <= 11'h007; 
        10'b0010111011: data <= 11'h006; 
        10'b0010111100: data <= 11'h006; 
        10'b0010111101: data <= 11'h006; 
        10'b0010111110: data <= 11'h004; 
        10'b0010111111: data <= 11'h001; 
        10'b0011000000: data <= 11'h7fd; 
        10'b0011000001: data <= 11'h7fd; 
        10'b0011000010: data <= 11'h7fe; 
        10'b0011000011: data <= 11'h000; 
        10'b0011000100: data <= 11'h001; 
        10'b0011000101: data <= 11'h000; 
        10'b0011000110: data <= 11'h000; 
        10'b0011000111: data <= 11'h7fe; 
        10'b0011001000: data <= 11'h7fd; 
        10'b0011001001: data <= 11'h000; 
        10'b0011001010: data <= 11'h7ff; 
        10'b0011001011: data <= 11'h000; 
        10'b0011001100: data <= 11'h7ff; 
        10'b0011001101: data <= 11'h000; 
        10'b0011001110: data <= 11'h000; 
        10'b0011001111: data <= 11'h002; 
        10'b0011010000: data <= 11'h005; 
        10'b0011010001: data <= 11'h005; 
        10'b0011010010: data <= 11'h002; 
        10'b0011010011: data <= 11'h003; 
        10'b0011010100: data <= 11'h004; 
        10'b0011010101: data <= 11'h008; 
        10'b0011010110: data <= 11'h006; 
        10'b0011010111: data <= 11'h005; 
        10'b0011011000: data <= 11'h002; 
        10'b0011011001: data <= 11'h004; 
        10'b0011011010: data <= 11'h004; 
        10'b0011011011: data <= 11'h002; 
        10'b0011011100: data <= 11'h7fe; 
        10'b0011011101: data <= 11'h7fd; 
        10'b0011011110: data <= 11'h7fe; 
        10'b0011011111: data <= 11'h000; 
        10'b0011100000: data <= 11'h001; 
        10'b0011100001: data <= 11'h000; 
        10'b0011100010: data <= 11'h000; 
        10'b0011100011: data <= 11'h000; 
        10'b0011100100: data <= 11'h7fe; 
        10'b0011100101: data <= 11'h7fe; 
        10'b0011100110: data <= 11'h7ff; 
        10'b0011100111: data <= 11'h7fe; 
        10'b0011101000: data <= 11'h7ff; 
        10'b0011101001: data <= 11'h7ff; 
        10'b0011101010: data <= 11'h002; 
        10'b0011101011: data <= 11'h003; 
        10'b0011101100: data <= 11'h001; 
        10'b0011101101: data <= 11'h001; 
        10'b0011101110: data <= 11'h001; 
        10'b0011101111: data <= 11'h004; 
        10'b0011110000: data <= 11'h00a; 
        10'b0011110001: data <= 11'h008; 
        10'b0011110010: data <= 11'h008; 
        10'b0011110011: data <= 11'h002; 
        10'b0011110100: data <= 11'h002; 
        10'b0011110101: data <= 11'h002; 
        10'b0011110110: data <= 11'h005; 
        10'b0011110111: data <= 11'h008; 
        10'b0011111000: data <= 11'h7ff; 
        10'b0011111001: data <= 11'h7fd; 
        10'b0011111010: data <= 11'h000; 
        10'b0011111011: data <= 11'h7ff; 
        10'b0011111100: data <= 11'h000; 
        10'b0011111101: data <= 11'h000; 
        10'b0011111110: data <= 11'h000; 
        10'b0011111111: data <= 11'h000; 
        10'b0100000000: data <= 11'h7fe; 
        10'b0100000001: data <= 11'h7fe; 
        10'b0100000010: data <= 11'h7fe; 
        10'b0100000011: data <= 11'h7ff; 
        10'b0100000100: data <= 11'h7ff; 
        10'b0100000101: data <= 11'h7ff; 
        10'b0100000110: data <= 11'h002; 
        10'b0100000111: data <= 11'h7ff; 
        10'b0100001000: data <= 11'h001; 
        10'b0100001001: data <= 11'h003; 
        10'b0100001010: data <= 11'h002; 
        10'b0100001011: data <= 11'h002; 
        10'b0100001100: data <= 11'h006; 
        10'b0100001101: data <= 11'h008; 
        10'b0100001110: data <= 11'h009; 
        10'b0100001111: data <= 11'h005; 
        10'b0100010000: data <= 11'h002; 
        10'b0100010001: data <= 11'h000; 
        10'b0100010010: data <= 11'h004; 
        10'b0100010011: data <= 11'h008; 
        10'b0100010100: data <= 11'h002; 
        10'b0100010101: data <= 11'h7fe; 
        10'b0100010110: data <= 11'h000; 
        10'b0100010111: data <= 11'h000; 
        10'b0100011000: data <= 11'h7ff; 
        10'b0100011001: data <= 11'h001; 
        10'b0100011010: data <= 11'h7ff; 
        10'b0100011011: data <= 11'h7fe; 
        10'b0100011100: data <= 11'h7fe; 
        10'b0100011101: data <= 11'h7ff; 
        10'b0100011110: data <= 11'h7ff; 
        10'b0100011111: data <= 11'h000; 
        10'b0100100000: data <= 11'h001; 
        10'b0100100001: data <= 11'h000; 
        10'b0100100010: data <= 11'h7ff; 
        10'b0100100011: data <= 11'h000; 
        10'b0100100100: data <= 11'h001; 
        10'b0100100101: data <= 11'h000; 
        10'b0100100110: data <= 11'h7fd; 
        10'b0100100111: data <= 11'h7fb; 
        10'b0100101000: data <= 11'h7fd; 
        10'b0100101001: data <= 11'h003; 
        10'b0100101010: data <= 11'h007; 
        10'b0100101011: data <= 11'h007; 
        10'b0100101100: data <= 11'h006; 
        10'b0100101101: data <= 11'h005; 
        10'b0100101110: data <= 11'h007; 
        10'b0100101111: data <= 11'h009; 
        10'b0100110000: data <= 11'h004; 
        10'b0100110001: data <= 11'h7fe; 
        10'b0100110010: data <= 11'h7fe; 
        10'b0100110011: data <= 11'h7ff; 
        10'b0100110100: data <= 11'h7ff; 
        10'b0100110101: data <= 11'h7ff; 
        10'b0100110110: data <= 11'h001; 
        10'b0100110111: data <= 11'h000; 
        10'b0100111000: data <= 11'h7fd; 
        10'b0100111001: data <= 11'h7ff; 
        10'b0100111010: data <= 11'h001; 
        10'b0100111011: data <= 11'h003; 
        10'b0100111100: data <= 11'h002; 
        10'b0100111101: data <= 11'h7ff; 
        10'b0100111110: data <= 11'h001; 
        10'b0100111111: data <= 11'h000; 
        10'b0101000000: data <= 11'h001; 
        10'b0101000001: data <= 11'h7ff; 
        10'b0101000010: data <= 11'h7f9; 
        10'b0101000011: data <= 11'h7f2; 
        10'b0101000100: data <= 11'h7f3; 
        10'b0101000101: data <= 11'h7fb; 
        10'b0101000110: data <= 11'h7ff; 
        10'b0101000111: data <= 11'h004; 
        10'b0101001000: data <= 11'h006; 
        10'b0101001001: data <= 11'h005; 
        10'b0101001010: data <= 11'h007; 
        10'b0101001011: data <= 11'h008; 
        10'b0101001100: data <= 11'h006; 
        10'b0101001101: data <= 11'h7ff; 
        10'b0101001110: data <= 11'h000; 
        10'b0101001111: data <= 11'h7ff; 
        10'b0101010000: data <= 11'h7ff; 
        10'b0101010001: data <= 11'h000; 
        10'b0101010010: data <= 11'h000; 
        10'b0101010011: data <= 11'h000; 
        10'b0101010100: data <= 11'h7fe; 
        10'b0101010101: data <= 11'h000; 
        10'b0101010110: data <= 11'h003; 
        10'b0101010111: data <= 11'h003; 
        10'b0101011000: data <= 11'h001; 
        10'b0101011001: data <= 11'h000; 
        10'b0101011010: data <= 11'h002; 
        10'b0101011011: data <= 11'h001; 
        10'b0101011100: data <= 11'h003; 
        10'b0101011101: data <= 11'h7fe; 
        10'b0101011110: data <= 11'h7f2; 
        10'b0101011111: data <= 11'h7ee; 
        10'b0101100000: data <= 11'h7ee; 
        10'b0101100001: data <= 11'h7f6; 
        10'b0101100010: data <= 11'h7fe; 
        10'b0101100011: data <= 11'h7ff; 
        10'b0101100100: data <= 11'h001; 
        10'b0101100101: data <= 11'h003; 
        10'b0101100110: data <= 11'h00a; 
        10'b0101100111: data <= 11'h009; 
        10'b0101101000: data <= 11'h006; 
        10'b0101101001: data <= 11'h000; 
        10'b0101101010: data <= 11'h7ff; 
        10'b0101101011: data <= 11'h7ff; 
        10'b0101101100: data <= 11'h7ff; 
        10'b0101101101: data <= 11'h000; 
        10'b0101101110: data <= 11'h000; 
        10'b0101101111: data <= 11'h7ff; 
        10'b0101110000: data <= 11'h7ff; 
        10'b0101110001: data <= 11'h002; 
        10'b0101110010: data <= 11'h003; 
        10'b0101110011: data <= 11'h004; 
        10'b0101110100: data <= 11'h003; 
        10'b0101110101: data <= 11'h002; 
        10'b0101110110: data <= 11'h003; 
        10'b0101110111: data <= 11'h003; 
        10'b0101111000: data <= 11'h002; 
        10'b0101111001: data <= 11'h7f7; 
        10'b0101111010: data <= 11'h7f1; 
        10'b0101111011: data <= 11'h7ee; 
        10'b0101111100: data <= 11'h7f1; 
        10'b0101111101: data <= 11'h7f8; 
        10'b0101111110: data <= 11'h7fc; 
        10'b0101111111: data <= 11'h7fb; 
        10'b0110000000: data <= 11'h7fc; 
        10'b0110000001: data <= 11'h002; 
        10'b0110000010: data <= 11'h006; 
        10'b0110000011: data <= 11'h00a; 
        10'b0110000100: data <= 11'h006; 
        10'b0110000101: data <= 11'h001; 
        10'b0110000110: data <= 11'h000; 
        10'b0110000111: data <= 11'h001; 
        10'b0110001000: data <= 11'h000; 
        10'b0110001001: data <= 11'h000; 
        10'b0110001010: data <= 11'h7ff; 
        10'b0110001011: data <= 11'h7ff; 
        10'b0110001100: data <= 11'h7fe; 
        10'b0110001101: data <= 11'h005; 
        10'b0110001110: data <= 11'h006; 
        10'b0110001111: data <= 11'h007; 
        10'b0110010000: data <= 11'h003; 
        10'b0110010001: data <= 11'h004; 
        10'b0110010010: data <= 11'h006; 
        10'b0110010011: data <= 11'h004; 
        10'b0110010100: data <= 11'h001; 
        10'b0110010101: data <= 11'h7f8; 
        10'b0110010110: data <= 11'h7ef; 
        10'b0110010111: data <= 11'h7ee; 
        10'b0110011000: data <= 11'h7f1; 
        10'b0110011001: data <= 11'h7f8; 
        10'b0110011010: data <= 11'h7fc; 
        10'b0110011011: data <= 11'h7fc; 
        10'b0110011100: data <= 11'h000; 
        10'b0110011101: data <= 11'h003; 
        10'b0110011110: data <= 11'h004; 
        10'b0110011111: data <= 11'h00a; 
        10'b0110100000: data <= 11'h005; 
        10'b0110100001: data <= 11'h7ff; 
        10'b0110100010: data <= 11'h7ff; 
        10'b0110100011: data <= 11'h7ff; 
        10'b0110100100: data <= 11'h001; 
        10'b0110100101: data <= 11'h000; 
        10'b0110100110: data <= 11'h7ff; 
        10'b0110100111: data <= 11'h000; 
        10'b0110101000: data <= 11'h000; 
        10'b0110101001: data <= 11'h006; 
        10'b0110101010: data <= 11'h005; 
        10'b0110101011: data <= 11'h006; 
        10'b0110101100: data <= 11'h004; 
        10'b0110101101: data <= 11'h006; 
        10'b0110101110: data <= 11'h007; 
        10'b0110101111: data <= 11'h002; 
        10'b0110110000: data <= 11'h7fa; 
        10'b0110110001: data <= 11'h7f2; 
        10'b0110110010: data <= 11'h7ed; 
        10'b0110110011: data <= 11'h7ee; 
        10'b0110110100: data <= 11'h7f4; 
        10'b0110110101: data <= 11'h7fa; 
        10'b0110110110: data <= 11'h7fe; 
        10'b0110110111: data <= 11'h7fe; 
        10'b0110111000: data <= 11'h002; 
        10'b0110111001: data <= 11'h002; 
        10'b0110111010: data <= 11'h006; 
        10'b0110111011: data <= 11'h007; 
        10'b0110111100: data <= 11'h004; 
        10'b0110111101: data <= 11'h000; 
        10'b0110111110: data <= 11'h000; 
        10'b0110111111: data <= 11'h7ff; 
        10'b0111000000: data <= 11'h000; 
        10'b0111000001: data <= 11'h001; 
        10'b0111000010: data <= 11'h7ff; 
        10'b0111000011: data <= 11'h7ff; 
        10'b0111000100: data <= 11'h001; 
        10'b0111000101: data <= 11'h006; 
        10'b0111000110: data <= 11'h007; 
        10'b0111000111: data <= 11'h006; 
        10'b0111001000: data <= 11'h004; 
        10'b0111001001: data <= 11'h004; 
        10'b0111001010: data <= 11'h007; 
        10'b0111001011: data <= 11'h7ff; 
        10'b0111001100: data <= 11'h7f5; 
        10'b0111001101: data <= 11'h7ed; 
        10'b0111001110: data <= 11'h7ed; 
        10'b0111001111: data <= 11'h7f1; 
        10'b0111010000: data <= 11'h7f8; 
        10'b0111010001: data <= 11'h7fc; 
        10'b0111010010: data <= 11'h000; 
        10'b0111010011: data <= 11'h001; 
        10'b0111010100: data <= 11'h003; 
        10'b0111010101: data <= 11'h004; 
        10'b0111010110: data <= 11'h006; 
        10'b0111010111: data <= 11'h005; 
        10'b0111011000: data <= 11'h002; 
        10'b0111011001: data <= 11'h000; 
        10'b0111011010: data <= 11'h7ff; 
        10'b0111011011: data <= 11'h7ff; 
        10'b0111011100: data <= 11'h7ff; 
        10'b0111011101: data <= 11'h000; 
        10'b0111011110: data <= 11'h7ff; 
        10'b0111011111: data <= 11'h7fe; 
        10'b0111100000: data <= 11'h000; 
        10'b0111100001: data <= 11'h004; 
        10'b0111100010: data <= 11'h005; 
        10'b0111100011: data <= 11'h005; 
        10'b0111100100: data <= 11'h002; 
        10'b0111100101: data <= 11'h004; 
        10'b0111100110: data <= 11'h006; 
        10'b0111100111: data <= 11'h7ff; 
        10'b0111101000: data <= 11'h7f3; 
        10'b0111101001: data <= 11'h7ed; 
        10'b0111101010: data <= 11'h7ef; 
        10'b0111101011: data <= 11'h7f6; 
        10'b0111101100: data <= 11'h7ff; 
        10'b0111101101: data <= 11'h003; 
        10'b0111101110: data <= 11'h004; 
        10'b0111101111: data <= 11'h003; 
        10'b0111110000: data <= 11'h004; 
        10'b0111110001: data <= 11'h003; 
        10'b0111110010: data <= 11'h003; 
        10'b0111110011: data <= 11'h003; 
        10'b0111110100: data <= 11'h000; 
        10'b0111110101: data <= 11'h000; 
        10'b0111110110: data <= 11'h000; 
        10'b0111110111: data <= 11'h7ff; 
        10'b0111111000: data <= 11'h7ff; 
        10'b0111111001: data <= 11'h000; 
        10'b0111111010: data <= 11'h000; 
        10'b0111111011: data <= 11'h7ff; 
        10'b0111111100: data <= 11'h7ff; 
        10'b0111111101: data <= 11'h003; 
        10'b0111111110: data <= 11'h005; 
        10'b0111111111: data <= 11'h003; 
        10'b1000000000: data <= 11'h002; 
        10'b1000000001: data <= 11'h005; 
        10'b1000000010: data <= 11'h00a; 
        10'b1000000011: data <= 11'h000; 
        10'b1000000100: data <= 11'h7f8; 
        10'b1000000101: data <= 11'h7f3; 
        10'b1000000110: data <= 11'h7f7; 
        10'b1000000111: data <= 11'h7fd; 
        10'b1000001000: data <= 11'h003; 
        10'b1000001001: data <= 11'h003; 
        10'b1000001010: data <= 11'h003; 
        10'b1000001011: data <= 11'h002; 
        10'b1000001100: data <= 11'h001; 
        10'b1000001101: data <= 11'h001; 
        10'b1000001110: data <= 11'h003; 
        10'b1000001111: data <= 11'h002; 
        10'b1000010000: data <= 11'h000; 
        10'b1000010001: data <= 11'h7ff; 
        10'b1000010010: data <= 11'h000; 
        10'b1000010011: data <= 11'h000; 
        10'b1000010100: data <= 11'h000; 
        10'b1000010101: data <= 11'h7ff; 
        10'b1000010110: data <= 11'h7ff; 
        10'b1000010111: data <= 11'h7fe; 
        10'b1000011000: data <= 11'h001; 
        10'b1000011001: data <= 11'h003; 
        10'b1000011010: data <= 11'h007; 
        10'b1000011011: data <= 11'h006; 
        10'b1000011100: data <= 11'h005; 
        10'b1000011101: data <= 11'h007; 
        10'b1000011110: data <= 11'h00a; 
        10'b1000011111: data <= 11'h007; 
        10'b1000100000: data <= 11'h002; 
        10'b1000100001: data <= 11'h7fd; 
        10'b1000100010: data <= 11'h7ff; 
        10'b1000100011: data <= 11'h7ff; 
        10'b1000100100: data <= 11'h002; 
        10'b1000100101: data <= 11'h7ff; 
        10'b1000100110: data <= 11'h7ff; 
        10'b1000100111: data <= 11'h7ff; 
        10'b1000101000: data <= 11'h002; 
        10'b1000101001: data <= 11'h001; 
        10'b1000101010: data <= 11'h003; 
        10'b1000101011: data <= 11'h000; 
        10'b1000101100: data <= 11'h000; 
        10'b1000101101: data <= 11'h7ff; 
        10'b1000101110: data <= 11'h7fe; 
        10'b1000101111: data <= 11'h001; 
        10'b1000110000: data <= 11'h001; 
        10'b1000110001: data <= 11'h001; 
        10'b1000110010: data <= 11'h000; 
        10'b1000110011: data <= 11'h7ff; 
        10'b1000110100: data <= 11'h7ff; 
        10'b1000110101: data <= 11'h003; 
        10'b1000110110: data <= 11'h006; 
        10'b1000110111: data <= 11'h004; 
        10'b1000111000: data <= 11'h005; 
        10'b1000111001: data <= 11'h006; 
        10'b1000111010: data <= 11'h00a; 
        10'b1000111011: data <= 11'h00a; 
        10'b1000111100: data <= 11'h005; 
        10'b1000111101: data <= 11'h001; 
        10'b1000111110: data <= 11'h7ff; 
        10'b1000111111: data <= 11'h001; 
        10'b1001000000: data <= 11'h001; 
        10'b1001000001: data <= 11'h7ff; 
        10'b1001000010: data <= 11'h7ff; 
        10'b1001000011: data <= 11'h7fe; 
        10'b1001000100: data <= 11'h001; 
        10'b1001000101: data <= 11'h001; 
        10'b1001000110: data <= 11'h002; 
        10'b1001000111: data <= 11'h001; 
        10'b1001001000: data <= 11'h7ff; 
        10'b1001001001: data <= 11'h000; 
        10'b1001001010: data <= 11'h7ff; 
        10'b1001001011: data <= 11'h7ff; 
        10'b1001001100: data <= 11'h7ff; 
        10'b1001001101: data <= 11'h7ff; 
        10'b1001001110: data <= 11'h000; 
        10'b1001001111: data <= 11'h7ff; 
        10'b1001010000: data <= 11'h7ff; 
        10'b1001010001: data <= 11'h001; 
        10'b1001010010: data <= 11'h003; 
        10'b1001010011: data <= 11'h006; 
        10'b1001010100: data <= 11'h004; 
        10'b1001010101: data <= 11'h004; 
        10'b1001010110: data <= 11'h008; 
        10'b1001010111: data <= 11'h009; 
        10'b1001011000: data <= 11'h006; 
        10'b1001011001: data <= 11'h002; 
        10'b1001011010: data <= 11'h001; 
        10'b1001011011: data <= 11'h000; 
        10'b1001011100: data <= 11'h000; 
        10'b1001011101: data <= 11'h7fd; 
        10'b1001011110: data <= 11'h7fe; 
        10'b1001011111: data <= 11'h7ff; 
        10'b1001100000: data <= 11'h001; 
        10'b1001100001: data <= 11'h000; 
        10'b1001100010: data <= 11'h7ff; 
        10'b1001100011: data <= 11'h7fe; 
        10'b1001100100: data <= 11'h000; 
        10'b1001100101: data <= 11'h7ff; 
        10'b1001100110: data <= 11'h7ff; 
        10'b1001100111: data <= 11'h7ff; 
        10'b1001101000: data <= 11'h7ff; 
        10'b1001101001: data <= 11'h000; 
        10'b1001101010: data <= 11'h000; 
        10'b1001101011: data <= 11'h7ff; 
        10'b1001101100: data <= 11'h7ff; 
        10'b1001101101: data <= 11'h000; 
        10'b1001101110: data <= 11'h003; 
        10'b1001101111: data <= 11'h002; 
        10'b1001110000: data <= 11'h006; 
        10'b1001110001: data <= 11'h005; 
        10'b1001110010: data <= 11'h006; 
        10'b1001110011: data <= 11'h007; 
        10'b1001110100: data <= 11'h006; 
        10'b1001110101: data <= 11'h007; 
        10'b1001110110: data <= 11'h003; 
        10'b1001110111: data <= 11'h003; 
        10'b1001111000: data <= 11'h002; 
        10'b1001111001: data <= 11'h7fe; 
        10'b1001111010: data <= 11'h7ff; 
        10'b1001111011: data <= 11'h000; 
        10'b1001111100: data <= 11'h7fe; 
        10'b1001111101: data <= 11'h7fe; 
        10'b1001111110: data <= 11'h7ff; 
        10'b1001111111: data <= 11'h7ff; 
        10'b1010000000: data <= 11'h000; 
        10'b1010000001: data <= 11'h7ff; 
        10'b1010000010: data <= 11'h7ff; 
        10'b1010000011: data <= 11'h000; 
        10'b1010000100: data <= 11'h7ff; 
        10'b1010000101: data <= 11'h000; 
        10'b1010000110: data <= 11'h000; 
        10'b1010000111: data <= 11'h7ff; 
        10'b1010001000: data <= 11'h7ff; 
        10'b1010001001: data <= 11'h000; 
        10'b1010001010: data <= 11'h000; 
        10'b1010001011: data <= 11'h002; 
        10'b1010001100: data <= 11'h002; 
        10'b1010001101: data <= 11'h006; 
        10'b1010001110: data <= 11'h007; 
        10'b1010001111: data <= 11'h009; 
        10'b1010010000: data <= 11'h008; 
        10'b1010010001: data <= 11'h005; 
        10'b1010010010: data <= 11'h004; 
        10'b1010010011: data <= 11'h002; 
        10'b1010010100: data <= 11'h001; 
        10'b1010010101: data <= 11'h000; 
        10'b1010010110: data <= 11'h7fd; 
        10'b1010010111: data <= 11'h7fc; 
        10'b1010011000: data <= 11'h7fd; 
        10'b1010011001: data <= 11'h7fe; 
        10'b1010011010: data <= 11'h7ff; 
        10'b1010011011: data <= 11'h000; 
        10'b1010011100: data <= 11'h000; 
        10'b1010011101: data <= 11'h000; 
        10'b1010011110: data <= 11'h7ff; 
        10'b1010011111: data <= 11'h7ff; 
        10'b1010100000: data <= 11'h7ff; 
        10'b1010100001: data <= 11'h000; 
        10'b1010100010: data <= 11'h7ff; 
        10'b1010100011: data <= 11'h000; 
        10'b1010100100: data <= 11'h000; 
        10'b1010100101: data <= 11'h000; 
        10'b1010100110: data <= 11'h7fe; 
        10'b1010100111: data <= 11'h7fe; 
        10'b1010101000: data <= 11'h7ff; 
        10'b1010101001: data <= 11'h7ff; 
        10'b1010101010: data <= 11'h001; 
        10'b1010101011: data <= 11'h001; 
        10'b1010101100: data <= 11'h002; 
        10'b1010101101: data <= 11'h003; 
        10'b1010101110: data <= 11'h002; 
        10'b1010101111: data <= 11'h7ff; 
        10'b1010110000: data <= 11'h7fe; 
        10'b1010110001: data <= 11'h7fd; 
        10'b1010110010: data <= 11'h7fe; 
        10'b1010110011: data <= 11'h7fd; 
        10'b1010110100: data <= 11'h7fd; 
        10'b1010110101: data <= 11'h7fd; 
        10'b1010110110: data <= 11'h7ff; 
        10'b1010110111: data <= 11'h7ff; 
        10'b1010111000: data <= 11'h7ff; 
        10'b1010111001: data <= 11'h7ff; 
        10'b1010111010: data <= 11'h000; 
        10'b1010111011: data <= 11'h7ff; 
        10'b1010111100: data <= 11'h7ff; 
        10'b1010111101: data <= 11'h001; 
        10'b1010111110: data <= 11'h000; 
        10'b1010111111: data <= 11'h001; 
        10'b1011000000: data <= 11'h001; 
        10'b1011000001: data <= 11'h000; 
        10'b1011000010: data <= 11'h7fe; 
        10'b1011000011: data <= 11'h7ff; 
        10'b1011000100: data <= 11'h7fd; 
        10'b1011000101: data <= 11'h7fd; 
        10'b1011000110: data <= 11'h7fd; 
        10'b1011000111: data <= 11'h7fc; 
        10'b1011001000: data <= 11'h7fb; 
        10'b1011001001: data <= 11'h7fb; 
        10'b1011001010: data <= 11'h7fb; 
        10'b1011001011: data <= 11'h7fb; 
        10'b1011001100: data <= 11'h7fb; 
        10'b1011001101: data <= 11'h7fd; 
        10'b1011001110: data <= 11'h7fe; 
        10'b1011001111: data <= 11'h7fe; 
        10'b1011010000: data <= 11'h7fe; 
        10'b1011010001: data <= 11'h7fe; 
        10'b1011010010: data <= 11'h7ff; 
        10'b1011010011: data <= 11'h001; 
        10'b1011010100: data <= 11'h000; 
        10'b1011010101: data <= 11'h7ff; 
        10'b1011010110: data <= 11'h7ff; 
        10'b1011010111: data <= 11'h000; 
        10'b1011011000: data <= 11'h001; 
        10'b1011011001: data <= 11'h001; 
        10'b1011011010: data <= 11'h7ff; 
        10'b1011011011: data <= 11'h000; 
        10'b1011011100: data <= 11'h7ff; 
        10'b1011011101: data <= 11'h7ff; 
        10'b1011011110: data <= 11'h7ff; 
        10'b1011011111: data <= 11'h000; 
        10'b1011100000: data <= 11'h7ff; 
        10'b1011100001: data <= 11'h7fe; 
        10'b1011100010: data <= 11'h7fe; 
        10'b1011100011: data <= 11'h7fe; 
        10'b1011100100: data <= 11'h7ff; 
        10'b1011100101: data <= 11'h7fe; 
        10'b1011100110: data <= 11'h7fe; 
        10'b1011100111: data <= 11'h7ff; 
        10'b1011101000: data <= 11'h7fe; 
        10'b1011101001: data <= 11'h7fe; 
        10'b1011101010: data <= 11'h7ff; 
        10'b1011101011: data <= 11'h7fe; 
        10'b1011101100: data <= 11'h7ff; 
        10'b1011101101: data <= 11'h7fe; 
        10'b1011101110: data <= 11'h7fe; 
        10'b1011101111: data <= 11'h001; 
        10'b1011110000: data <= 11'h7ff; 
        10'b1011110001: data <= 11'h000; 
        10'b1011110010: data <= 11'h001; 
        10'b1011110011: data <= 11'h000; 
        10'b1011110100: data <= 11'h7ff; 
        10'b1011110101: data <= 11'h000; 
        10'b1011110110: data <= 11'h000; 
        10'b1011110111: data <= 11'h7ff; 
        10'b1011111000: data <= 11'h001; 
        10'b1011111001: data <= 11'h000; 
        10'b1011111010: data <= 11'h000; 
        10'b1011111011: data <= 11'h7ff; 
        10'b1011111100: data <= 11'h001; 
        10'b1011111101: data <= 11'h001; 
        10'b1011111110: data <= 11'h000; 
        10'b1011111111: data <= 11'h000; 
        10'b1100000000: data <= 11'h000; 
        10'b1100000001: data <= 11'h7ff; 
        10'b1100000010: data <= 11'h000; 
        10'b1100000011: data <= 11'h7ff; 
        10'b1100000100: data <= 11'h000; 
        10'b1100000101: data <= 11'h7ff; 
        10'b1100000110: data <= 11'h000; 
        10'b1100000111: data <= 11'h7ff; 
        10'b1100001000: data <= 11'h7ff; 
        10'b1100001001: data <= 11'h7ff; 
        10'b1100001010: data <= 11'h7fe; 
        10'b1100001011: data <= 11'h000; 
        10'b1100001100: data <= 11'h000; 
        10'b1100001101: data <= 11'h7ff; 
        10'b1100001110: data <= 11'h7ff; 
        10'b1100001111: data <= 11'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 6) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 12'hffe; 
        10'b0000000001: data <= 12'h001; 
        10'b0000000010: data <= 12'hfff; 
        10'b0000000011: data <= 12'h000; 
        10'b0000000100: data <= 12'h001; 
        10'b0000000101: data <= 12'h000; 
        10'b0000000110: data <= 12'hfff; 
        10'b0000000111: data <= 12'hfff; 
        10'b0000001000: data <= 12'h000; 
        10'b0000001001: data <= 12'hfff; 
        10'b0000001010: data <= 12'h002; 
        10'b0000001011: data <= 12'h000; 
        10'b0000001100: data <= 12'h001; 
        10'b0000001101: data <= 12'hffe; 
        10'b0000001110: data <= 12'h000; 
        10'b0000001111: data <= 12'hffd; 
        10'b0000010000: data <= 12'hffe; 
        10'b0000010001: data <= 12'hfff; 
        10'b0000010010: data <= 12'hffe; 
        10'b0000010011: data <= 12'h002; 
        10'b0000010100: data <= 12'hffe; 
        10'b0000010101: data <= 12'hfff; 
        10'b0000010110: data <= 12'hffe; 
        10'b0000010111: data <= 12'h000; 
        10'b0000011000: data <= 12'h001; 
        10'b0000011001: data <= 12'hfff; 
        10'b0000011010: data <= 12'h000; 
        10'b0000011011: data <= 12'h000; 
        10'b0000011100: data <= 12'h001; 
        10'b0000011101: data <= 12'h001; 
        10'b0000011110: data <= 12'h000; 
        10'b0000011111: data <= 12'hffe; 
        10'b0000100000: data <= 12'hffd; 
        10'b0000100001: data <= 12'h000; 
        10'b0000100010: data <= 12'hffe; 
        10'b0000100011: data <= 12'hfff; 
        10'b0000100100: data <= 12'hffe; 
        10'b0000100101: data <= 12'hffd; 
        10'b0000100110: data <= 12'hffe; 
        10'b0000100111: data <= 12'h000; 
        10'b0000101000: data <= 12'h002; 
        10'b0000101001: data <= 12'hffe; 
        10'b0000101010: data <= 12'hfff; 
        10'b0000101011: data <= 12'h001; 
        10'b0000101100: data <= 12'hffe; 
        10'b0000101101: data <= 12'hffd; 
        10'b0000101110: data <= 12'h001; 
        10'b0000101111: data <= 12'h001; 
        10'b0000110000: data <= 12'hffe; 
        10'b0000110001: data <= 12'h001; 
        10'b0000110010: data <= 12'hffe; 
        10'b0000110011: data <= 12'hffe; 
        10'b0000110100: data <= 12'h000; 
        10'b0000110101: data <= 12'h000; 
        10'b0000110110: data <= 12'hfff; 
        10'b0000110111: data <= 12'h001; 
        10'b0000111000: data <= 12'hffd; 
        10'b0000111001: data <= 12'hffe; 
        10'b0000111010: data <= 12'hffe; 
        10'b0000111011: data <= 12'h001; 
        10'b0000111100: data <= 12'h000; 
        10'b0000111101: data <= 12'hffd; 
        10'b0000111110: data <= 12'hfff; 
        10'b0000111111: data <= 12'h001; 
        10'b0001000000: data <= 12'hfff; 
        10'b0001000001: data <= 12'hffe; 
        10'b0001000010: data <= 12'hffe; 
        10'b0001000011: data <= 12'hffd; 
        10'b0001000100: data <= 12'hffd; 
        10'b0001000101: data <= 12'hfff; 
        10'b0001000110: data <= 12'hffd; 
        10'b0001000111: data <= 12'hffc; 
        10'b0001001000: data <= 12'hffd; 
        10'b0001001001: data <= 12'hfff; 
        10'b0001001010: data <= 12'hffd; 
        10'b0001001011: data <= 12'hffc; 
        10'b0001001100: data <= 12'hfff; 
        10'b0001001101: data <= 12'h001; 
        10'b0001001110: data <= 12'h000; 
        10'b0001001111: data <= 12'hffe; 
        10'b0001010000: data <= 12'h001; 
        10'b0001010001: data <= 12'hffd; 
        10'b0001010010: data <= 12'hfff; 
        10'b0001010011: data <= 12'h001; 
        10'b0001010100: data <= 12'hffd; 
        10'b0001010101: data <= 12'hfff; 
        10'b0001010110: data <= 12'h002; 
        10'b0001010111: data <= 12'hffd; 
        10'b0001011000: data <= 12'hffe; 
        10'b0001011001: data <= 12'h001; 
        10'b0001011010: data <= 12'h000; 
        10'b0001011011: data <= 12'h000; 
        10'b0001011100: data <= 12'h000; 
        10'b0001011101: data <= 12'hfff; 
        10'b0001011110: data <= 12'hfff; 
        10'b0001011111: data <= 12'hffc; 
        10'b0001100000: data <= 12'hffb; 
        10'b0001100001: data <= 12'hffd; 
        10'b0001100010: data <= 12'hffc; 
        10'b0001100011: data <= 12'hffc; 
        10'b0001100100: data <= 12'h001; 
        10'b0001100101: data <= 12'h000; 
        10'b0001100110: data <= 12'hffb; 
        10'b0001100111: data <= 12'hffc; 
        10'b0001101000: data <= 12'hffa; 
        10'b0001101001: data <= 12'hffc; 
        10'b0001101010: data <= 12'hffb; 
        10'b0001101011: data <= 12'hffd; 
        10'b0001101100: data <= 12'hffe; 
        10'b0001101101: data <= 12'h001; 
        10'b0001101110: data <= 12'h001; 
        10'b0001101111: data <= 12'hfff; 
        10'b0001110000: data <= 12'h000; 
        10'b0001110001: data <= 12'hffd; 
        10'b0001110010: data <= 12'hffe; 
        10'b0001110011: data <= 12'hffd; 
        10'b0001110100: data <= 12'hffd; 
        10'b0001110101: data <= 12'h000; 
        10'b0001110110: data <= 12'hfff; 
        10'b0001110111: data <= 12'hffd; 
        10'b0001111000: data <= 12'hfff; 
        10'b0001111001: data <= 12'hfff; 
        10'b0001111010: data <= 12'hffc; 
        10'b0001111011: data <= 12'hffc; 
        10'b0001111100: data <= 12'hffc; 
        10'b0001111101: data <= 12'hffc; 
        10'b0001111110: data <= 12'hfff; 
        10'b0001111111: data <= 12'h000; 
        10'b0010000000: data <= 12'hffd; 
        10'b0010000001: data <= 12'hffd; 
        10'b0010000010: data <= 12'hffd; 
        10'b0010000011: data <= 12'hffc; 
        10'b0010000100: data <= 12'hffe; 
        10'b0010000101: data <= 12'hffa; 
        10'b0010000110: data <= 12'hffe; 
        10'b0010000111: data <= 12'h000; 
        10'b0010001000: data <= 12'hffd; 
        10'b0010001001: data <= 12'hfff; 
        10'b0010001010: data <= 12'hfff; 
        10'b0010001011: data <= 12'h000; 
        10'b0010001100: data <= 12'h001; 
        10'b0010001101: data <= 12'hfff; 
        10'b0010001110: data <= 12'h000; 
        10'b0010001111: data <= 12'hffe; 
        10'b0010010000: data <= 12'hfff; 
        10'b0010010001: data <= 12'hfff; 
        10'b0010010010: data <= 12'hfff; 
        10'b0010010011: data <= 12'hffe; 
        10'b0010010100: data <= 12'hfff; 
        10'b0010010101: data <= 12'hffd; 
        10'b0010010110: data <= 12'hfff; 
        10'b0010010111: data <= 12'h001; 
        10'b0010011000: data <= 12'h004; 
        10'b0010011001: data <= 12'h008; 
        10'b0010011010: data <= 12'h00a; 
        10'b0010011011: data <= 12'h00a; 
        10'b0010011100: data <= 12'h00b; 
        10'b0010011101: data <= 12'h00c; 
        10'b0010011110: data <= 12'h00c; 
        10'b0010011111: data <= 12'h004; 
        10'b0010100000: data <= 12'h001; 
        10'b0010100001: data <= 12'h002; 
        10'b0010100010: data <= 12'hfff; 
        10'b0010100011: data <= 12'h000; 
        10'b0010100100: data <= 12'hffb; 
        10'b0010100101: data <= 12'hffc; 
        10'b0010100110: data <= 12'h000; 
        10'b0010100111: data <= 12'hffe; 
        10'b0010101000: data <= 12'hfff; 
        10'b0010101001: data <= 12'hfff; 
        10'b0010101010: data <= 12'h000; 
        10'b0010101011: data <= 12'hfff; 
        10'b0010101100: data <= 12'h000; 
        10'b0010101101: data <= 12'h000; 
        10'b0010101110: data <= 12'h000; 
        10'b0010101111: data <= 12'h000; 
        10'b0010110000: data <= 12'hffd; 
        10'b0010110001: data <= 12'hffb; 
        10'b0010110010: data <= 12'h002; 
        10'b0010110011: data <= 12'h000; 
        10'b0010110100: data <= 12'h007; 
        10'b0010110101: data <= 12'h006; 
        10'b0010110110: data <= 12'h006; 
        10'b0010110111: data <= 12'h008; 
        10'b0010111000: data <= 12'h00a; 
        10'b0010111001: data <= 12'h00f; 
        10'b0010111010: data <= 12'h00e; 
        10'b0010111011: data <= 12'h00c; 
        10'b0010111100: data <= 12'h00b; 
        10'b0010111101: data <= 12'h00d; 
        10'b0010111110: data <= 12'h007; 
        10'b0010111111: data <= 12'h003; 
        10'b0011000000: data <= 12'hffa; 
        10'b0011000001: data <= 12'hffa; 
        10'b0011000010: data <= 12'hffc; 
        10'b0011000011: data <= 12'h001; 
        10'b0011000100: data <= 12'h001; 
        10'b0011000101: data <= 12'h000; 
        10'b0011000110: data <= 12'h000; 
        10'b0011000111: data <= 12'hffd; 
        10'b0011001000: data <= 12'hffb; 
        10'b0011001001: data <= 12'h000; 
        10'b0011001010: data <= 12'hffe; 
        10'b0011001011: data <= 12'h000; 
        10'b0011001100: data <= 12'hffe; 
        10'b0011001101: data <= 12'hfff; 
        10'b0011001110: data <= 12'h000; 
        10'b0011001111: data <= 12'h005; 
        10'b0011010000: data <= 12'h00a; 
        10'b0011010001: data <= 12'h009; 
        10'b0011010010: data <= 12'h004; 
        10'b0011010011: data <= 12'h006; 
        10'b0011010100: data <= 12'h008; 
        10'b0011010101: data <= 12'h010; 
        10'b0011010110: data <= 12'h00c; 
        10'b0011010111: data <= 12'h00a; 
        10'b0011011000: data <= 12'h004; 
        10'b0011011001: data <= 12'h008; 
        10'b0011011010: data <= 12'h009; 
        10'b0011011011: data <= 12'h004; 
        10'b0011011100: data <= 12'hffd; 
        10'b0011011101: data <= 12'hffa; 
        10'b0011011110: data <= 12'hffb; 
        10'b0011011111: data <= 12'h000; 
        10'b0011100000: data <= 12'h002; 
        10'b0011100001: data <= 12'h001; 
        10'b0011100010: data <= 12'hfff; 
        10'b0011100011: data <= 12'h000; 
        10'b0011100100: data <= 12'hffc; 
        10'b0011100101: data <= 12'hffd; 
        10'b0011100110: data <= 12'hffe; 
        10'b0011100111: data <= 12'hffd; 
        10'b0011101000: data <= 12'hffe; 
        10'b0011101001: data <= 12'hffe; 
        10'b0011101010: data <= 12'h005; 
        10'b0011101011: data <= 12'h005; 
        10'b0011101100: data <= 12'h003; 
        10'b0011101101: data <= 12'h001; 
        10'b0011101110: data <= 12'h002; 
        10'b0011101111: data <= 12'h007; 
        10'b0011110000: data <= 12'h015; 
        10'b0011110001: data <= 12'h010; 
        10'b0011110010: data <= 12'h00f; 
        10'b0011110011: data <= 12'h005; 
        10'b0011110100: data <= 12'h004; 
        10'b0011110101: data <= 12'h004; 
        10'b0011110110: data <= 12'h009; 
        10'b0011110111: data <= 12'h010; 
        10'b0011111000: data <= 12'hffe; 
        10'b0011111001: data <= 12'hffb; 
        10'b0011111010: data <= 12'hfff; 
        10'b0011111011: data <= 12'hffd; 
        10'b0011111100: data <= 12'h000; 
        10'b0011111101: data <= 12'h000; 
        10'b0011111110: data <= 12'h000; 
        10'b0011111111: data <= 12'h000; 
        10'b0100000000: data <= 12'hffb; 
        10'b0100000001: data <= 12'hffd; 
        10'b0100000010: data <= 12'hffb; 
        10'b0100000011: data <= 12'hffd; 
        10'b0100000100: data <= 12'hffd; 
        10'b0100000101: data <= 12'hfff; 
        10'b0100000110: data <= 12'h003; 
        10'b0100000111: data <= 12'hffd; 
        10'b0100001000: data <= 12'h002; 
        10'b0100001001: data <= 12'h005; 
        10'b0100001010: data <= 12'h005; 
        10'b0100001011: data <= 12'h004; 
        10'b0100001100: data <= 12'h00b; 
        10'b0100001101: data <= 12'h00f; 
        10'b0100001110: data <= 12'h011; 
        10'b0100001111: data <= 12'h00a; 
        10'b0100010000: data <= 12'h003; 
        10'b0100010001: data <= 12'hfff; 
        10'b0100010010: data <= 12'h007; 
        10'b0100010011: data <= 12'h010; 
        10'b0100010100: data <= 12'h005; 
        10'b0100010101: data <= 12'hffc; 
        10'b0100010110: data <= 12'h000; 
        10'b0100010111: data <= 12'h000; 
        10'b0100011000: data <= 12'hffd; 
        10'b0100011001: data <= 12'h001; 
        10'b0100011010: data <= 12'hffe; 
        10'b0100011011: data <= 12'hffc; 
        10'b0100011100: data <= 12'hffc; 
        10'b0100011101: data <= 12'hffd; 
        10'b0100011110: data <= 12'hffe; 
        10'b0100011111: data <= 12'h000; 
        10'b0100100000: data <= 12'h002; 
        10'b0100100001: data <= 12'h000; 
        10'b0100100010: data <= 12'hffd; 
        10'b0100100011: data <= 12'h001; 
        10'b0100100100: data <= 12'h001; 
        10'b0100100101: data <= 12'hfff; 
        10'b0100100110: data <= 12'hffb; 
        10'b0100100111: data <= 12'hff7; 
        10'b0100101000: data <= 12'hffa; 
        10'b0100101001: data <= 12'h005; 
        10'b0100101010: data <= 12'h00e; 
        10'b0100101011: data <= 12'h00e; 
        10'b0100101100: data <= 12'h00d; 
        10'b0100101101: data <= 12'h009; 
        10'b0100101110: data <= 12'h00e; 
        10'b0100101111: data <= 12'h013; 
        10'b0100110000: data <= 12'h009; 
        10'b0100110001: data <= 12'hffc; 
        10'b0100110010: data <= 12'hffc; 
        10'b0100110011: data <= 12'hffd; 
        10'b0100110100: data <= 12'hffe; 
        10'b0100110101: data <= 12'hffd; 
        10'b0100110110: data <= 12'h001; 
        10'b0100110111: data <= 12'hfff; 
        10'b0100111000: data <= 12'hff9; 
        10'b0100111001: data <= 12'hfff; 
        10'b0100111010: data <= 12'h001; 
        10'b0100111011: data <= 12'h005; 
        10'b0100111100: data <= 12'h004; 
        10'b0100111101: data <= 12'hffe; 
        10'b0100111110: data <= 12'h001; 
        10'b0100111111: data <= 12'h000; 
        10'b0101000000: data <= 12'h003; 
        10'b0101000001: data <= 12'hffe; 
        10'b0101000010: data <= 12'hff1; 
        10'b0101000011: data <= 12'hfe5; 
        10'b0101000100: data <= 12'hfe6; 
        10'b0101000101: data <= 12'hff6; 
        10'b0101000110: data <= 12'hfff; 
        10'b0101000111: data <= 12'h007; 
        10'b0101001000: data <= 12'h00c; 
        10'b0101001001: data <= 12'h00b; 
        10'b0101001010: data <= 12'h00f; 
        10'b0101001011: data <= 12'h011; 
        10'b0101001100: data <= 12'h00c; 
        10'b0101001101: data <= 12'hffe; 
        10'b0101001110: data <= 12'h000; 
        10'b0101001111: data <= 12'hffd; 
        10'b0101010000: data <= 12'hffe; 
        10'b0101010001: data <= 12'hfff; 
        10'b0101010010: data <= 12'hfff; 
        10'b0101010011: data <= 12'hfff; 
        10'b0101010100: data <= 12'hffc; 
        10'b0101010101: data <= 12'h001; 
        10'b0101010110: data <= 12'h006; 
        10'b0101010111: data <= 12'h006; 
        10'b0101011000: data <= 12'h003; 
        10'b0101011001: data <= 12'hfff; 
        10'b0101011010: data <= 12'h004; 
        10'b0101011011: data <= 12'h003; 
        10'b0101011100: data <= 12'h005; 
        10'b0101011101: data <= 12'hffc; 
        10'b0101011110: data <= 12'hfe3; 
        10'b0101011111: data <= 12'hfdc; 
        10'b0101100000: data <= 12'hfdc; 
        10'b0101100001: data <= 12'hfec; 
        10'b0101100010: data <= 12'hffd; 
        10'b0101100011: data <= 12'hfff; 
        10'b0101100100: data <= 12'h002; 
        10'b0101100101: data <= 12'h005; 
        10'b0101100110: data <= 12'h013; 
        10'b0101100111: data <= 12'h011; 
        10'b0101101000: data <= 12'h00c; 
        10'b0101101001: data <= 12'h000; 
        10'b0101101010: data <= 12'hffe; 
        10'b0101101011: data <= 12'hffe; 
        10'b0101101100: data <= 12'hffd; 
        10'b0101101101: data <= 12'h000; 
        10'b0101101110: data <= 12'h001; 
        10'b0101101111: data <= 12'hffd; 
        10'b0101110000: data <= 12'hfff; 
        10'b0101110001: data <= 12'h004; 
        10'b0101110010: data <= 12'h007; 
        10'b0101110011: data <= 12'h009; 
        10'b0101110100: data <= 12'h007; 
        10'b0101110101: data <= 12'h005; 
        10'b0101110110: data <= 12'h006; 
        10'b0101110111: data <= 12'h005; 
        10'b0101111000: data <= 12'h004; 
        10'b0101111001: data <= 12'hfee; 
        10'b0101111010: data <= 12'hfe3; 
        10'b0101111011: data <= 12'hfdb; 
        10'b0101111100: data <= 12'hfe2; 
        10'b0101111101: data <= 12'hff1; 
        10'b0101111110: data <= 12'hff9; 
        10'b0101111111: data <= 12'hff6; 
        10'b0110000000: data <= 12'hff8; 
        10'b0110000001: data <= 12'h003; 
        10'b0110000010: data <= 12'h00c; 
        10'b0110000011: data <= 12'h014; 
        10'b0110000100: data <= 12'h00b; 
        10'b0110000101: data <= 12'h002; 
        10'b0110000110: data <= 12'h000; 
        10'b0110000111: data <= 12'h001; 
        10'b0110001000: data <= 12'h000; 
        10'b0110001001: data <= 12'h001; 
        10'b0110001010: data <= 12'hffe; 
        10'b0110001011: data <= 12'hffe; 
        10'b0110001100: data <= 12'hffd; 
        10'b0110001101: data <= 12'h009; 
        10'b0110001110: data <= 12'h00c; 
        10'b0110001111: data <= 12'h00e; 
        10'b0110010000: data <= 12'h007; 
        10'b0110010001: data <= 12'h008; 
        10'b0110010010: data <= 12'h00c; 
        10'b0110010011: data <= 12'h007; 
        10'b0110010100: data <= 12'h002; 
        10'b0110010101: data <= 12'hff1; 
        10'b0110010110: data <= 12'hfde; 
        10'b0110010111: data <= 12'hfdb; 
        10'b0110011000: data <= 12'hfe3; 
        10'b0110011001: data <= 12'hff0; 
        10'b0110011010: data <= 12'hff9; 
        10'b0110011011: data <= 12'hff7; 
        10'b0110011100: data <= 12'h001; 
        10'b0110011101: data <= 12'h007; 
        10'b0110011110: data <= 12'h008; 
        10'b0110011111: data <= 12'h014; 
        10'b0110100000: data <= 12'h00a; 
        10'b0110100001: data <= 12'hffe; 
        10'b0110100010: data <= 12'hfff; 
        10'b0110100011: data <= 12'hffe; 
        10'b0110100100: data <= 12'h001; 
        10'b0110100101: data <= 12'h001; 
        10'b0110100110: data <= 12'hffe; 
        10'b0110100111: data <= 12'h000; 
        10'b0110101000: data <= 12'h000; 
        10'b0110101001: data <= 12'h00d; 
        10'b0110101010: data <= 12'h009; 
        10'b0110101011: data <= 12'h00d; 
        10'b0110101100: data <= 12'h009; 
        10'b0110101101: data <= 12'h00c; 
        10'b0110101110: data <= 12'h00f; 
        10'b0110101111: data <= 12'h004; 
        10'b0110110000: data <= 12'hff5; 
        10'b0110110001: data <= 12'hfe3; 
        10'b0110110010: data <= 12'hfda; 
        10'b0110110011: data <= 12'hfdb; 
        10'b0110110100: data <= 12'hfe7; 
        10'b0110110101: data <= 12'hff4; 
        10'b0110110110: data <= 12'hffc; 
        10'b0110110111: data <= 12'hffc; 
        10'b0110111000: data <= 12'h004; 
        10'b0110111001: data <= 12'h003; 
        10'b0110111010: data <= 12'h00d; 
        10'b0110111011: data <= 12'h00f; 
        10'b0110111100: data <= 12'h008; 
        10'b0110111101: data <= 12'hfff; 
        10'b0110111110: data <= 12'h000; 
        10'b0110111111: data <= 12'hffe; 
        10'b0111000000: data <= 12'h000; 
        10'b0111000001: data <= 12'h001; 
        10'b0111000010: data <= 12'hffd; 
        10'b0111000011: data <= 12'hffe; 
        10'b0111000100: data <= 12'h002; 
        10'b0111000101: data <= 12'h00c; 
        10'b0111000110: data <= 12'h00f; 
        10'b0111000111: data <= 12'h00b; 
        10'b0111001000: data <= 12'h008; 
        10'b0111001001: data <= 12'h008; 
        10'b0111001010: data <= 12'h00d; 
        10'b0111001011: data <= 12'hffe; 
        10'b0111001100: data <= 12'hfea; 
        10'b0111001101: data <= 12'hfda; 
        10'b0111001110: data <= 12'hfdb; 
        10'b0111001111: data <= 12'hfe3; 
        10'b0111010000: data <= 12'hff0; 
        10'b0111010001: data <= 12'hff9; 
        10'b0111010010: data <= 12'h000; 
        10'b0111010011: data <= 12'h002; 
        10'b0111010100: data <= 12'h006; 
        10'b0111010101: data <= 12'h008; 
        10'b0111010110: data <= 12'h00b; 
        10'b0111010111: data <= 12'h00b; 
        10'b0111011000: data <= 12'h004; 
        10'b0111011001: data <= 12'h000; 
        10'b0111011010: data <= 12'hfff; 
        10'b0111011011: data <= 12'hffe; 
        10'b0111011100: data <= 12'hfff; 
        10'b0111011101: data <= 12'h000; 
        10'b0111011110: data <= 12'hffe; 
        10'b0111011111: data <= 12'hffb; 
        10'b0111100000: data <= 12'h000; 
        10'b0111100001: data <= 12'h008; 
        10'b0111100010: data <= 12'h00a; 
        10'b0111100011: data <= 12'h00a; 
        10'b0111100100: data <= 12'h003; 
        10'b0111100101: data <= 12'h008; 
        10'b0111100110: data <= 12'h00d; 
        10'b0111100111: data <= 12'hffe; 
        10'b0111101000: data <= 12'hfe6; 
        10'b0111101001: data <= 12'hfda; 
        10'b0111101010: data <= 12'hfdf; 
        10'b0111101011: data <= 12'hfec; 
        10'b0111101100: data <= 12'hffd; 
        10'b0111101101: data <= 12'h005; 
        10'b0111101110: data <= 12'h007; 
        10'b0111101111: data <= 12'h007; 
        10'b0111110000: data <= 12'h009; 
        10'b0111110001: data <= 12'h006; 
        10'b0111110010: data <= 12'h005; 
        10'b0111110011: data <= 12'h006; 
        10'b0111110100: data <= 12'h000; 
        10'b0111110101: data <= 12'hfff; 
        10'b0111110110: data <= 12'h000; 
        10'b0111110111: data <= 12'hffe; 
        10'b0111111000: data <= 12'hfff; 
        10'b0111111001: data <= 12'h000; 
        10'b0111111010: data <= 12'hfff; 
        10'b0111111011: data <= 12'hffe; 
        10'b0111111100: data <= 12'hfff; 
        10'b0111111101: data <= 12'h005; 
        10'b0111111110: data <= 12'h00b; 
        10'b0111111111: data <= 12'h006; 
        10'b1000000000: data <= 12'h004; 
        10'b1000000001: data <= 12'h00b; 
        10'b1000000010: data <= 12'h015; 
        10'b1000000011: data <= 12'h001; 
        10'b1000000100: data <= 12'hfef; 
        10'b1000000101: data <= 12'hfe5; 
        10'b1000000110: data <= 12'hfed; 
        10'b1000000111: data <= 12'hffa; 
        10'b1000001000: data <= 12'h006; 
        10'b1000001001: data <= 12'h006; 
        10'b1000001010: data <= 12'h007; 
        10'b1000001011: data <= 12'h004; 
        10'b1000001100: data <= 12'h002; 
        10'b1000001101: data <= 12'h003; 
        10'b1000001110: data <= 12'h006; 
        10'b1000001111: data <= 12'h004; 
        10'b1000010000: data <= 12'h000; 
        10'b1000010001: data <= 12'hffe; 
        10'b1000010010: data <= 12'h000; 
        10'b1000010011: data <= 12'hfff; 
        10'b1000010100: data <= 12'hfff; 
        10'b1000010101: data <= 12'hfff; 
        10'b1000010110: data <= 12'hfff; 
        10'b1000010111: data <= 12'hffb; 
        10'b1000011000: data <= 12'h002; 
        10'b1000011001: data <= 12'h006; 
        10'b1000011010: data <= 12'h00e; 
        10'b1000011011: data <= 12'h00d; 
        10'b1000011100: data <= 12'h00a; 
        10'b1000011101: data <= 12'h00d; 
        10'b1000011110: data <= 12'h015; 
        10'b1000011111: data <= 12'h00f; 
        10'b1000100000: data <= 12'h003; 
        10'b1000100001: data <= 12'hff9; 
        10'b1000100010: data <= 12'hffd; 
        10'b1000100011: data <= 12'hffe; 
        10'b1000100100: data <= 12'h003; 
        10'b1000100101: data <= 12'hfff; 
        10'b1000100110: data <= 12'hffd; 
        10'b1000100111: data <= 12'hffe; 
        10'b1000101000: data <= 12'h003; 
        10'b1000101001: data <= 12'h003; 
        10'b1000101010: data <= 12'h006; 
        10'b1000101011: data <= 12'hfff; 
        10'b1000101100: data <= 12'h001; 
        10'b1000101101: data <= 12'hfff; 
        10'b1000101110: data <= 12'hffd; 
        10'b1000101111: data <= 12'h001; 
        10'b1000110000: data <= 12'h001; 
        10'b1000110001: data <= 12'h001; 
        10'b1000110010: data <= 12'hfff; 
        10'b1000110011: data <= 12'hffe; 
        10'b1000110100: data <= 12'hfff; 
        10'b1000110101: data <= 12'h006; 
        10'b1000110110: data <= 12'h00b; 
        10'b1000110111: data <= 12'h008; 
        10'b1000111000: data <= 12'h00a; 
        10'b1000111001: data <= 12'h00d; 
        10'b1000111010: data <= 12'h014; 
        10'b1000111011: data <= 12'h014; 
        10'b1000111100: data <= 12'h00a; 
        10'b1000111101: data <= 12'h003; 
        10'b1000111110: data <= 12'hffe; 
        10'b1000111111: data <= 12'h001; 
        10'b1001000000: data <= 12'h001; 
        10'b1001000001: data <= 12'hffd; 
        10'b1001000010: data <= 12'hffe; 
        10'b1001000011: data <= 12'hffd; 
        10'b1001000100: data <= 12'h002; 
        10'b1001000101: data <= 12'h002; 
        10'b1001000110: data <= 12'h003; 
        10'b1001000111: data <= 12'h001; 
        10'b1001001000: data <= 12'hffe; 
        10'b1001001001: data <= 12'h000; 
        10'b1001001010: data <= 12'hffe; 
        10'b1001001011: data <= 12'hfff; 
        10'b1001001100: data <= 12'hffe; 
        10'b1001001101: data <= 12'hffd; 
        10'b1001001110: data <= 12'hfff; 
        10'b1001001111: data <= 12'hffe; 
        10'b1001010000: data <= 12'hfff; 
        10'b1001010001: data <= 12'h002; 
        10'b1001010010: data <= 12'h007; 
        10'b1001010011: data <= 12'h00b; 
        10'b1001010100: data <= 12'h008; 
        10'b1001010101: data <= 12'h009; 
        10'b1001010110: data <= 12'h011; 
        10'b1001010111: data <= 12'h013; 
        10'b1001011000: data <= 12'h00d; 
        10'b1001011001: data <= 12'h005; 
        10'b1001011010: data <= 12'h002; 
        10'b1001011011: data <= 12'h000; 
        10'b1001011100: data <= 12'h000; 
        10'b1001011101: data <= 12'hffb; 
        10'b1001011110: data <= 12'hffc; 
        10'b1001011111: data <= 12'hffe; 
        10'b1001100000: data <= 12'h002; 
        10'b1001100001: data <= 12'h000; 
        10'b1001100010: data <= 12'hffe; 
        10'b1001100011: data <= 12'hffc; 
        10'b1001100100: data <= 12'hfff; 
        10'b1001100101: data <= 12'hfff; 
        10'b1001100110: data <= 12'hffe; 
        10'b1001100111: data <= 12'hffe; 
        10'b1001101000: data <= 12'hffe; 
        10'b1001101001: data <= 12'h000; 
        10'b1001101010: data <= 12'h000; 
        10'b1001101011: data <= 12'hfff; 
        10'b1001101100: data <= 12'hffe; 
        10'b1001101101: data <= 12'h001; 
        10'b1001101110: data <= 12'h005; 
        10'b1001101111: data <= 12'h004; 
        10'b1001110000: data <= 12'h00d; 
        10'b1001110001: data <= 12'h00a; 
        10'b1001110010: data <= 12'h00b; 
        10'b1001110011: data <= 12'h00d; 
        10'b1001110100: data <= 12'h00b; 
        10'b1001110101: data <= 12'h00f; 
        10'b1001110110: data <= 12'h006; 
        10'b1001110111: data <= 12'h007; 
        10'b1001111000: data <= 12'h004; 
        10'b1001111001: data <= 12'hffd; 
        10'b1001111010: data <= 12'hffe; 
        10'b1001111011: data <= 12'h000; 
        10'b1001111100: data <= 12'hffd; 
        10'b1001111101: data <= 12'hffc; 
        10'b1001111110: data <= 12'hffe; 
        10'b1001111111: data <= 12'hffe; 
        10'b1010000000: data <= 12'hfff; 
        10'b1010000001: data <= 12'hfff; 
        10'b1010000010: data <= 12'hfff; 
        10'b1010000011: data <= 12'hfff; 
        10'b1010000100: data <= 12'hffe; 
        10'b1010000101: data <= 12'hfff; 
        10'b1010000110: data <= 12'h000; 
        10'b1010000111: data <= 12'hffd; 
        10'b1010001000: data <= 12'hffd; 
        10'b1010001001: data <= 12'hfff; 
        10'b1010001010: data <= 12'h000; 
        10'b1010001011: data <= 12'h003; 
        10'b1010001100: data <= 12'h005; 
        10'b1010001101: data <= 12'h00c; 
        10'b1010001110: data <= 12'h00e; 
        10'b1010001111: data <= 12'h011; 
        10'b1010010000: data <= 12'h011; 
        10'b1010010001: data <= 12'h00a; 
        10'b1010010010: data <= 12'h008; 
        10'b1010010011: data <= 12'h005; 
        10'b1010010100: data <= 12'h002; 
        10'b1010010101: data <= 12'h000; 
        10'b1010010110: data <= 12'hffa; 
        10'b1010010111: data <= 12'hff8; 
        10'b1010011000: data <= 12'hffa; 
        10'b1010011001: data <= 12'hffd; 
        10'b1010011010: data <= 12'hffd; 
        10'b1010011011: data <= 12'h000; 
        10'b1010011100: data <= 12'hfff; 
        10'b1010011101: data <= 12'h001; 
        10'b1010011110: data <= 12'hfff; 
        10'b1010011111: data <= 12'hffd; 
        10'b1010100000: data <= 12'hfff; 
        10'b1010100001: data <= 12'hfff; 
        10'b1010100010: data <= 12'hffd; 
        10'b1010100011: data <= 12'h000; 
        10'b1010100100: data <= 12'hfff; 
        10'b1010100101: data <= 12'hfff; 
        10'b1010100110: data <= 12'hffd; 
        10'b1010100111: data <= 12'hffc; 
        10'b1010101000: data <= 12'hffe; 
        10'b1010101001: data <= 12'hffe; 
        10'b1010101010: data <= 12'h003; 
        10'b1010101011: data <= 12'h002; 
        10'b1010101100: data <= 12'h005; 
        10'b1010101101: data <= 12'h007; 
        10'b1010101110: data <= 12'h004; 
        10'b1010101111: data <= 12'hffd; 
        10'b1010110000: data <= 12'hffc; 
        10'b1010110001: data <= 12'hffb; 
        10'b1010110010: data <= 12'hffc; 
        10'b1010110011: data <= 12'hffa; 
        10'b1010110100: data <= 12'hffa; 
        10'b1010110101: data <= 12'hffa; 
        10'b1010110110: data <= 12'hfff; 
        10'b1010110111: data <= 12'hfff; 
        10'b1010111000: data <= 12'hffe; 
        10'b1010111001: data <= 12'hffe; 
        10'b1010111010: data <= 12'h000; 
        10'b1010111011: data <= 12'hffe; 
        10'b1010111100: data <= 12'hffe; 
        10'b1010111101: data <= 12'h002; 
        10'b1010111110: data <= 12'hfff; 
        10'b1010111111: data <= 12'h001; 
        10'b1011000000: data <= 12'h002; 
        10'b1011000001: data <= 12'h000; 
        10'b1011000010: data <= 12'hffd; 
        10'b1011000011: data <= 12'hfff; 
        10'b1011000100: data <= 12'hffa; 
        10'b1011000101: data <= 12'hffa; 
        10'b1011000110: data <= 12'hff9; 
        10'b1011000111: data <= 12'hff7; 
        10'b1011001000: data <= 12'hff6; 
        10'b1011001001: data <= 12'hff7; 
        10'b1011001010: data <= 12'hff5; 
        10'b1011001011: data <= 12'hff6; 
        10'b1011001100: data <= 12'hff7; 
        10'b1011001101: data <= 12'hffa; 
        10'b1011001110: data <= 12'hffb; 
        10'b1011001111: data <= 12'hffc; 
        10'b1011010000: data <= 12'hffc; 
        10'b1011010001: data <= 12'hffc; 
        10'b1011010010: data <= 12'hfff; 
        10'b1011010011: data <= 12'h001; 
        10'b1011010100: data <= 12'h001; 
        10'b1011010101: data <= 12'hfff; 
        10'b1011010110: data <= 12'hfff; 
        10'b1011010111: data <= 12'hfff; 
        10'b1011011000: data <= 12'h001; 
        10'b1011011001: data <= 12'h001; 
        10'b1011011010: data <= 12'hfff; 
        10'b1011011011: data <= 12'h000; 
        10'b1011011100: data <= 12'hffe; 
        10'b1011011101: data <= 12'hfff; 
        10'b1011011110: data <= 12'hffd; 
        10'b1011011111: data <= 12'h001; 
        10'b1011100000: data <= 12'hfff; 
        10'b1011100001: data <= 12'hffb; 
        10'b1011100010: data <= 12'hffb; 
        10'b1011100011: data <= 12'hffc; 
        10'b1011100100: data <= 12'hffe; 
        10'b1011100101: data <= 12'hffc; 
        10'b1011100110: data <= 12'hffc; 
        10'b1011100111: data <= 12'hffe; 
        10'b1011101000: data <= 12'hffc; 
        10'b1011101001: data <= 12'hffc; 
        10'b1011101010: data <= 12'hffd; 
        10'b1011101011: data <= 12'hffd; 
        10'b1011101100: data <= 12'hffe; 
        10'b1011101101: data <= 12'hffc; 
        10'b1011101110: data <= 12'hffd; 
        10'b1011101111: data <= 12'h001; 
        10'b1011110000: data <= 12'hffe; 
        10'b1011110001: data <= 12'h000; 
        10'b1011110010: data <= 12'h001; 
        10'b1011110011: data <= 12'h000; 
        10'b1011110100: data <= 12'hffe; 
        10'b1011110101: data <= 12'h001; 
        10'b1011110110: data <= 12'h000; 
        10'b1011110111: data <= 12'hfff; 
        10'b1011111000: data <= 12'h001; 
        10'b1011111001: data <= 12'h000; 
        10'b1011111010: data <= 12'h000; 
        10'b1011111011: data <= 12'hffd; 
        10'b1011111100: data <= 12'h001; 
        10'b1011111101: data <= 12'h001; 
        10'b1011111110: data <= 12'h000; 
        10'b1011111111: data <= 12'h001; 
        10'b1100000000: data <= 12'hfff; 
        10'b1100000001: data <= 12'hffe; 
        10'b1100000010: data <= 12'h001; 
        10'b1100000011: data <= 12'hffe; 
        10'b1100000100: data <= 12'hfff; 
        10'b1100000101: data <= 12'hffe; 
        10'b1100000110: data <= 12'h000; 
        10'b1100000111: data <= 12'hffe; 
        10'b1100001000: data <= 12'hffd; 
        10'b1100001001: data <= 12'hffd; 
        10'b1100001010: data <= 12'hffc; 
        10'b1100001011: data <= 12'hfff; 
        10'b1100001100: data <= 12'h001; 
        10'b1100001101: data <= 12'hffe; 
        10'b1100001110: data <= 12'hffd; 
        10'b1100001111: data <= 12'h001; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 7) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 13'h1ffc; 
        10'b0000000001: data <= 13'h0002; 
        10'b0000000010: data <= 13'h1fff; 
        10'b0000000011: data <= 13'h1fff; 
        10'b0000000100: data <= 13'h0003; 
        10'b0000000101: data <= 13'h0000; 
        10'b0000000110: data <= 13'h1ffd; 
        10'b0000000111: data <= 13'h1ffd; 
        10'b0000001000: data <= 13'h1fff; 
        10'b0000001001: data <= 13'h1fff; 
        10'b0000001010: data <= 13'h0003; 
        10'b0000001011: data <= 13'h0000; 
        10'b0000001100: data <= 13'h0001; 
        10'b0000001101: data <= 13'h1ffc; 
        10'b0000001110: data <= 13'h0000; 
        10'b0000001111: data <= 13'h1ffa; 
        10'b0000010000: data <= 13'h1ffb; 
        10'b0000010001: data <= 13'h1fff; 
        10'b0000010010: data <= 13'h1ffb; 
        10'b0000010011: data <= 13'h0003; 
        10'b0000010100: data <= 13'h1ffb; 
        10'b0000010101: data <= 13'h1fff; 
        10'b0000010110: data <= 13'h1ffb; 
        10'b0000010111: data <= 13'h1fff; 
        10'b0000011000: data <= 13'h0002; 
        10'b0000011001: data <= 13'h1fff; 
        10'b0000011010: data <= 13'h0000; 
        10'b0000011011: data <= 13'h0000; 
        10'b0000011100: data <= 13'h0002; 
        10'b0000011101: data <= 13'h0002; 
        10'b0000011110: data <= 13'h0001; 
        10'b0000011111: data <= 13'h1ffb; 
        10'b0000100000: data <= 13'h1ffb; 
        10'b0000100001: data <= 13'h0000; 
        10'b0000100010: data <= 13'h1ffc; 
        10'b0000100011: data <= 13'h1fff; 
        10'b0000100100: data <= 13'h1ffd; 
        10'b0000100101: data <= 13'h1ffa; 
        10'b0000100110: data <= 13'h1ffc; 
        10'b0000100111: data <= 13'h0000; 
        10'b0000101000: data <= 13'h0003; 
        10'b0000101001: data <= 13'h1ffb; 
        10'b0000101010: data <= 13'h1ffd; 
        10'b0000101011: data <= 13'h0002; 
        10'b0000101100: data <= 13'h1ffc; 
        10'b0000101101: data <= 13'h1ffb; 
        10'b0000101110: data <= 13'h0001; 
        10'b0000101111: data <= 13'h0002; 
        10'b0000110000: data <= 13'h1ffc; 
        10'b0000110001: data <= 13'h0001; 
        10'b0000110010: data <= 13'h1ffc; 
        10'b0000110011: data <= 13'h1ffc; 
        10'b0000110100: data <= 13'h1fff; 
        10'b0000110101: data <= 13'h0000; 
        10'b0000110110: data <= 13'h1fff; 
        10'b0000110111: data <= 13'h0003; 
        10'b0000111000: data <= 13'h1ffb; 
        10'b0000111001: data <= 13'h1ffd; 
        10'b0000111010: data <= 13'h1ffd; 
        10'b0000111011: data <= 13'h0001; 
        10'b0000111100: data <= 13'h0000; 
        10'b0000111101: data <= 13'h1ffb; 
        10'b0000111110: data <= 13'h1fff; 
        10'b0000111111: data <= 13'h0003; 
        10'b0001000000: data <= 13'h1ffe; 
        10'b0001000001: data <= 13'h1ffc; 
        10'b0001000010: data <= 13'h1ffc; 
        10'b0001000011: data <= 13'h1ffa; 
        10'b0001000100: data <= 13'h1ff9; 
        10'b0001000101: data <= 13'h1ffe; 
        10'b0001000110: data <= 13'h1ff9; 
        10'b0001000111: data <= 13'h1ff7; 
        10'b0001001000: data <= 13'h1ff9; 
        10'b0001001001: data <= 13'h1ffe; 
        10'b0001001010: data <= 13'h1ffa; 
        10'b0001001011: data <= 13'h1ff9; 
        10'b0001001100: data <= 13'h1fff; 
        10'b0001001101: data <= 13'h0002; 
        10'b0001001110: data <= 13'h0000; 
        10'b0001001111: data <= 13'h1ffc; 
        10'b0001010000: data <= 13'h0003; 
        10'b0001010001: data <= 13'h1ffa; 
        10'b0001010010: data <= 13'h1fff; 
        10'b0001010011: data <= 13'h0001; 
        10'b0001010100: data <= 13'h1ffb; 
        10'b0001010101: data <= 13'h1fff; 
        10'b0001010110: data <= 13'h0003; 
        10'b0001010111: data <= 13'h1ffb; 
        10'b0001011000: data <= 13'h1ffc; 
        10'b0001011001: data <= 13'h0002; 
        10'b0001011010: data <= 13'h0001; 
        10'b0001011011: data <= 13'h0000; 
        10'b0001011100: data <= 13'h0000; 
        10'b0001011101: data <= 13'h1fff; 
        10'b0001011110: data <= 13'h1ffe; 
        10'b0001011111: data <= 13'h1ff9; 
        10'b0001100000: data <= 13'h1ff6; 
        10'b0001100001: data <= 13'h1ffb; 
        10'b0001100010: data <= 13'h1ff8; 
        10'b0001100011: data <= 13'h1ff7; 
        10'b0001100100: data <= 13'h0001; 
        10'b0001100101: data <= 13'h0001; 
        10'b0001100110: data <= 13'h1ff6; 
        10'b0001100111: data <= 13'h1ff8; 
        10'b0001101000: data <= 13'h1ff4; 
        10'b0001101001: data <= 13'h1ff8; 
        10'b0001101010: data <= 13'h1ff6; 
        10'b0001101011: data <= 13'h1ff9; 
        10'b0001101100: data <= 13'h1ffb; 
        10'b0001101101: data <= 13'h0002; 
        10'b0001101110: data <= 13'h0002; 
        10'b0001101111: data <= 13'h1ffd; 
        10'b0001110000: data <= 13'h0001; 
        10'b0001110001: data <= 13'h1ffb; 
        10'b0001110010: data <= 13'h1ffc; 
        10'b0001110011: data <= 13'h1ffb; 
        10'b0001110100: data <= 13'h1ffa; 
        10'b0001110101: data <= 13'h1fff; 
        10'b0001110110: data <= 13'h1ffe; 
        10'b0001110111: data <= 13'h1ffb; 
        10'b0001111000: data <= 13'h1ffe; 
        10'b0001111001: data <= 13'h1fff; 
        10'b0001111010: data <= 13'h1ff7; 
        10'b0001111011: data <= 13'h1ff7; 
        10'b0001111100: data <= 13'h1ff8; 
        10'b0001111101: data <= 13'h1ff8; 
        10'b0001111110: data <= 13'h1ffe; 
        10'b0001111111: data <= 13'h1fff; 
        10'b0010000000: data <= 13'h1ff9; 
        10'b0010000001: data <= 13'h1ffa; 
        10'b0010000010: data <= 13'h1ffa; 
        10'b0010000011: data <= 13'h1ff7; 
        10'b0010000100: data <= 13'h1ffc; 
        10'b0010000101: data <= 13'h1ff4; 
        10'b0010000110: data <= 13'h1ffc; 
        10'b0010000111: data <= 13'h1fff; 
        10'b0010001000: data <= 13'h1ffb; 
        10'b0010001001: data <= 13'h1ffe; 
        10'b0010001010: data <= 13'h1ffd; 
        10'b0010001011: data <= 13'h0000; 
        10'b0010001100: data <= 13'h0001; 
        10'b0010001101: data <= 13'h1ffd; 
        10'b0010001110: data <= 13'h0000; 
        10'b0010001111: data <= 13'h1ffb; 
        10'b0010010000: data <= 13'h1fff; 
        10'b0010010001: data <= 13'h1ffe; 
        10'b0010010010: data <= 13'h1ffe; 
        10'b0010010011: data <= 13'h1ffc; 
        10'b0010010100: data <= 13'h1ffe; 
        10'b0010010101: data <= 13'h1ffa; 
        10'b0010010110: data <= 13'h1ffd; 
        10'b0010010111: data <= 13'h0002; 
        10'b0010011000: data <= 13'h0008; 
        10'b0010011001: data <= 13'h0010; 
        10'b0010011010: data <= 13'h0014; 
        10'b0010011011: data <= 13'h0014; 
        10'b0010011100: data <= 13'h0016; 
        10'b0010011101: data <= 13'h0018; 
        10'b0010011110: data <= 13'h0019; 
        10'b0010011111: data <= 13'h0009; 
        10'b0010100000: data <= 13'h0002; 
        10'b0010100001: data <= 13'h0004; 
        10'b0010100010: data <= 13'h1ffe; 
        10'b0010100011: data <= 13'h0000; 
        10'b0010100100: data <= 13'h1ff5; 
        10'b0010100101: data <= 13'h1ff8; 
        10'b0010100110: data <= 13'h1fff; 
        10'b0010100111: data <= 13'h1ffc; 
        10'b0010101000: data <= 13'h1ffe; 
        10'b0010101001: data <= 13'h1fff; 
        10'b0010101010: data <= 13'h0001; 
        10'b0010101011: data <= 13'h1ffe; 
        10'b0010101100: data <= 13'h0000; 
        10'b0010101101: data <= 13'h0000; 
        10'b0010101110: data <= 13'h0001; 
        10'b0010101111: data <= 13'h0000; 
        10'b0010110000: data <= 13'h1ffb; 
        10'b0010110001: data <= 13'h1ff7; 
        10'b0010110010: data <= 13'h0005; 
        10'b0010110011: data <= 13'h1fff; 
        10'b0010110100: data <= 13'h000e; 
        10'b0010110101: data <= 13'h000c; 
        10'b0010110110: data <= 13'h000b; 
        10'b0010110111: data <= 13'h0011; 
        10'b0010111000: data <= 13'h0015; 
        10'b0010111001: data <= 13'h001d; 
        10'b0010111010: data <= 13'h001b; 
        10'b0010111011: data <= 13'h0017; 
        10'b0010111100: data <= 13'h0016; 
        10'b0010111101: data <= 13'h001a; 
        10'b0010111110: data <= 13'h000f; 
        10'b0010111111: data <= 13'h0005; 
        10'b0011000000: data <= 13'h1ff5; 
        10'b0011000001: data <= 13'h1ff4; 
        10'b0011000010: data <= 13'h1ff8; 
        10'b0011000011: data <= 13'h0001; 
        10'b0011000100: data <= 13'h0003; 
        10'b0011000101: data <= 13'h0000; 
        10'b0011000110: data <= 13'h1fff; 
        10'b0011000111: data <= 13'h1ff9; 
        10'b0011001000: data <= 13'h1ff5; 
        10'b0011001001: data <= 13'h1fff; 
        10'b0011001010: data <= 13'h1ffc; 
        10'b0011001011: data <= 13'h0000; 
        10'b0011001100: data <= 13'h1ffb; 
        10'b0011001101: data <= 13'h1fff; 
        10'b0011001110: data <= 13'h0001; 
        10'b0011001111: data <= 13'h000a; 
        10'b0011010000: data <= 13'h0014; 
        10'b0011010001: data <= 13'h0013; 
        10'b0011010010: data <= 13'h0008; 
        10'b0011010011: data <= 13'h000c; 
        10'b0011010100: data <= 13'h0011; 
        10'b0011010101: data <= 13'h001f; 
        10'b0011010110: data <= 13'h0017; 
        10'b0011010111: data <= 13'h0014; 
        10'b0011011000: data <= 13'h0008; 
        10'b0011011001: data <= 13'h0010; 
        10'b0011011010: data <= 13'h0011; 
        10'b0011011011: data <= 13'h0009; 
        10'b0011011100: data <= 13'h1ff9; 
        10'b0011011101: data <= 13'h1ff5; 
        10'b0011011110: data <= 13'h1ff6; 
        10'b0011011111: data <= 13'h1fff; 
        10'b0011100000: data <= 13'h0003; 
        10'b0011100001: data <= 13'h0001; 
        10'b0011100010: data <= 13'h1fff; 
        10'b0011100011: data <= 13'h0000; 
        10'b0011100100: data <= 13'h1ff8; 
        10'b0011100101: data <= 13'h1ffa; 
        10'b0011100110: data <= 13'h1ffb; 
        10'b0011100111: data <= 13'h1ffa; 
        10'b0011101000: data <= 13'h1ffd; 
        10'b0011101001: data <= 13'h1ffd; 
        10'b0011101010: data <= 13'h000a; 
        10'b0011101011: data <= 13'h000a; 
        10'b0011101100: data <= 13'h0005; 
        10'b0011101101: data <= 13'h0002; 
        10'b0011101110: data <= 13'h0004; 
        10'b0011101111: data <= 13'h000e; 
        10'b0011110000: data <= 13'h0029; 
        10'b0011110001: data <= 13'h0021; 
        10'b0011110010: data <= 13'h001f; 
        10'b0011110011: data <= 13'h000a; 
        10'b0011110100: data <= 13'h0008; 
        10'b0011110101: data <= 13'h0007; 
        10'b0011110110: data <= 13'h0012; 
        10'b0011110111: data <= 13'h0020; 
        10'b0011111000: data <= 13'h1ffd; 
        10'b0011111001: data <= 13'h1ff6; 
        10'b0011111010: data <= 13'h1fff; 
        10'b0011111011: data <= 13'h1ffa; 
        10'b0011111100: data <= 13'h1fff; 
        10'b0011111101: data <= 13'h1fff; 
        10'b0011111110: data <= 13'h0001; 
        10'b0011111111: data <= 13'h0001; 
        10'b0100000000: data <= 13'h1ff6; 
        10'b0100000001: data <= 13'h1ff9; 
        10'b0100000010: data <= 13'h1ff6; 
        10'b0100000011: data <= 13'h1ffa; 
        10'b0100000100: data <= 13'h1ffa; 
        10'b0100000101: data <= 13'h1ffd; 
        10'b0100000110: data <= 13'h0007; 
        10'b0100000111: data <= 13'h1ffa; 
        10'b0100001000: data <= 13'h0003; 
        10'b0100001001: data <= 13'h000a; 
        10'b0100001010: data <= 13'h0009; 
        10'b0100001011: data <= 13'h0008; 
        10'b0100001100: data <= 13'h0017; 
        10'b0100001101: data <= 13'h001e; 
        10'b0100001110: data <= 13'h0023; 
        10'b0100001111: data <= 13'h0014; 
        10'b0100010000: data <= 13'h0006; 
        10'b0100010001: data <= 13'h1fff; 
        10'b0100010010: data <= 13'h000f; 
        10'b0100010011: data <= 13'h0020; 
        10'b0100010100: data <= 13'h0009; 
        10'b0100010101: data <= 13'h1ff8; 
        10'b0100010110: data <= 13'h0000; 
        10'b0100010111: data <= 13'h1fff; 
        10'b0100011000: data <= 13'h1ffb; 
        10'b0100011001: data <= 13'h0002; 
        10'b0100011010: data <= 13'h1ffc; 
        10'b0100011011: data <= 13'h1ff8; 
        10'b0100011100: data <= 13'h1ff9; 
        10'b0100011101: data <= 13'h1ffa; 
        10'b0100011110: data <= 13'h1ffb; 
        10'b0100011111: data <= 13'h0001; 
        10'b0100100000: data <= 13'h0003; 
        10'b0100100001: data <= 13'h1fff; 
        10'b0100100010: data <= 13'h1ffb; 
        10'b0100100011: data <= 13'h0002; 
        10'b0100100100: data <= 13'h0002; 
        10'b0100100101: data <= 13'h1fff; 
        10'b0100100110: data <= 13'h1ff5; 
        10'b0100100111: data <= 13'h1fed; 
        10'b0100101000: data <= 13'h1ff5; 
        10'b0100101001: data <= 13'h000b; 
        10'b0100101010: data <= 13'h001c; 
        10'b0100101011: data <= 13'h001d; 
        10'b0100101100: data <= 13'h0019; 
        10'b0100101101: data <= 13'h0012; 
        10'b0100101110: data <= 13'h001b; 
        10'b0100101111: data <= 13'h0025; 
        10'b0100110000: data <= 13'h0012; 
        10'b0100110001: data <= 13'h1ff9; 
        10'b0100110010: data <= 13'h1ff9; 
        10'b0100110011: data <= 13'h1ffa; 
        10'b0100110100: data <= 13'h1ffc; 
        10'b0100110101: data <= 13'h1ffb; 
        10'b0100110110: data <= 13'h0002; 
        10'b0100110111: data <= 13'h1ffe; 
        10'b0100111000: data <= 13'h1ff2; 
        10'b0100111001: data <= 13'h1ffd; 
        10'b0100111010: data <= 13'h0002; 
        10'b0100111011: data <= 13'h000b; 
        10'b0100111100: data <= 13'h0008; 
        10'b0100111101: data <= 13'h1ffd; 
        10'b0100111110: data <= 13'h0003; 
        10'b0100111111: data <= 13'h0000; 
        10'b0101000000: data <= 13'h0005; 
        10'b0101000001: data <= 13'h1ffc; 
        10'b0101000010: data <= 13'h1fe2; 
        10'b0101000011: data <= 13'h1fc9; 
        10'b0101000100: data <= 13'h1fcd; 
        10'b0101000101: data <= 13'h1fec; 
        10'b0101000110: data <= 13'h1ffd; 
        10'b0101000111: data <= 13'h000f; 
        10'b0101001000: data <= 13'h0017; 
        10'b0101001001: data <= 13'h0016; 
        10'b0101001010: data <= 13'h001d; 
        10'b0101001011: data <= 13'h0021; 
        10'b0101001100: data <= 13'h0018; 
        10'b0101001101: data <= 13'h1ffb; 
        10'b0101001110: data <= 13'h0000; 
        10'b0101001111: data <= 13'h1ffa; 
        10'b0101010000: data <= 13'h1ffc; 
        10'b0101010001: data <= 13'h1fff; 
        10'b0101010010: data <= 13'h1ffe; 
        10'b0101010011: data <= 13'h1ffe; 
        10'b0101010100: data <= 13'h1ff8; 
        10'b0101010101: data <= 13'h0001; 
        10'b0101010110: data <= 13'h000b; 
        10'b0101010111: data <= 13'h000c; 
        10'b0101011000: data <= 13'h0006; 
        10'b0101011001: data <= 13'h1ffe; 
        10'b0101011010: data <= 13'h0008; 
        10'b0101011011: data <= 13'h0006; 
        10'b0101011100: data <= 13'h000b; 
        10'b0101011101: data <= 13'h1ff7; 
        10'b0101011110: data <= 13'h1fc6; 
        10'b0101011111: data <= 13'h1fb8; 
        10'b0101100000: data <= 13'h1fb9; 
        10'b0101100001: data <= 13'h1fd9; 
        10'b0101100010: data <= 13'h1ff9; 
        10'b0101100011: data <= 13'h1ffd; 
        10'b0101100100: data <= 13'h0004; 
        10'b0101100101: data <= 13'h000a; 
        10'b0101100110: data <= 13'h0026; 
        10'b0101100111: data <= 13'h0023; 
        10'b0101101000: data <= 13'h0018; 
        10'b0101101001: data <= 13'h0001; 
        10'b0101101010: data <= 13'h1ffc; 
        10'b0101101011: data <= 13'h1ffc; 
        10'b0101101100: data <= 13'h1ffa; 
        10'b0101101101: data <= 13'h0000; 
        10'b0101101110: data <= 13'h0002; 
        10'b0101101111: data <= 13'h1ffb; 
        10'b0101110000: data <= 13'h1ffe; 
        10'b0101110001: data <= 13'h0007; 
        10'b0101110010: data <= 13'h000e; 
        10'b0101110011: data <= 13'h0012; 
        10'b0101110100: data <= 13'h000e; 
        10'b0101110101: data <= 13'h0009; 
        10'b0101110110: data <= 13'h000d; 
        10'b0101110111: data <= 13'h000a; 
        10'b0101111000: data <= 13'h0007; 
        10'b0101111001: data <= 13'h1fdd; 
        10'b0101111010: data <= 13'h1fc6; 
        10'b0101111011: data <= 13'h1fb6; 
        10'b0101111100: data <= 13'h1fc3; 
        10'b0101111101: data <= 13'h1fe2; 
        10'b0101111110: data <= 13'h1ff1; 
        10'b0101111111: data <= 13'h1fec; 
        10'b0110000000: data <= 13'h1ff1; 
        10'b0110000001: data <= 13'h0007; 
        10'b0110000010: data <= 13'h0019; 
        10'b0110000011: data <= 13'h0027; 
        10'b0110000100: data <= 13'h0016; 
        10'b0110000101: data <= 13'h0004; 
        10'b0110000110: data <= 13'h0000; 
        10'b0110000111: data <= 13'h0002; 
        10'b0110001000: data <= 13'h1fff; 
        10'b0110001001: data <= 13'h0002; 
        10'b0110001010: data <= 13'h1ffc; 
        10'b0110001011: data <= 13'h1ffd; 
        10'b0110001100: data <= 13'h1ff9; 
        10'b0110001101: data <= 13'h0012; 
        10'b0110001110: data <= 13'h0018; 
        10'b0110001111: data <= 13'h001d; 
        10'b0110010000: data <= 13'h000e; 
        10'b0110010001: data <= 13'h0011; 
        10'b0110010010: data <= 13'h0019; 
        10'b0110010011: data <= 13'h000e; 
        10'b0110010100: data <= 13'h0003; 
        10'b0110010101: data <= 13'h1fe1; 
        10'b0110010110: data <= 13'h1fbc; 
        10'b0110010111: data <= 13'h1fb6; 
        10'b0110011000: data <= 13'h1fc5; 
        10'b0110011001: data <= 13'h1fe0; 
        10'b0110011010: data <= 13'h1ff2; 
        10'b0110011011: data <= 13'h1fef; 
        10'b0110011100: data <= 13'h0002; 
        10'b0110011101: data <= 13'h000e; 
        10'b0110011110: data <= 13'h0011; 
        10'b0110011111: data <= 13'h0028; 
        10'b0110100000: data <= 13'h0015; 
        10'b0110100001: data <= 13'h1ffc; 
        10'b0110100010: data <= 13'h1ffe; 
        10'b0110100011: data <= 13'h1ffc; 
        10'b0110100100: data <= 13'h0002; 
        10'b0110100101: data <= 13'h0001; 
        10'b0110100110: data <= 13'h1ffc; 
        10'b0110100111: data <= 13'h1fff; 
        10'b0110101000: data <= 13'h0000; 
        10'b0110101001: data <= 13'h001a; 
        10'b0110101010: data <= 13'h0013; 
        10'b0110101011: data <= 13'h001a; 
        10'b0110101100: data <= 13'h0012; 
        10'b0110101101: data <= 13'h0018; 
        10'b0110101110: data <= 13'h001e; 
        10'b0110101111: data <= 13'h0008; 
        10'b0110110000: data <= 13'h1fe9; 
        10'b0110110001: data <= 13'h1fc7; 
        10'b0110110010: data <= 13'h1fb3; 
        10'b0110110011: data <= 13'h1fb7; 
        10'b0110110100: data <= 13'h1fcf; 
        10'b0110110101: data <= 13'h1fe8; 
        10'b0110110110: data <= 13'h1ff7; 
        10'b0110110111: data <= 13'h1ff7; 
        10'b0110111000: data <= 13'h0007; 
        10'b0110111001: data <= 13'h0007; 
        10'b0110111010: data <= 13'h0019; 
        10'b0110111011: data <= 13'h001e; 
        10'b0110111100: data <= 13'h000f; 
        10'b0110111101: data <= 13'h1ffe; 
        10'b0110111110: data <= 13'h0000; 
        10'b0110111111: data <= 13'h1ffc; 
        10'b0111000000: data <= 13'h0001; 
        10'b0111000001: data <= 13'h0003; 
        10'b0111000010: data <= 13'h1ffa; 
        10'b0111000011: data <= 13'h1ffd; 
        10'b0111000100: data <= 13'h0004; 
        10'b0111000101: data <= 13'h0017; 
        10'b0111000110: data <= 13'h001d; 
        10'b0111000111: data <= 13'h0017; 
        10'b0111001000: data <= 13'h0010; 
        10'b0111001001: data <= 13'h0010; 
        10'b0111001010: data <= 13'h001b; 
        10'b0111001011: data <= 13'h1ffc; 
        10'b0111001100: data <= 13'h1fd4; 
        10'b0111001101: data <= 13'h1fb4; 
        10'b0111001110: data <= 13'h1fb6; 
        10'b0111001111: data <= 13'h1fc5; 
        10'b0111010000: data <= 13'h1fe0; 
        10'b0111010001: data <= 13'h1ff1; 
        10'b0111010010: data <= 13'h0000; 
        10'b0111010011: data <= 13'h0005; 
        10'b0111010100: data <= 13'h000b; 
        10'b0111010101: data <= 13'h0010; 
        10'b0111010110: data <= 13'h0017; 
        10'b0111010111: data <= 13'h0016; 
        10'b0111011000: data <= 13'h0008; 
        10'b0111011001: data <= 13'h0000; 
        10'b0111011010: data <= 13'h1ffd; 
        10'b0111011011: data <= 13'h1ffc; 
        10'b0111011100: data <= 13'h1ffe; 
        10'b0111011101: data <= 13'h0001; 
        10'b0111011110: data <= 13'h1ffb; 
        10'b0111011111: data <= 13'h1ff6; 
        10'b0111100000: data <= 13'h0001; 
        10'b0111100001: data <= 13'h0011; 
        10'b0111100010: data <= 13'h0015; 
        10'b0111100011: data <= 13'h0014; 
        10'b0111100100: data <= 13'h0006; 
        10'b0111100101: data <= 13'h0010; 
        10'b0111100110: data <= 13'h001a; 
        10'b0111100111: data <= 13'h1ffc; 
        10'b0111101000: data <= 13'h1fcc; 
        10'b0111101001: data <= 13'h1fb5; 
        10'b0111101010: data <= 13'h1fbe; 
        10'b0111101011: data <= 13'h1fd9; 
        10'b0111101100: data <= 13'h1ffb; 
        10'b0111101101: data <= 13'h000a; 
        10'b0111101110: data <= 13'h000e; 
        10'b0111101111: data <= 13'h000d; 
        10'b0111110000: data <= 13'h0011; 
        10'b0111110001: data <= 13'h000d; 
        10'b0111110010: data <= 13'h000a; 
        10'b0111110011: data <= 13'h000c; 
        10'b0111110100: data <= 13'h1fff; 
        10'b0111110101: data <= 13'h1ffe; 
        10'b0111110110: data <= 13'h0001; 
        10'b0111110111: data <= 13'h1ffc; 
        10'b0111111000: data <= 13'h1ffd; 
        10'b0111111001: data <= 13'h0001; 
        10'b0111111010: data <= 13'h1ffe; 
        10'b0111111011: data <= 13'h1ffc; 
        10'b0111111100: data <= 13'h1ffe; 
        10'b0111111101: data <= 13'h000b; 
        10'b0111111110: data <= 13'h0016; 
        10'b0111111111: data <= 13'h000d; 
        10'b1000000000: data <= 13'h0008; 
        10'b1000000001: data <= 13'h0016; 
        10'b1000000010: data <= 13'h0029; 
        10'b1000000011: data <= 13'h0002; 
        10'b1000000100: data <= 13'h1fdf; 
        10'b1000000101: data <= 13'h1fca; 
        10'b1000000110: data <= 13'h1fda; 
        10'b1000000111: data <= 13'h1ff5; 
        10'b1000001000: data <= 13'h000c; 
        10'b1000001001: data <= 13'h000d; 
        10'b1000001010: data <= 13'h000e; 
        10'b1000001011: data <= 13'h0007; 
        10'b1000001100: data <= 13'h0004; 
        10'b1000001101: data <= 13'h0006; 
        10'b1000001110: data <= 13'h000b; 
        10'b1000001111: data <= 13'h0007; 
        10'b1000010000: data <= 13'h1fff; 
        10'b1000010001: data <= 13'h1ffd; 
        10'b1000010010: data <= 13'h0000; 
        10'b1000010011: data <= 13'h1ffe; 
        10'b1000010100: data <= 13'h1ffe; 
        10'b1000010101: data <= 13'h1ffe; 
        10'b1000010110: data <= 13'h1ffe; 
        10'b1000010111: data <= 13'h1ff7; 
        10'b1000011000: data <= 13'h0004; 
        10'b1000011001: data <= 13'h000c; 
        10'b1000011010: data <= 13'h001c; 
        10'b1000011011: data <= 13'h0019; 
        10'b1000011100: data <= 13'h0014; 
        10'b1000011101: data <= 13'h001a; 
        10'b1000011110: data <= 13'h0029; 
        10'b1000011111: data <= 13'h001d; 
        10'b1000100000: data <= 13'h0006; 
        10'b1000100001: data <= 13'h1ff3; 
        10'b1000100010: data <= 13'h1ffa; 
        10'b1000100011: data <= 13'h1ffc; 
        10'b1000100100: data <= 13'h0006; 
        10'b1000100101: data <= 13'h1ffd; 
        10'b1000100110: data <= 13'h1ffb; 
        10'b1000100111: data <= 13'h1ffd; 
        10'b1000101000: data <= 13'h0007; 
        10'b1000101001: data <= 13'h0006; 
        10'b1000101010: data <= 13'h000c; 
        10'b1000101011: data <= 13'h1ffe; 
        10'b1000101100: data <= 13'h0002; 
        10'b1000101101: data <= 13'h1ffd; 
        10'b1000101110: data <= 13'h1ffa; 
        10'b1000101111: data <= 13'h0002; 
        10'b1000110000: data <= 13'h0002; 
        10'b1000110001: data <= 13'h0003; 
        10'b1000110010: data <= 13'h1ffe; 
        10'b1000110011: data <= 13'h1ffc; 
        10'b1000110100: data <= 13'h1ffd; 
        10'b1000110101: data <= 13'h000c; 
        10'b1000110110: data <= 13'h0016; 
        10'b1000110111: data <= 13'h0011; 
        10'b1000111000: data <= 13'h0014; 
        10'b1000111001: data <= 13'h0019; 
        10'b1000111010: data <= 13'h0027; 
        10'b1000111011: data <= 13'h0027; 
        10'b1000111100: data <= 13'h0014; 
        10'b1000111101: data <= 13'h0006; 
        10'b1000111110: data <= 13'h1ffc; 
        10'b1000111111: data <= 13'h0003; 
        10'b1001000000: data <= 13'h0003; 
        10'b1001000001: data <= 13'h1ffa; 
        10'b1001000010: data <= 13'h1ffc; 
        10'b1001000011: data <= 13'h1ffa; 
        10'b1001000100: data <= 13'h0003; 
        10'b1001000101: data <= 13'h0004; 
        10'b1001000110: data <= 13'h0006; 
        10'b1001000111: data <= 13'h0002; 
        10'b1001001000: data <= 13'h1ffd; 
        10'b1001001001: data <= 13'h1fff; 
        10'b1001001010: data <= 13'h1ffb; 
        10'b1001001011: data <= 13'h1ffd; 
        10'b1001001100: data <= 13'h1ffc; 
        10'b1001001101: data <= 13'h1ffb; 
        10'b1001001110: data <= 13'h1ffe; 
        10'b1001001111: data <= 13'h1ffc; 
        10'b1001010000: data <= 13'h1ffe; 
        10'b1001010001: data <= 13'h0003; 
        10'b1001010010: data <= 13'h000e; 
        10'b1001010011: data <= 13'h0017; 
        10'b1001010100: data <= 13'h0010; 
        10'b1001010101: data <= 13'h0011; 
        10'b1001010110: data <= 13'h0022; 
        10'b1001010111: data <= 13'h0026; 
        10'b1001011000: data <= 13'h0019; 
        10'b1001011001: data <= 13'h000a; 
        10'b1001011010: data <= 13'h0004; 
        10'b1001011011: data <= 13'h0001; 
        10'b1001011100: data <= 13'h1fff; 
        10'b1001011101: data <= 13'h1ff6; 
        10'b1001011110: data <= 13'h1ff8; 
        10'b1001011111: data <= 13'h1ffb; 
        10'b1001100000: data <= 13'h0004; 
        10'b1001100001: data <= 13'h0000; 
        10'b1001100010: data <= 13'h1ffb; 
        10'b1001100011: data <= 13'h1ff8; 
        10'b1001100100: data <= 13'h1ffe; 
        10'b1001100101: data <= 13'h1ffe; 
        10'b1001100110: data <= 13'h1ffc; 
        10'b1001100111: data <= 13'h1ffd; 
        10'b1001101000: data <= 13'h1ffc; 
        10'b1001101001: data <= 13'h0000; 
        10'b1001101010: data <= 13'h0000; 
        10'b1001101011: data <= 13'h1ffd; 
        10'b1001101100: data <= 13'h1ffb; 
        10'b1001101101: data <= 13'h0002; 
        10'b1001101110: data <= 13'h000a; 
        10'b1001101111: data <= 13'h0009; 
        10'b1001110000: data <= 13'h0019; 
        10'b1001110001: data <= 13'h0015; 
        10'b1001110010: data <= 13'h0017; 
        10'b1001110011: data <= 13'h001b; 
        10'b1001110100: data <= 13'h0017; 
        10'b1001110101: data <= 13'h001e; 
        10'b1001110110: data <= 13'h000d; 
        10'b1001110111: data <= 13'h000d; 
        10'b1001111000: data <= 13'h0007; 
        10'b1001111001: data <= 13'h1ffa; 
        10'b1001111010: data <= 13'h1ffb; 
        10'b1001111011: data <= 13'h0000; 
        10'b1001111100: data <= 13'h1ff9; 
        10'b1001111101: data <= 13'h1ff9; 
        10'b1001111110: data <= 13'h1ffd; 
        10'b1001111111: data <= 13'h1ffc; 
        10'b1010000000: data <= 13'h1fff; 
        10'b1010000001: data <= 13'h1ffe; 
        10'b1010000010: data <= 13'h1ffd; 
        10'b1010000011: data <= 13'h1ffe; 
        10'b1010000100: data <= 13'h1ffc; 
        10'b1010000101: data <= 13'h1fff; 
        10'b1010000110: data <= 13'h0000; 
        10'b1010000111: data <= 13'h1ffb; 
        10'b1010001000: data <= 13'h1ffa; 
        10'b1010001001: data <= 13'h1ffe; 
        10'b1010001010: data <= 13'h1fff; 
        10'b1010001011: data <= 13'h0007; 
        10'b1010001100: data <= 13'h000a; 
        10'b1010001101: data <= 13'h0017; 
        10'b1010001110: data <= 13'h001c; 
        10'b1010001111: data <= 13'h0022; 
        10'b1010010000: data <= 13'h0022; 
        10'b1010010001: data <= 13'h0014; 
        10'b1010010010: data <= 13'h0011; 
        10'b1010010011: data <= 13'h0009; 
        10'b1010010100: data <= 13'h0004; 
        10'b1010010101: data <= 13'h0000; 
        10'b1010010110: data <= 13'h1ff3; 
        10'b1010010111: data <= 13'h1ff0; 
        10'b1010011000: data <= 13'h1ff3; 
        10'b1010011001: data <= 13'h1ffa; 
        10'b1010011010: data <= 13'h1ffb; 
        10'b1010011011: data <= 13'h1fff; 
        10'b1010011100: data <= 13'h1ffe; 
        10'b1010011101: data <= 13'h0002; 
        10'b1010011110: data <= 13'h1ffd; 
        10'b1010011111: data <= 13'h1ffa; 
        10'b1010100000: data <= 13'h1ffd; 
        10'b1010100001: data <= 13'h1fff; 
        10'b1010100010: data <= 13'h1ffa; 
        10'b1010100011: data <= 13'h0000; 
        10'b1010100100: data <= 13'h1ffe; 
        10'b1010100101: data <= 13'h1fff; 
        10'b1010100110: data <= 13'h1ff9; 
        10'b1010100111: data <= 13'h1ff7; 
        10'b1010101000: data <= 13'h1ffb; 
        10'b1010101001: data <= 13'h1ffc; 
        10'b1010101010: data <= 13'h0005; 
        10'b1010101011: data <= 13'h0004; 
        10'b1010101100: data <= 13'h0009; 
        10'b1010101101: data <= 13'h000e; 
        10'b1010101110: data <= 13'h0007; 
        10'b1010101111: data <= 13'h1ffa; 
        10'b1010110000: data <= 13'h1ff7; 
        10'b1010110001: data <= 13'h1ff6; 
        10'b1010110010: data <= 13'h1ff7; 
        10'b1010110011: data <= 13'h1ff4; 
        10'b1010110100: data <= 13'h1ff4; 
        10'b1010110101: data <= 13'h1ff5; 
        10'b1010110110: data <= 13'h1ffe; 
        10'b1010110111: data <= 13'h1ffd; 
        10'b1010111000: data <= 13'h1ffb; 
        10'b1010111001: data <= 13'h1ffd; 
        10'b1010111010: data <= 13'h0000; 
        10'b1010111011: data <= 13'h1ffc; 
        10'b1010111100: data <= 13'h1ffd; 
        10'b1010111101: data <= 13'h0003; 
        10'b1010111110: data <= 13'h1ffe; 
        10'b1010111111: data <= 13'h0003; 
        10'b1011000000: data <= 13'h0003; 
        10'b1011000001: data <= 13'h0000; 
        10'b1011000010: data <= 13'h1ffa; 
        10'b1011000011: data <= 13'h1ffd; 
        10'b1011000100: data <= 13'h1ff4; 
        10'b1011000101: data <= 13'h1ff5; 
        10'b1011000110: data <= 13'h1ff2; 
        10'b1011000111: data <= 13'h1fee; 
        10'b1011001000: data <= 13'h1fec; 
        10'b1011001001: data <= 13'h1fed; 
        10'b1011001010: data <= 13'h1fea; 
        10'b1011001011: data <= 13'h1fec; 
        10'b1011001100: data <= 13'h1fed; 
        10'b1011001101: data <= 13'h1ff5; 
        10'b1011001110: data <= 13'h1ff7; 
        10'b1011001111: data <= 13'h1ff8; 
        10'b1011010000: data <= 13'h1ff7; 
        10'b1011010001: data <= 13'h1ff8; 
        10'b1011010010: data <= 13'h1ffd; 
        10'b1011010011: data <= 13'h0003; 
        10'b1011010100: data <= 13'h0001; 
        10'b1011010101: data <= 13'h1ffe; 
        10'b1011010110: data <= 13'h1ffd; 
        10'b1011010111: data <= 13'h1fff; 
        10'b1011011000: data <= 13'h0003; 
        10'b1011011001: data <= 13'h0002; 
        10'b1011011010: data <= 13'h1ffe; 
        10'b1011011011: data <= 13'h0000; 
        10'b1011011100: data <= 13'h1ffd; 
        10'b1011011101: data <= 13'h1ffd; 
        10'b1011011110: data <= 13'h1ffb; 
        10'b1011011111: data <= 13'h0001; 
        10'b1011100000: data <= 13'h1ffd; 
        10'b1011100001: data <= 13'h1ff6; 
        10'b1011100010: data <= 13'h1ff6; 
        10'b1011100011: data <= 13'h1ff7; 
        10'b1011100100: data <= 13'h1ffc; 
        10'b1011100101: data <= 13'h1ff7; 
        10'b1011100110: data <= 13'h1ff8; 
        10'b1011100111: data <= 13'h1ffd; 
        10'b1011101000: data <= 13'h1ff7; 
        10'b1011101001: data <= 13'h1ff9; 
        10'b1011101010: data <= 13'h1ffb; 
        10'b1011101011: data <= 13'h1ff9; 
        10'b1011101100: data <= 13'h1ffd; 
        10'b1011101101: data <= 13'h1ff8; 
        10'b1011101110: data <= 13'h1ff9; 
        10'b1011101111: data <= 13'h0003; 
        10'b1011110000: data <= 13'h1ffc; 
        10'b1011110001: data <= 13'h0001; 
        10'b1011110010: data <= 13'h0002; 
        10'b1011110011: data <= 13'h1fff; 
        10'b1011110100: data <= 13'h1ffb; 
        10'b1011110101: data <= 13'h0002; 
        10'b1011110110: data <= 13'h1fff; 
        10'b1011110111: data <= 13'h1ffd; 
        10'b1011111000: data <= 13'h0002; 
        10'b1011111001: data <= 13'h0000; 
        10'b1011111010: data <= 13'h0001; 
        10'b1011111011: data <= 13'h1ffa; 
        10'b1011111100: data <= 13'h0003; 
        10'b1011111101: data <= 13'h0003; 
        10'b1011111110: data <= 13'h0001; 
        10'b1011111111: data <= 13'h0002; 
        10'b1100000000: data <= 13'h1fff; 
        10'b1100000001: data <= 13'h1ffd; 
        10'b1100000010: data <= 13'h0002; 
        10'b1100000011: data <= 13'h1ffb; 
        10'b1100000100: data <= 13'h1ffe; 
        10'b1100000101: data <= 13'h1ffd; 
        10'b1100000110: data <= 13'h1fff; 
        10'b1100000111: data <= 13'h1ffd; 
        10'b1100001000: data <= 13'h1ffa; 
        10'b1100001001: data <= 13'h1ffb; 
        10'b1100001010: data <= 13'h1ff9; 
        10'b1100001011: data <= 13'h1ffe; 
        10'b1100001100: data <= 13'h0001; 
        10'b1100001101: data <= 13'h1ffb; 
        10'b1100001110: data <= 13'h1ffa; 
        10'b1100001111: data <= 13'h0002; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 8) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 14'h3ff8; 
        10'b0000000001: data <= 14'h0005; 
        10'b0000000010: data <= 14'h3ffd; 
        10'b0000000011: data <= 14'h3fff; 
        10'b0000000100: data <= 14'h0006; 
        10'b0000000101: data <= 14'h3fff; 
        10'b0000000110: data <= 14'h3ffb; 
        10'b0000000111: data <= 14'h3ffa; 
        10'b0000001000: data <= 14'h3fff; 
        10'b0000001001: data <= 14'h3ffd; 
        10'b0000001010: data <= 14'h0006; 
        10'b0000001011: data <= 14'h0000; 
        10'b0000001100: data <= 14'h0003; 
        10'b0000001101: data <= 14'h3ff8; 
        10'b0000001110: data <= 14'h0000; 
        10'b0000001111: data <= 14'h3ff5; 
        10'b0000010000: data <= 14'h3ff7; 
        10'b0000010001: data <= 14'h3ffe; 
        10'b0000010010: data <= 14'h3ff7; 
        10'b0000010011: data <= 14'h0006; 
        10'b0000010100: data <= 14'h3ff7; 
        10'b0000010101: data <= 14'h3ffd; 
        10'b0000010110: data <= 14'h3ff6; 
        10'b0000010111: data <= 14'h3fff; 
        10'b0000011000: data <= 14'h0003; 
        10'b0000011001: data <= 14'h3ffe; 
        10'b0000011010: data <= 14'h0000; 
        10'b0000011011: data <= 14'h0000; 
        10'b0000011100: data <= 14'h0004; 
        10'b0000011101: data <= 14'h0004; 
        10'b0000011110: data <= 14'h0001; 
        10'b0000011111: data <= 14'h3ff6; 
        10'b0000100000: data <= 14'h3ff6; 
        10'b0000100001: data <= 14'h0001; 
        10'b0000100010: data <= 14'h3ff8; 
        10'b0000100011: data <= 14'h3ffe; 
        10'b0000100100: data <= 14'h3ffa; 
        10'b0000100101: data <= 14'h3ff5; 
        10'b0000100110: data <= 14'h3ff9; 
        10'b0000100111: data <= 14'h0001; 
        10'b0000101000: data <= 14'h0007; 
        10'b0000101001: data <= 14'h3ff6; 
        10'b0000101010: data <= 14'h3ffb; 
        10'b0000101011: data <= 14'h0003; 
        10'b0000101100: data <= 14'h3ff8; 
        10'b0000101101: data <= 14'h3ff5; 
        10'b0000101110: data <= 14'h0002; 
        10'b0000101111: data <= 14'h0005; 
        10'b0000110000: data <= 14'h3ff8; 
        10'b0000110001: data <= 14'h0002; 
        10'b0000110010: data <= 14'h3ff9; 
        10'b0000110011: data <= 14'h3ff7; 
        10'b0000110100: data <= 14'h3ffe; 
        10'b0000110101: data <= 14'h0001; 
        10'b0000110110: data <= 14'h3ffd; 
        10'b0000110111: data <= 14'h0006; 
        10'b0000111000: data <= 14'h3ff6; 
        10'b0000111001: data <= 14'h3ffa; 
        10'b0000111010: data <= 14'h3ff9; 
        10'b0000111011: data <= 14'h0003; 
        10'b0000111100: data <= 14'h0001; 
        10'b0000111101: data <= 14'h3ff5; 
        10'b0000111110: data <= 14'h3ffd; 
        10'b0000111111: data <= 14'h0006; 
        10'b0001000000: data <= 14'h3ffd; 
        10'b0001000001: data <= 14'h3ff8; 
        10'b0001000010: data <= 14'h3ff9; 
        10'b0001000011: data <= 14'h3ff3; 
        10'b0001000100: data <= 14'h3ff3; 
        10'b0001000101: data <= 14'h3ffb; 
        10'b0001000110: data <= 14'h3ff2; 
        10'b0001000111: data <= 14'h3fee; 
        10'b0001001000: data <= 14'h3ff3; 
        10'b0001001001: data <= 14'h3ffd; 
        10'b0001001010: data <= 14'h3ff5; 
        10'b0001001011: data <= 14'h3ff2; 
        10'b0001001100: data <= 14'h3ffe; 
        10'b0001001101: data <= 14'h0004; 
        10'b0001001110: data <= 14'h0001; 
        10'b0001001111: data <= 14'h3ff8; 
        10'b0001010000: data <= 14'h0005; 
        10'b0001010001: data <= 14'h3ff5; 
        10'b0001010010: data <= 14'h3ffd; 
        10'b0001010011: data <= 14'h0003; 
        10'b0001010100: data <= 14'h3ff5; 
        10'b0001010101: data <= 14'h3ffd; 
        10'b0001010110: data <= 14'h0006; 
        10'b0001010111: data <= 14'h3ff6; 
        10'b0001011000: data <= 14'h3ff9; 
        10'b0001011001: data <= 14'h0005; 
        10'b0001011010: data <= 14'h0002; 
        10'b0001011011: data <= 14'h0000; 
        10'b0001011100: data <= 14'h0001; 
        10'b0001011101: data <= 14'h3ffd; 
        10'b0001011110: data <= 14'h3ffc; 
        10'b0001011111: data <= 14'h3ff2; 
        10'b0001100000: data <= 14'h3fed; 
        10'b0001100001: data <= 14'h3ff5; 
        10'b0001100010: data <= 14'h3ff1; 
        10'b0001100011: data <= 14'h3fef; 
        10'b0001100100: data <= 14'h0003; 
        10'b0001100101: data <= 14'h0001; 
        10'b0001100110: data <= 14'h3fed; 
        10'b0001100111: data <= 14'h3ff0; 
        10'b0001101000: data <= 14'h3fe9; 
        10'b0001101001: data <= 14'h3fef; 
        10'b0001101010: data <= 14'h3fec; 
        10'b0001101011: data <= 14'h3ff2; 
        10'b0001101100: data <= 14'h3ff6; 
        10'b0001101101: data <= 14'h0004; 
        10'b0001101110: data <= 14'h0004; 
        10'b0001101111: data <= 14'h3ffa; 
        10'b0001110000: data <= 14'h0001; 
        10'b0001110001: data <= 14'h3ff5; 
        10'b0001110010: data <= 14'h3ff8; 
        10'b0001110011: data <= 14'h3ff5; 
        10'b0001110100: data <= 14'h3ff4; 
        10'b0001110101: data <= 14'h3ffe; 
        10'b0001110110: data <= 14'h3ffd; 
        10'b0001110111: data <= 14'h3ff5; 
        10'b0001111000: data <= 14'h3ffc; 
        10'b0001111001: data <= 14'h3ffe; 
        10'b0001111010: data <= 14'h3fef; 
        10'b0001111011: data <= 14'h3fef; 
        10'b0001111100: data <= 14'h3fef; 
        10'b0001111101: data <= 14'h3ff0; 
        10'b0001111110: data <= 14'h3ffc; 
        10'b0001111111: data <= 14'h3ffe; 
        10'b0010000000: data <= 14'h3ff3; 
        10'b0010000001: data <= 14'h3ff4; 
        10'b0010000010: data <= 14'h3ff3; 
        10'b0010000011: data <= 14'h3fee; 
        10'b0010000100: data <= 14'h3ff9; 
        10'b0010000101: data <= 14'h3fe9; 
        10'b0010000110: data <= 14'h3ff7; 
        10'b0010000111: data <= 14'h3fff; 
        10'b0010001000: data <= 14'h3ff6; 
        10'b0010001001: data <= 14'h3ffb; 
        10'b0010001010: data <= 14'h3ffa; 
        10'b0010001011: data <= 14'h3fff; 
        10'b0010001100: data <= 14'h0003; 
        10'b0010001101: data <= 14'h3ffb; 
        10'b0010001110: data <= 14'h0000; 
        10'b0010001111: data <= 14'h3ff7; 
        10'b0010010000: data <= 14'h3ffd; 
        10'b0010010001: data <= 14'h3ffb; 
        10'b0010010010: data <= 14'h3ffd; 
        10'b0010010011: data <= 14'h3ff9; 
        10'b0010010100: data <= 14'h3ffd; 
        10'b0010010101: data <= 14'h3ff3; 
        10'b0010010110: data <= 14'h3ffa; 
        10'b0010010111: data <= 14'h0004; 
        10'b0010011000: data <= 14'h000f; 
        10'b0010011001: data <= 14'h0021; 
        10'b0010011010: data <= 14'h0027; 
        10'b0010011011: data <= 14'h0027; 
        10'b0010011100: data <= 14'h002c; 
        10'b0010011101: data <= 14'h002f; 
        10'b0010011110: data <= 14'h0032; 
        10'b0010011111: data <= 14'h0012; 
        10'b0010100000: data <= 14'h0003; 
        10'b0010100001: data <= 14'h0008; 
        10'b0010100010: data <= 14'h3ffc; 
        10'b0010100011: data <= 14'h3fff; 
        10'b0010100100: data <= 14'h3feb; 
        10'b0010100101: data <= 14'h3ff1; 
        10'b0010100110: data <= 14'h3fff; 
        10'b0010100111: data <= 14'h3ff8; 
        10'b0010101000: data <= 14'h3ffc; 
        10'b0010101001: data <= 14'h3ffe; 
        10'b0010101010: data <= 14'h0001; 
        10'b0010101011: data <= 14'h3ffc; 
        10'b0010101100: data <= 14'h0000; 
        10'b0010101101: data <= 14'h0001; 
        10'b0010101110: data <= 14'h0001; 
        10'b0010101111: data <= 14'h0000; 
        10'b0010110000: data <= 14'h3ff5; 
        10'b0010110001: data <= 14'h3fee; 
        10'b0010110010: data <= 14'h000a; 
        10'b0010110011: data <= 14'h3ffe; 
        10'b0010110100: data <= 14'h001b; 
        10'b0010110101: data <= 14'h0018; 
        10'b0010110110: data <= 14'h0017; 
        10'b0010110111: data <= 14'h0022; 
        10'b0010111000: data <= 14'h0029; 
        10'b0010111001: data <= 14'h003b; 
        10'b0010111010: data <= 14'h0037; 
        10'b0010111011: data <= 14'h002f; 
        10'b0010111100: data <= 14'h002d; 
        10'b0010111101: data <= 14'h0033; 
        10'b0010111110: data <= 14'h001d; 
        10'b0010111111: data <= 14'h000a; 
        10'b0011000000: data <= 14'h3fea; 
        10'b0011000001: data <= 14'h3fe9; 
        10'b0011000010: data <= 14'h3ff0; 
        10'b0011000011: data <= 14'h0002; 
        10'b0011000100: data <= 14'h0005; 
        10'b0011000101: data <= 14'h0001; 
        10'b0011000110: data <= 14'h3fff; 
        10'b0011000111: data <= 14'h3ff2; 
        10'b0011001000: data <= 14'h3feb; 
        10'b0011001001: data <= 14'h3ffe; 
        10'b0011001010: data <= 14'h3ff7; 
        10'b0011001011: data <= 14'h0000; 
        10'b0011001100: data <= 14'h3ff6; 
        10'b0011001101: data <= 14'h3ffd; 
        10'b0011001110: data <= 14'h0002; 
        10'b0011001111: data <= 14'h0013; 
        10'b0011010000: data <= 14'h0028; 
        10'b0011010001: data <= 14'h0025; 
        10'b0011010010: data <= 14'h000f; 
        10'b0011010011: data <= 14'h0018; 
        10'b0011010100: data <= 14'h0022; 
        10'b0011010101: data <= 14'h003f; 
        10'b0011010110: data <= 14'h002e; 
        10'b0011010111: data <= 14'h0029; 
        10'b0011011000: data <= 14'h0011; 
        10'b0011011001: data <= 14'h0020; 
        10'b0011011010: data <= 14'h0023; 
        10'b0011011011: data <= 14'h0012; 
        10'b0011011100: data <= 14'h3ff2; 
        10'b0011011101: data <= 14'h3fea; 
        10'b0011011110: data <= 14'h3fec; 
        10'b0011011111: data <= 14'h3fff; 
        10'b0011100000: data <= 14'h0006; 
        10'b0011100001: data <= 14'h0002; 
        10'b0011100010: data <= 14'h3ffd; 
        10'b0011100011: data <= 14'h0000; 
        10'b0011100100: data <= 14'h3ff0; 
        10'b0011100101: data <= 14'h3ff4; 
        10'b0011100110: data <= 14'h3ff6; 
        10'b0011100111: data <= 14'h3ff4; 
        10'b0011101000: data <= 14'h3ffa; 
        10'b0011101001: data <= 14'h3ff9; 
        10'b0011101010: data <= 14'h0013; 
        10'b0011101011: data <= 14'h0014; 
        10'b0011101100: data <= 14'h000a; 
        10'b0011101101: data <= 14'h0004; 
        10'b0011101110: data <= 14'h0007; 
        10'b0011101111: data <= 14'h001c; 
        10'b0011110000: data <= 14'h0053; 
        10'b0011110001: data <= 14'h0042; 
        10'b0011110010: data <= 14'h003d; 
        10'b0011110011: data <= 14'h0013; 
        10'b0011110100: data <= 14'h0010; 
        10'b0011110101: data <= 14'h000f; 
        10'b0011110110: data <= 14'h0024; 
        10'b0011110111: data <= 14'h003f; 
        10'b0011111000: data <= 14'h3ff9; 
        10'b0011111001: data <= 14'h3feb; 
        10'b0011111010: data <= 14'h3ffe; 
        10'b0011111011: data <= 14'h3ff5; 
        10'b0011111100: data <= 14'h3ffe; 
        10'b0011111101: data <= 14'h3fff; 
        10'b0011111110: data <= 14'h0002; 
        10'b0011111111: data <= 14'h0001; 
        10'b0100000000: data <= 14'h3fed; 
        10'b0100000001: data <= 14'h3ff2; 
        10'b0100000010: data <= 14'h3fec; 
        10'b0100000011: data <= 14'h3ff5; 
        10'b0100000100: data <= 14'h3ff5; 
        10'b0100000101: data <= 14'h3ffa; 
        10'b0100000110: data <= 14'h000e; 
        10'b0100000111: data <= 14'h3ff4; 
        10'b0100001000: data <= 14'h0007; 
        10'b0100001001: data <= 14'h0015; 
        10'b0100001010: data <= 14'h0012; 
        10'b0100001011: data <= 14'h0010; 
        10'b0100001100: data <= 14'h002d; 
        10'b0100001101: data <= 14'h003c; 
        10'b0100001110: data <= 14'h0045; 
        10'b0100001111: data <= 14'h0028; 
        10'b0100010000: data <= 14'h000c; 
        10'b0100010001: data <= 14'h3ffe; 
        10'b0100010010: data <= 14'h001e; 
        10'b0100010011: data <= 14'h0040; 
        10'b0100010100: data <= 14'h0013; 
        10'b0100010101: data <= 14'h3ff0; 
        10'b0100010110: data <= 14'h0000; 
        10'b0100010111: data <= 14'h3ffe; 
        10'b0100011000: data <= 14'h3ff6; 
        10'b0100011001: data <= 14'h0005; 
        10'b0100011010: data <= 14'h3ff7; 
        10'b0100011011: data <= 14'h3ff0; 
        10'b0100011100: data <= 14'h3ff2; 
        10'b0100011101: data <= 14'h3ff5; 
        10'b0100011110: data <= 14'h3ff6; 
        10'b0100011111: data <= 14'h0001; 
        10'b0100100000: data <= 14'h0007; 
        10'b0100100001: data <= 14'h3ffe; 
        10'b0100100010: data <= 14'h3ff5; 
        10'b0100100011: data <= 14'h0004; 
        10'b0100100100: data <= 14'h0004; 
        10'b0100100101: data <= 14'h3ffd; 
        10'b0100100110: data <= 14'h3fea; 
        10'b0100100111: data <= 14'h3fdb; 
        10'b0100101000: data <= 14'h3fea; 
        10'b0100101001: data <= 14'h0016; 
        10'b0100101010: data <= 14'h0037; 
        10'b0100101011: data <= 14'h0039; 
        10'b0100101100: data <= 14'h0033; 
        10'b0100101101: data <= 14'h0025; 
        10'b0100101110: data <= 14'h0036; 
        10'b0100101111: data <= 14'h004a; 
        10'b0100110000: data <= 14'h0023; 
        10'b0100110001: data <= 14'h3ff1; 
        10'b0100110010: data <= 14'h3ff1; 
        10'b0100110011: data <= 14'h3ff5; 
        10'b0100110100: data <= 14'h3ff8; 
        10'b0100110101: data <= 14'h3ff6; 
        10'b0100110110: data <= 14'h0004; 
        10'b0100110111: data <= 14'h3ffd; 
        10'b0100111000: data <= 14'h3fe4; 
        10'b0100111001: data <= 14'h3ffa; 
        10'b0100111010: data <= 14'h0004; 
        10'b0100111011: data <= 14'h0015; 
        10'b0100111100: data <= 14'h0010; 
        10'b0100111101: data <= 14'h3ffa; 
        10'b0100111110: data <= 14'h0006; 
        10'b0100111111: data <= 14'h0001; 
        10'b0101000000: data <= 14'h000b; 
        10'b0101000001: data <= 14'h3ff9; 
        10'b0101000010: data <= 14'h3fc5; 
        10'b0101000011: data <= 14'h3f93; 
        10'b0101000100: data <= 14'h3f99; 
        10'b0101000101: data <= 14'h3fd8; 
        10'b0101000110: data <= 14'h3ffb; 
        10'b0101000111: data <= 14'h001d; 
        10'b0101001000: data <= 14'h002e; 
        10'b0101001001: data <= 14'h002b; 
        10'b0101001010: data <= 14'h003b; 
        10'b0101001011: data <= 14'h0043; 
        10'b0101001100: data <= 14'h0030; 
        10'b0101001101: data <= 14'h3ff7; 
        10'b0101001110: data <= 14'h3fff; 
        10'b0101001111: data <= 14'h3ff4; 
        10'b0101010000: data <= 14'h3ff8; 
        10'b0101010001: data <= 14'h3ffd; 
        10'b0101010010: data <= 14'h3ffc; 
        10'b0101010011: data <= 14'h3ffd; 
        10'b0101010100: data <= 14'h3ff0; 
        10'b0101010101: data <= 14'h0003; 
        10'b0101010110: data <= 14'h0017; 
        10'b0101010111: data <= 14'h0018; 
        10'b0101011000: data <= 14'h000c; 
        10'b0101011001: data <= 14'h3ffd; 
        10'b0101011010: data <= 14'h0010; 
        10'b0101011011: data <= 14'h000c; 
        10'b0101011100: data <= 14'h0015; 
        10'b0101011101: data <= 14'h3fee; 
        10'b0101011110: data <= 14'h3f8c; 
        10'b0101011111: data <= 14'h3f70; 
        10'b0101100000: data <= 14'h3f71; 
        10'b0101100001: data <= 14'h3fb2; 
        10'b0101100010: data <= 14'h3ff2; 
        10'b0101100011: data <= 14'h3ffa; 
        10'b0101100100: data <= 14'h0007; 
        10'b0101100101: data <= 14'h0014; 
        10'b0101100110: data <= 14'h004c; 
        10'b0101100111: data <= 14'h0046; 
        10'b0101101000: data <= 14'h0030; 
        10'b0101101001: data <= 14'h0002; 
        10'b0101101010: data <= 14'h3ff8; 
        10'b0101101011: data <= 14'h3ff8; 
        10'b0101101100: data <= 14'h3ff5; 
        10'b0101101101: data <= 14'h0000; 
        10'b0101101110: data <= 14'h0004; 
        10'b0101101111: data <= 14'h3ff5; 
        10'b0101110000: data <= 14'h3ffc; 
        10'b0101110001: data <= 14'h000e; 
        10'b0101110010: data <= 14'h001c; 
        10'b0101110011: data <= 14'h0024; 
        10'b0101110100: data <= 14'h001b; 
        10'b0101110101: data <= 14'h0013; 
        10'b0101110110: data <= 14'h001a; 
        10'b0101110111: data <= 14'h0014; 
        10'b0101111000: data <= 14'h000f; 
        10'b0101111001: data <= 14'h3fb9; 
        10'b0101111010: data <= 14'h3f8c; 
        10'b0101111011: data <= 14'h3f6c; 
        10'b0101111100: data <= 14'h3f87; 
        10'b0101111101: data <= 14'h3fc4; 
        10'b0101111110: data <= 14'h3fe3; 
        10'b0101111111: data <= 14'h3fd9; 
        10'b0110000000: data <= 14'h3fe2; 
        10'b0110000001: data <= 14'h000d; 
        10'b0110000010: data <= 14'h0032; 
        10'b0110000011: data <= 14'h004e; 
        10'b0110000100: data <= 14'h002d; 
        10'b0110000101: data <= 14'h0007; 
        10'b0110000110: data <= 14'h0000; 
        10'b0110000111: data <= 14'h0004; 
        10'b0110001000: data <= 14'h3ffe; 
        10'b0110001001: data <= 14'h0003; 
        10'b0110001010: data <= 14'h3ff7; 
        10'b0110001011: data <= 14'h3ffa; 
        10'b0110001100: data <= 14'h3ff2; 
        10'b0110001101: data <= 14'h0025; 
        10'b0110001110: data <= 14'h0030; 
        10'b0110001111: data <= 14'h003a; 
        10'b0110010000: data <= 14'h001c; 
        10'b0110010001: data <= 14'h0021; 
        10'b0110010010: data <= 14'h0031; 
        10'b0110010011: data <= 14'h001c; 
        10'b0110010100: data <= 14'h0007; 
        10'b0110010101: data <= 14'h3fc3; 
        10'b0110010110: data <= 14'h3f77; 
        10'b0110010111: data <= 14'h3f6c; 
        10'b0110011000: data <= 14'h3f8a; 
        10'b0110011001: data <= 14'h3fc0; 
        10'b0110011010: data <= 14'h3fe4; 
        10'b0110011011: data <= 14'h3fde; 
        10'b0110011100: data <= 14'h0003; 
        10'b0110011101: data <= 14'h001c; 
        10'b0110011110: data <= 14'h0021; 
        10'b0110011111: data <= 14'h004f; 
        10'b0110100000: data <= 14'h0029; 
        10'b0110100001: data <= 14'h3ff8; 
        10'b0110100010: data <= 14'h3ffc; 
        10'b0110100011: data <= 14'h3ff7; 
        10'b0110100100: data <= 14'h0005; 
        10'b0110100101: data <= 14'h0003; 
        10'b0110100110: data <= 14'h3ff8; 
        10'b0110100111: data <= 14'h3ffe; 
        10'b0110101000: data <= 14'h3fff; 
        10'b0110101001: data <= 14'h0034; 
        10'b0110101010: data <= 14'h0026; 
        10'b0110101011: data <= 14'h0034; 
        10'b0110101100: data <= 14'h0024; 
        10'b0110101101: data <= 14'h002f; 
        10'b0110101110: data <= 14'h003c; 
        10'b0110101111: data <= 14'h0011; 
        10'b0110110000: data <= 14'h3fd3; 
        10'b0110110001: data <= 14'h3f8d; 
        10'b0110110010: data <= 14'h3f67; 
        10'b0110110011: data <= 14'h3f6e; 
        10'b0110110100: data <= 14'h3f9d; 
        10'b0110110101: data <= 14'h3fd0; 
        10'b0110110110: data <= 14'h3fee; 
        10'b0110110111: data <= 14'h3fef; 
        10'b0110111000: data <= 14'h000f; 
        10'b0110111001: data <= 14'h000d; 
        10'b0110111010: data <= 14'h0032; 
        10'b0110111011: data <= 14'h003b; 
        10'b0110111100: data <= 14'h001f; 
        10'b0110111101: data <= 14'h3ffd; 
        10'b0110111110: data <= 14'h0001; 
        10'b0110111111: data <= 14'h3ff8; 
        10'b0111000000: data <= 14'h0001; 
        10'b0111000001: data <= 14'h0006; 
        10'b0111000010: data <= 14'h3ff4; 
        10'b0111000011: data <= 14'h3ffa; 
        10'b0111000100: data <= 14'h0009; 
        10'b0111000101: data <= 14'h002f; 
        10'b0111000110: data <= 14'h003a; 
        10'b0111000111: data <= 14'h002d; 
        10'b0111001000: data <= 14'h001f; 
        10'b0111001001: data <= 14'h0020; 
        10'b0111001010: data <= 14'h0035; 
        10'b0111001011: data <= 14'h3ff9; 
        10'b0111001100: data <= 14'h3fa8; 
        10'b0111001101: data <= 14'h3f68; 
        10'b0111001110: data <= 14'h3f6c; 
        10'b0111001111: data <= 14'h3f8a; 
        10'b0111010000: data <= 14'h3fc1; 
        10'b0111010001: data <= 14'h3fe3; 
        10'b0111010010: data <= 14'h0000; 
        10'b0111010011: data <= 14'h000a; 
        10'b0111010100: data <= 14'h0016; 
        10'b0111010101: data <= 14'h0021; 
        10'b0111010110: data <= 14'h002d; 
        10'b0111010111: data <= 14'h002b; 
        10'b0111011000: data <= 14'h0010; 
        10'b0111011001: data <= 14'h0001; 
        10'b0111011010: data <= 14'h3ffb; 
        10'b0111011011: data <= 14'h3ff9; 
        10'b0111011100: data <= 14'h3ffc; 
        10'b0111011101: data <= 14'h0001; 
        10'b0111011110: data <= 14'h3ff6; 
        10'b0111011111: data <= 14'h3fed; 
        10'b0111100000: data <= 14'h0002; 
        10'b0111100001: data <= 14'h0021; 
        10'b0111100010: data <= 14'h002a; 
        10'b0111100011: data <= 14'h0029; 
        10'b0111100100: data <= 14'h000d; 
        10'b0111100101: data <= 14'h0021; 
        10'b0111100110: data <= 14'h0034; 
        10'b0111100111: data <= 14'h3ff8; 
        10'b0111101000: data <= 14'h3f97; 
        10'b0111101001: data <= 14'h3f6a; 
        10'b0111101010: data <= 14'h3f7c; 
        10'b0111101011: data <= 14'h3fb1; 
        10'b0111101100: data <= 14'h3ff6; 
        10'b0111101101: data <= 14'h0014; 
        10'b0111101110: data <= 14'h001d; 
        10'b0111101111: data <= 14'h001b; 
        10'b0111110000: data <= 14'h0022; 
        10'b0111110001: data <= 14'h001a; 
        10'b0111110010: data <= 14'h0015; 
        10'b0111110011: data <= 14'h0017; 
        10'b0111110100: data <= 14'h3fff; 
        10'b0111110101: data <= 14'h3ffd; 
        10'b0111110110: data <= 14'h0002; 
        10'b0111110111: data <= 14'h3ff8; 
        10'b0111111000: data <= 14'h3ffa; 
        10'b0111111001: data <= 14'h0002; 
        10'b0111111010: data <= 14'h3ffc; 
        10'b0111111011: data <= 14'h3ff9; 
        10'b0111111100: data <= 14'h3ffc; 
        10'b0111111101: data <= 14'h0015; 
        10'b0111111110: data <= 14'h002b; 
        10'b0111111111: data <= 14'h0019; 
        10'b1000000000: data <= 14'h000f; 
        10'b1000000001: data <= 14'h002b; 
        10'b1000000010: data <= 14'h0053; 
        10'b1000000011: data <= 14'h0003; 
        10'b1000000100: data <= 14'h3fbd; 
        10'b1000000101: data <= 14'h3f94; 
        10'b1000000110: data <= 14'h3fb5; 
        10'b1000000111: data <= 14'h3fe9; 
        10'b1000001000: data <= 14'h0018; 
        10'b1000001001: data <= 14'h001a; 
        10'b1000001010: data <= 14'h001b; 
        10'b1000001011: data <= 14'h000e; 
        10'b1000001100: data <= 14'h0007; 
        10'b1000001101: data <= 14'h000c; 
        10'b1000001110: data <= 14'h0017; 
        10'b1000001111: data <= 14'h000e; 
        10'b1000010000: data <= 14'h3ffe; 
        10'b1000010001: data <= 14'h3ff9; 
        10'b1000010010: data <= 14'h0001; 
        10'b1000010011: data <= 14'h3ffc; 
        10'b1000010100: data <= 14'h3ffd; 
        10'b1000010101: data <= 14'h3ffb; 
        10'b1000010110: data <= 14'h3ffc; 
        10'b1000010111: data <= 14'h3fed; 
        10'b1000011000: data <= 14'h0008; 
        10'b1000011001: data <= 14'h0017; 
        10'b1000011010: data <= 14'h0038; 
        10'b1000011011: data <= 14'h0033; 
        10'b1000011100: data <= 14'h0028; 
        10'b1000011101: data <= 14'h0035; 
        10'b1000011110: data <= 14'h0053; 
        10'b1000011111: data <= 14'h003a; 
        10'b1000100000: data <= 14'h000c; 
        10'b1000100001: data <= 14'h3fe5; 
        10'b1000100010: data <= 14'h3ff4; 
        10'b1000100011: data <= 14'h3ff8; 
        10'b1000100100: data <= 14'h000d; 
        10'b1000100101: data <= 14'h3ffa; 
        10'b1000100110: data <= 14'h3ff5; 
        10'b1000100111: data <= 14'h3ff9; 
        10'b1000101000: data <= 14'h000d; 
        10'b1000101001: data <= 14'h000c; 
        10'b1000101010: data <= 14'h0017; 
        10'b1000101011: data <= 14'h3ffd; 
        10'b1000101100: data <= 14'h0003; 
        10'b1000101101: data <= 14'h3ffb; 
        10'b1000101110: data <= 14'h3ff4; 
        10'b1000101111: data <= 14'h0004; 
        10'b1000110000: data <= 14'h0004; 
        10'b1000110001: data <= 14'h0005; 
        10'b1000110010: data <= 14'h3ffc; 
        10'b1000110011: data <= 14'h3ff7; 
        10'b1000110100: data <= 14'h3ffb; 
        10'b1000110101: data <= 14'h0018; 
        10'b1000110110: data <= 14'h002d; 
        10'b1000110111: data <= 14'h0021; 
        10'b1000111000: data <= 14'h0029; 
        10'b1000111001: data <= 14'h0032; 
        10'b1000111010: data <= 14'h004e; 
        10'b1000111011: data <= 14'h004e; 
        10'b1000111100: data <= 14'h0027; 
        10'b1000111101: data <= 14'h000c; 
        10'b1000111110: data <= 14'h3ff8; 
        10'b1000111111: data <= 14'h0006; 
        10'b1001000000: data <= 14'h0005; 
        10'b1001000001: data <= 14'h3ff5; 
        10'b1001000010: data <= 14'h3ff7; 
        10'b1001000011: data <= 14'h3ff4; 
        10'b1001000100: data <= 14'h0006; 
        10'b1001000101: data <= 14'h0008; 
        10'b1001000110: data <= 14'h000c; 
        10'b1001000111: data <= 14'h0004; 
        10'b1001001000: data <= 14'h3ff9; 
        10'b1001001001: data <= 14'h3ffe; 
        10'b1001001010: data <= 14'h3ff6; 
        10'b1001001011: data <= 14'h3ffb; 
        10'b1001001100: data <= 14'h3ff9; 
        10'b1001001101: data <= 14'h3ff5; 
        10'b1001001110: data <= 14'h3ffc; 
        10'b1001001111: data <= 14'h3ff9; 
        10'b1001010000: data <= 14'h3ffc; 
        10'b1001010001: data <= 14'h0006; 
        10'b1001010010: data <= 14'h001c; 
        10'b1001010011: data <= 14'h002d; 
        10'b1001010100: data <= 14'h0020; 
        10'b1001010101: data <= 14'h0022; 
        10'b1001010110: data <= 14'h0043; 
        10'b1001010111: data <= 14'h004c; 
        10'b1001011000: data <= 14'h0032; 
        10'b1001011001: data <= 14'h0013; 
        10'b1001011010: data <= 14'h0007; 
        10'b1001011011: data <= 14'h0001; 
        10'b1001011100: data <= 14'h3fff; 
        10'b1001011101: data <= 14'h3feb; 
        10'b1001011110: data <= 14'h3ff0; 
        10'b1001011111: data <= 14'h3ff7; 
        10'b1001100000: data <= 14'h0008; 
        10'b1001100001: data <= 14'h3fff; 
        10'b1001100010: data <= 14'h3ff7; 
        10'b1001100011: data <= 14'h3ff1; 
        10'b1001100100: data <= 14'h3ffc; 
        10'b1001100101: data <= 14'h3ffb; 
        10'b1001100110: data <= 14'h3ff9; 
        10'b1001100111: data <= 14'h3ffa; 
        10'b1001101000: data <= 14'h3ff7; 
        10'b1001101001: data <= 14'h0001; 
        10'b1001101010: data <= 14'h0001; 
        10'b1001101011: data <= 14'h3ffb; 
        10'b1001101100: data <= 14'h3ff7; 
        10'b1001101101: data <= 14'h0003; 
        10'b1001101110: data <= 14'h0014; 
        10'b1001101111: data <= 14'h0011; 
        10'b1001110000: data <= 14'h0033; 
        10'b1001110001: data <= 14'h0029; 
        10'b1001110010: data <= 14'h002d; 
        10'b1001110011: data <= 14'h0036; 
        10'b1001110100: data <= 14'h002e; 
        10'b1001110101: data <= 14'h003b; 
        10'b1001110110: data <= 14'h001a; 
        10'b1001110111: data <= 14'h001a; 
        10'b1001111000: data <= 14'h000e; 
        10'b1001111001: data <= 14'h3ff4; 
        10'b1001111010: data <= 14'h3ff6; 
        10'b1001111011: data <= 14'h3fff; 
        10'b1001111100: data <= 14'h3ff2; 
        10'b1001111101: data <= 14'h3ff2; 
        10'b1001111110: data <= 14'h3ff9; 
        10'b1001111111: data <= 14'h3ff9; 
        10'b1010000000: data <= 14'h3ffd; 
        10'b1010000001: data <= 14'h3ffb; 
        10'b1010000010: data <= 14'h3ffa; 
        10'b1010000011: data <= 14'h3ffd; 
        10'b1010000100: data <= 14'h3ff7; 
        10'b1010000101: data <= 14'h3ffe; 
        10'b1010000110: data <= 14'h0000; 
        10'b1010000111: data <= 14'h3ff5; 
        10'b1010001000: data <= 14'h3ff5; 
        10'b1010001001: data <= 14'h3ffd; 
        10'b1010001010: data <= 14'h3fff; 
        10'b1010001011: data <= 14'h000e; 
        10'b1010001100: data <= 14'h0014; 
        10'b1010001101: data <= 14'h002f; 
        10'b1010001110: data <= 14'h0038; 
        10'b1010001111: data <= 14'h0045; 
        10'b1010010000: data <= 14'h0044; 
        10'b1010010001: data <= 14'h0029; 
        10'b1010010010: data <= 14'h0021; 
        10'b1010010011: data <= 14'h0012; 
        10'b1010010100: data <= 14'h0008; 
        10'b1010010101: data <= 14'h3fff; 
        10'b1010010110: data <= 14'h3fe6; 
        10'b1010010111: data <= 14'h3fe0; 
        10'b1010011000: data <= 14'h3fe7; 
        10'b1010011001: data <= 14'h3ff4; 
        10'b1010011010: data <= 14'h3ff6; 
        10'b1010011011: data <= 14'h3fff; 
        10'b1010011100: data <= 14'h3ffc; 
        10'b1010011101: data <= 14'h0003; 
        10'b1010011110: data <= 14'h3ffb; 
        10'b1010011111: data <= 14'h3ff5; 
        10'b1010100000: data <= 14'h3ffb; 
        10'b1010100001: data <= 14'h3ffe; 
        10'b1010100010: data <= 14'h3ff5; 
        10'b1010100011: data <= 14'h0000; 
        10'b1010100100: data <= 14'h3ffd; 
        10'b1010100101: data <= 14'h3ffd; 
        10'b1010100110: data <= 14'h3ff3; 
        10'b1010100111: data <= 14'h3fee; 
        10'b1010101000: data <= 14'h3ff6; 
        10'b1010101001: data <= 14'h3ff7; 
        10'b1010101010: data <= 14'h000a; 
        10'b1010101011: data <= 14'h0008; 
        10'b1010101100: data <= 14'h0013; 
        10'b1010101101: data <= 14'h001c; 
        10'b1010101110: data <= 14'h000f; 
        10'b1010101111: data <= 14'h3ff5; 
        10'b1010110000: data <= 14'h3fef; 
        10'b1010110001: data <= 14'h3feb; 
        10'b1010110010: data <= 14'h3fee; 
        10'b1010110011: data <= 14'h3fe7; 
        10'b1010110100: data <= 14'h3fe8; 
        10'b1010110101: data <= 14'h3fea; 
        10'b1010110110: data <= 14'h3ffc; 
        10'b1010110111: data <= 14'h3ffa; 
        10'b1010111000: data <= 14'h3ff7; 
        10'b1010111001: data <= 14'h3ff9; 
        10'b1010111010: data <= 14'h0001; 
        10'b1010111011: data <= 14'h3ff8; 
        10'b1010111100: data <= 14'h3ff9; 
        10'b1010111101: data <= 14'h0006; 
        10'b1010111110: data <= 14'h3ffd; 
        10'b1010111111: data <= 14'h0005; 
        10'b1011000000: data <= 14'h0006; 
        10'b1011000001: data <= 14'h0000; 
        10'b1011000010: data <= 14'h3ff4; 
        10'b1011000011: data <= 14'h3ffb; 
        10'b1011000100: data <= 14'h3fe9; 
        10'b1011000101: data <= 14'h3fea; 
        10'b1011000110: data <= 14'h3fe4; 
        10'b1011000111: data <= 14'h3fdc; 
        10'b1011001000: data <= 14'h3fd7; 
        10'b1011001001: data <= 14'h3fdb; 
        10'b1011001010: data <= 14'h3fd5; 
        10'b1011001011: data <= 14'h3fd9; 
        10'b1011001100: data <= 14'h3fdb; 
        10'b1011001101: data <= 14'h3fea; 
        10'b1011001110: data <= 14'h3fee; 
        10'b1011001111: data <= 14'h3ff0; 
        10'b1011010000: data <= 14'h3fef; 
        10'b1011010001: data <= 14'h3ff0; 
        10'b1011010010: data <= 14'h3ffb; 
        10'b1011010011: data <= 14'h0006; 
        10'b1011010100: data <= 14'h0003; 
        10'b1011010101: data <= 14'h3ffc; 
        10'b1011010110: data <= 14'h3ffa; 
        10'b1011010111: data <= 14'h3ffe; 
        10'b1011011000: data <= 14'h0005; 
        10'b1011011001: data <= 14'h0005; 
        10'b1011011010: data <= 14'h3ffb; 
        10'b1011011011: data <= 14'h0000; 
        10'b1011011100: data <= 14'h3ffa; 
        10'b1011011101: data <= 14'h3ffb; 
        10'b1011011110: data <= 14'h3ff5; 
        10'b1011011111: data <= 14'h0002; 
        10'b1011100000: data <= 14'h3ffa; 
        10'b1011100001: data <= 14'h3fec; 
        10'b1011100010: data <= 14'h3fec; 
        10'b1011100011: data <= 14'h3fee; 
        10'b1011100100: data <= 14'h3ff9; 
        10'b1011100101: data <= 14'h3fee; 
        10'b1011100110: data <= 14'h3fef; 
        10'b1011100111: data <= 14'h3ffa; 
        10'b1011101000: data <= 14'h3fee; 
        10'b1011101001: data <= 14'h3ff1; 
        10'b1011101010: data <= 14'h3ff5; 
        10'b1011101011: data <= 14'h3ff2; 
        10'b1011101100: data <= 14'h3ff9; 
        10'b1011101101: data <= 14'h3ff0; 
        10'b1011101110: data <= 14'h3ff2; 
        10'b1011101111: data <= 14'h0005; 
        10'b1011110000: data <= 14'h3ff7; 
        10'b1011110001: data <= 14'h0002; 
        10'b1011110010: data <= 14'h0004; 
        10'b1011110011: data <= 14'h3fff; 
        10'b1011110100: data <= 14'h3ff7; 
        10'b1011110101: data <= 14'h0004; 
        10'b1011110110: data <= 14'h3ffe; 
        10'b1011110111: data <= 14'h3ffb; 
        10'b1011111000: data <= 14'h0005; 
        10'b1011111001: data <= 14'h0001; 
        10'b1011111010: data <= 14'h0002; 
        10'b1011111011: data <= 14'h3ff5; 
        10'b1011111100: data <= 14'h0006; 
        10'b1011111101: data <= 14'h0005; 
        10'b1011111110: data <= 14'h0002; 
        10'b1011111111: data <= 14'h0004; 
        10'b1100000000: data <= 14'h3ffd; 
        10'b1100000001: data <= 14'h3ff9; 
        10'b1100000010: data <= 14'h0004; 
        10'b1100000011: data <= 14'h3ff6; 
        10'b1100000100: data <= 14'h3ffc; 
        10'b1100000101: data <= 14'h3ff9; 
        10'b1100000110: data <= 14'h3ffe; 
        10'b1100000111: data <= 14'h3ffa; 
        10'b1100001000: data <= 14'h3ff4; 
        10'b1100001001: data <= 14'h3ff6; 
        10'b1100001010: data <= 14'h3ff1; 
        10'b1100001011: data <= 14'h3ffd; 
        10'b1100001100: data <= 14'h0002; 
        10'b1100001101: data <= 14'h3ff7; 
        10'b1100001110: data <= 14'h3ff4; 
        10'b1100001111: data <= 14'h0003; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 9) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 15'h7fef; 
        10'b0000000001: data <= 15'h0009; 
        10'b0000000010: data <= 15'h7ffb; 
        10'b0000000011: data <= 15'h7ffe; 
        10'b0000000100: data <= 15'h000b; 
        10'b0000000101: data <= 15'h7fff; 
        10'b0000000110: data <= 15'h7ff5; 
        10'b0000000111: data <= 15'h7ff5; 
        10'b0000001000: data <= 15'h7ffd; 
        10'b0000001001: data <= 15'h7ffa; 
        10'b0000001010: data <= 15'h000c; 
        10'b0000001011: data <= 15'h7fff; 
        10'b0000001100: data <= 15'h0006; 
        10'b0000001101: data <= 15'h7ff0; 
        10'b0000001110: data <= 15'h7fff; 
        10'b0000001111: data <= 15'h7fea; 
        10'b0000010000: data <= 15'h7fee; 
        10'b0000010001: data <= 15'h7ffb; 
        10'b0000010010: data <= 15'h7fed; 
        10'b0000010011: data <= 15'h000c; 
        10'b0000010100: data <= 15'h7fed; 
        10'b0000010101: data <= 15'h7ffa; 
        10'b0000010110: data <= 15'h7fec; 
        10'b0000010111: data <= 15'h7ffe; 
        10'b0000011000: data <= 15'h0006; 
        10'b0000011001: data <= 15'h7ffc; 
        10'b0000011010: data <= 15'h7fff; 
        10'b0000011011: data <= 15'h7fff; 
        10'b0000011100: data <= 15'h0007; 
        10'b0000011101: data <= 15'h0009; 
        10'b0000011110: data <= 15'h0003; 
        10'b0000011111: data <= 15'h7fed; 
        10'b0000100000: data <= 15'h7fec; 
        10'b0000100001: data <= 15'h0001; 
        10'b0000100010: data <= 15'h7ff0; 
        10'b0000100011: data <= 15'h7ffb; 
        10'b0000100100: data <= 15'h7ff3; 
        10'b0000100101: data <= 15'h7fe9; 
        10'b0000100110: data <= 15'h7ff1; 
        10'b0000100111: data <= 15'h0001; 
        10'b0000101000: data <= 15'h000e; 
        10'b0000101001: data <= 15'h7fed; 
        10'b0000101010: data <= 15'h7ff6; 
        10'b0000101011: data <= 15'h0006; 
        10'b0000101100: data <= 15'h7ff0; 
        10'b0000101101: data <= 15'h7fea; 
        10'b0000101110: data <= 15'h0004; 
        10'b0000101111: data <= 15'h000a; 
        10'b0000110000: data <= 15'h7fef; 
        10'b0000110001: data <= 15'h0005; 
        10'b0000110010: data <= 15'h7ff2; 
        10'b0000110011: data <= 15'h7fee; 
        10'b0000110100: data <= 15'h7ffc; 
        10'b0000110101: data <= 15'h0001; 
        10'b0000110110: data <= 15'h7ffa; 
        10'b0000110111: data <= 15'h000c; 
        10'b0000111000: data <= 15'h7feb; 
        10'b0000111001: data <= 15'h7ff3; 
        10'b0000111010: data <= 15'h7ff2; 
        10'b0000111011: data <= 15'h0006; 
        10'b0000111100: data <= 15'h0002; 
        10'b0000111101: data <= 15'h7feb; 
        10'b0000111110: data <= 15'h7ffb; 
        10'b0000111111: data <= 15'h000b; 
        10'b0001000000: data <= 15'h7ff9; 
        10'b0001000001: data <= 15'h7ff1; 
        10'b0001000010: data <= 15'h7ff1; 
        10'b0001000011: data <= 15'h7fe7; 
        10'b0001000100: data <= 15'h7fe5; 
        10'b0001000101: data <= 15'h7ff7; 
        10'b0001000110: data <= 15'h7fe4; 
        10'b0001000111: data <= 15'h7fdc; 
        10'b0001001000: data <= 15'h7fe6; 
        10'b0001001001: data <= 15'h7ff9; 
        10'b0001001010: data <= 15'h7fea; 
        10'b0001001011: data <= 15'h7fe3; 
        10'b0001001100: data <= 15'h7ffb; 
        10'b0001001101: data <= 15'h0009; 
        10'b0001001110: data <= 15'h0002; 
        10'b0001001111: data <= 15'h7ff0; 
        10'b0001010000: data <= 15'h000b; 
        10'b0001010001: data <= 15'h7fe9; 
        10'b0001010010: data <= 15'h7ffa; 
        10'b0001010011: data <= 15'h0005; 
        10'b0001010100: data <= 15'h7feb; 
        10'b0001010101: data <= 15'h7ffb; 
        10'b0001010110: data <= 15'h000c; 
        10'b0001010111: data <= 15'h7feb; 
        10'b0001011000: data <= 15'h7ff1; 
        10'b0001011001: data <= 15'h000a; 
        10'b0001011010: data <= 15'h0004; 
        10'b0001011011: data <= 15'h0000; 
        10'b0001011100: data <= 15'h0002; 
        10'b0001011101: data <= 15'h7ffb; 
        10'b0001011110: data <= 15'h7ff9; 
        10'b0001011111: data <= 15'h7fe4; 
        10'b0001100000: data <= 15'h7fd9; 
        10'b0001100001: data <= 15'h7fea; 
        10'b0001100010: data <= 15'h7fe2; 
        10'b0001100011: data <= 15'h7fde; 
        10'b0001100100: data <= 15'h0006; 
        10'b0001100101: data <= 15'h0003; 
        10'b0001100110: data <= 15'h7fda; 
        10'b0001100111: data <= 15'h7fdf; 
        10'b0001101000: data <= 15'h7fd1; 
        10'b0001101001: data <= 15'h7fdf; 
        10'b0001101010: data <= 15'h7fd8; 
        10'b0001101011: data <= 15'h7fe4; 
        10'b0001101100: data <= 15'h7fed; 
        10'b0001101101: data <= 15'h0007; 
        10'b0001101110: data <= 15'h0007; 
        10'b0001101111: data <= 15'h7ff5; 
        10'b0001110000: data <= 15'h0003; 
        10'b0001110001: data <= 15'h7fea; 
        10'b0001110010: data <= 15'h7ff1; 
        10'b0001110011: data <= 15'h7feb; 
        10'b0001110100: data <= 15'h7fe8; 
        10'b0001110101: data <= 15'h7ffd; 
        10'b0001110110: data <= 15'h7ffa; 
        10'b0001110111: data <= 15'h7feb; 
        10'b0001111000: data <= 15'h7ff9; 
        10'b0001111001: data <= 15'h7ffb; 
        10'b0001111010: data <= 15'h7fdd; 
        10'b0001111011: data <= 15'h7fde; 
        10'b0001111100: data <= 15'h7fde; 
        10'b0001111101: data <= 15'h7fe0; 
        10'b0001111110: data <= 15'h7ff7; 
        10'b0001111111: data <= 15'h7ffd; 
        10'b0010000000: data <= 15'h7fe5; 
        10'b0010000001: data <= 15'h7fe7; 
        10'b0010000010: data <= 15'h7fe6; 
        10'b0010000011: data <= 15'h7fdc; 
        10'b0010000100: data <= 15'h7ff1; 
        10'b0010000101: data <= 15'h7fd2; 
        10'b0010000110: data <= 15'h7fee; 
        10'b0010000111: data <= 15'h7ffd; 
        10'b0010001000: data <= 15'h7fec; 
        10'b0010001001: data <= 15'h7ff7; 
        10'b0010001010: data <= 15'h7ff4; 
        10'b0010001011: data <= 15'h7ffe; 
        10'b0010001100: data <= 15'h0006; 
        10'b0010001101: data <= 15'h7ff6; 
        10'b0010001110: data <= 15'h0000; 
        10'b0010001111: data <= 15'h7fed; 
        10'b0010010000: data <= 15'h7ffb; 
        10'b0010010001: data <= 15'h7ff7; 
        10'b0010010010: data <= 15'h7ff9; 
        10'b0010010011: data <= 15'h7ff2; 
        10'b0010010100: data <= 15'h7ffa; 
        10'b0010010101: data <= 15'h7fe6; 
        10'b0010010110: data <= 15'h7ff4; 
        10'b0010010111: data <= 15'h0008; 
        10'b0010011000: data <= 15'h001e; 
        10'b0010011001: data <= 15'h0041; 
        10'b0010011010: data <= 15'h004f; 
        10'b0010011011: data <= 15'h004e; 
        10'b0010011100: data <= 15'h0058; 
        10'b0010011101: data <= 15'h005e; 
        10'b0010011110: data <= 15'h0064; 
        10'b0010011111: data <= 15'h0023; 
        10'b0010100000: data <= 15'h0006; 
        10'b0010100001: data <= 15'h0010; 
        10'b0010100010: data <= 15'h7ff8; 
        10'b0010100011: data <= 15'h7fff; 
        10'b0010100100: data <= 15'h7fd5; 
        10'b0010100101: data <= 15'h7fe1; 
        10'b0010100110: data <= 15'h7ffe; 
        10'b0010100111: data <= 15'h7ff0; 
        10'b0010101000: data <= 15'h7ff7; 
        10'b0010101001: data <= 15'h7ffc; 
        10'b0010101010: data <= 15'h0002; 
        10'b0010101011: data <= 15'h7ff9; 
        10'b0010101100: data <= 15'h0000; 
        10'b0010101101: data <= 15'h0001; 
        10'b0010101110: data <= 15'h0002; 
        10'b0010101111: data <= 15'h7fff; 
        10'b0010110000: data <= 15'h7feb; 
        10'b0010110001: data <= 15'h7fdc; 
        10'b0010110010: data <= 15'h0014; 
        10'b0010110011: data <= 15'h7ffd; 
        10'b0010110100: data <= 15'h0036; 
        10'b0010110101: data <= 15'h0030; 
        10'b0010110110: data <= 15'h002e; 
        10'b0010110111: data <= 15'h0044; 
        10'b0010111000: data <= 15'h0053; 
        10'b0010111001: data <= 15'h0075; 
        10'b0010111010: data <= 15'h006d; 
        10'b0010111011: data <= 15'h005d; 
        10'b0010111100: data <= 15'h005a; 
        10'b0010111101: data <= 15'h0066; 
        10'b0010111110: data <= 15'h003a; 
        10'b0010111111: data <= 15'h0015; 
        10'b0011000000: data <= 15'h7fd4; 
        10'b0011000001: data <= 15'h7fd2; 
        10'b0011000010: data <= 15'h7fe1; 
        10'b0011000011: data <= 15'h0005; 
        10'b0011000100: data <= 15'h000b; 
        10'b0011000101: data <= 15'h0002; 
        10'b0011000110: data <= 15'h7ffe; 
        10'b0011000111: data <= 15'h7fe5; 
        10'b0011001000: data <= 15'h7fd6; 
        10'b0011001001: data <= 15'h7ffc; 
        10'b0011001010: data <= 15'h7fef; 
        10'b0011001011: data <= 15'h0000; 
        10'b0011001100: data <= 15'h7fec; 
        10'b0011001101: data <= 15'h7ffa; 
        10'b0011001110: data <= 15'h0004; 
        10'b0011001111: data <= 15'h0027; 
        10'b0011010000: data <= 15'h0050; 
        10'b0011010001: data <= 15'h004a; 
        10'b0011010010: data <= 15'h001e; 
        10'b0011010011: data <= 15'h002f; 
        10'b0011010100: data <= 15'h0043; 
        10'b0011010101: data <= 15'h007e; 
        10'b0011010110: data <= 15'h005d; 
        10'b0011010111: data <= 15'h0051; 
        10'b0011011000: data <= 15'h0021; 
        10'b0011011001: data <= 15'h0040; 
        10'b0011011010: data <= 15'h0046; 
        10'b0011011011: data <= 15'h0024; 
        10'b0011011100: data <= 15'h7fe5; 
        10'b0011011101: data <= 15'h7fd3; 
        10'b0011011110: data <= 15'h7fd8; 
        10'b0011011111: data <= 15'h7ffe; 
        10'b0011100000: data <= 15'h000c; 
        10'b0011100001: data <= 15'h0004; 
        10'b0011100010: data <= 15'h7ffb; 
        10'b0011100011: data <= 15'h0000; 
        10'b0011100100: data <= 15'h7fe1; 
        10'b0011100101: data <= 15'h7fe8; 
        10'b0011100110: data <= 15'h7fec; 
        10'b0011100111: data <= 15'h7fe8; 
        10'b0011101000: data <= 15'h7ff3; 
        10'b0011101001: data <= 15'h7ff2; 
        10'b0011101010: data <= 15'h0026; 
        10'b0011101011: data <= 15'h0028; 
        10'b0011101100: data <= 15'h0015; 
        10'b0011101101: data <= 15'h0009; 
        10'b0011101110: data <= 15'h000e; 
        10'b0011101111: data <= 15'h0039; 
        10'b0011110000: data <= 15'h00a5; 
        10'b0011110001: data <= 15'h0083; 
        10'b0011110010: data <= 15'h007a; 
        10'b0011110011: data <= 15'h0026; 
        10'b0011110100: data <= 15'h0020; 
        10'b0011110101: data <= 15'h001e; 
        10'b0011110110: data <= 15'h0048; 
        10'b0011110111: data <= 15'h007e; 
        10'b0011111000: data <= 15'h7ff2; 
        10'b0011111001: data <= 15'h7fd6; 
        10'b0011111010: data <= 15'h7ffc; 
        10'b0011111011: data <= 15'h7fea; 
        10'b0011111100: data <= 15'h7ffd; 
        10'b0011111101: data <= 15'h7ffe; 
        10'b0011111110: data <= 15'h0004; 
        10'b0011111111: data <= 15'h0003; 
        10'b0100000000: data <= 15'h7fd9; 
        10'b0100000001: data <= 15'h7fe4; 
        10'b0100000010: data <= 15'h7fd8; 
        10'b0100000011: data <= 15'h7fe9; 
        10'b0100000100: data <= 15'h7fe9; 
        10'b0100000101: data <= 15'h7ff4; 
        10'b0100000110: data <= 15'h001b; 
        10'b0100000111: data <= 15'h7fe9; 
        10'b0100001000: data <= 15'h000e; 
        10'b0100001001: data <= 15'h0029; 
        10'b0100001010: data <= 15'h0025; 
        10'b0100001011: data <= 15'h001f; 
        10'b0100001100: data <= 15'h005a; 
        10'b0100001101: data <= 15'h0079; 
        10'b0100001110: data <= 15'h008b; 
        10'b0100001111: data <= 15'h0050; 
        10'b0100010000: data <= 15'h0018; 
        10'b0100010001: data <= 15'h7ffb; 
        10'b0100010010: data <= 15'h003b; 
        10'b0100010011: data <= 15'h0080; 
        10'b0100010100: data <= 15'h0025; 
        10'b0100010101: data <= 15'h7fe0; 
        10'b0100010110: data <= 15'h0000; 
        10'b0100010111: data <= 15'h7ffc; 
        10'b0100011000: data <= 15'h7fec; 
        10'b0100011001: data <= 15'h000a; 
        10'b0100011010: data <= 15'h7fef; 
        10'b0100011011: data <= 15'h7fe1; 
        10'b0100011100: data <= 15'h7fe4; 
        10'b0100011101: data <= 15'h7fe9; 
        10'b0100011110: data <= 15'h7fed; 
        10'b0100011111: data <= 15'h0003; 
        10'b0100100000: data <= 15'h000d; 
        10'b0100100001: data <= 15'h7ffd; 
        10'b0100100010: data <= 15'h7fea; 
        10'b0100100011: data <= 15'h0007; 
        10'b0100100100: data <= 15'h0009; 
        10'b0100100101: data <= 15'h7ffb; 
        10'b0100100110: data <= 15'h7fd4; 
        10'b0100100111: data <= 15'h7fb5; 
        10'b0100101000: data <= 15'h7fd3; 
        10'b0100101001: data <= 15'h002b; 
        10'b0100101010: data <= 15'h006e; 
        10'b0100101011: data <= 15'h0072; 
        10'b0100101100: data <= 15'h0065; 
        10'b0100101101: data <= 15'h0049; 
        10'b0100101110: data <= 15'h006d; 
        10'b0100101111: data <= 15'h0095; 
        10'b0100110000: data <= 15'h0047; 
        10'b0100110001: data <= 15'h7fe3; 
        10'b0100110010: data <= 15'h7fe3; 
        10'b0100110011: data <= 15'h7fea; 
        10'b0100110100: data <= 15'h7ff1; 
        10'b0100110101: data <= 15'h7fec; 
        10'b0100110110: data <= 15'h0009; 
        10'b0100110111: data <= 15'h7ffa; 
        10'b0100111000: data <= 15'h7fc8; 
        10'b0100111001: data <= 15'h7ff4; 
        10'b0100111010: data <= 15'h0009; 
        10'b0100111011: data <= 15'h002a; 
        10'b0100111100: data <= 15'h0020; 
        10'b0100111101: data <= 15'h7ff4; 
        10'b0100111110: data <= 15'h000b; 
        10'b0100111111: data <= 15'h0001; 
        10'b0101000000: data <= 15'h0016; 
        10'b0101000001: data <= 15'h7ff1; 
        10'b0101000010: data <= 15'h7f8a; 
        10'b0101000011: data <= 15'h7f25; 
        10'b0101000100: data <= 15'h7f32; 
        10'b0101000101: data <= 15'h7fb0; 
        10'b0101000110: data <= 15'h7ff5; 
        10'b0101000111: data <= 15'h003a; 
        10'b0101001000: data <= 15'h005d; 
        10'b0101001001: data <= 15'h0056; 
        10'b0101001010: data <= 15'h0075; 
        10'b0101001011: data <= 15'h0085; 
        10'b0101001100: data <= 15'h0060; 
        10'b0101001101: data <= 15'h7fee; 
        10'b0101001110: data <= 15'h7fff; 
        10'b0101001111: data <= 15'h7fe8; 
        10'b0101010000: data <= 15'h7ff0; 
        10'b0101010001: data <= 15'h7ffb; 
        10'b0101010010: data <= 15'h7ff9; 
        10'b0101010011: data <= 15'h7ffa; 
        10'b0101010100: data <= 15'h7fe1; 
        10'b0101010101: data <= 15'h0005; 
        10'b0101010110: data <= 15'h002e; 
        10'b0101010111: data <= 15'h0030; 
        10'b0101011000: data <= 15'h0017; 
        10'b0101011001: data <= 15'h7ffa; 
        10'b0101011010: data <= 15'h0021; 
        10'b0101011011: data <= 15'h0017; 
        10'b0101011100: data <= 15'h002b; 
        10'b0101011101: data <= 15'h7fdd; 
        10'b0101011110: data <= 15'h7f18; 
        10'b0101011111: data <= 15'h7ee1; 
        10'b0101100000: data <= 15'h7ee2; 
        10'b0101100001: data <= 15'h7f64; 
        10'b0101100010: data <= 15'h7fe4; 
        10'b0101100011: data <= 15'h7ff5; 
        10'b0101100100: data <= 15'h000e; 
        10'b0101100101: data <= 15'h0028; 
        10'b0101100110: data <= 15'h0098; 
        10'b0101100111: data <= 15'h008b; 
        10'b0101101000: data <= 15'h0061; 
        10'b0101101001: data <= 15'h0003; 
        10'b0101101010: data <= 15'h7ff1; 
        10'b0101101011: data <= 15'h7ff1; 
        10'b0101101100: data <= 15'h7fe9; 
        10'b0101101101: data <= 15'h7fff; 
        10'b0101101110: data <= 15'h0008; 
        10'b0101101111: data <= 15'h7fea; 
        10'b0101110000: data <= 15'h7ff8; 
        10'b0101110001: data <= 15'h001c; 
        10'b0101110010: data <= 15'h0038; 
        10'b0101110011: data <= 15'h0048; 
        10'b0101110100: data <= 15'h0036; 
        10'b0101110101: data <= 15'h0026; 
        10'b0101110110: data <= 15'h0034; 
        10'b0101110111: data <= 15'h0028; 
        10'b0101111000: data <= 15'h001d; 
        10'b0101111001: data <= 15'h7f73; 
        10'b0101111010: data <= 15'h7f18; 
        10'b0101111011: data <= 15'h7ed9; 
        10'b0101111100: data <= 15'h7f0e; 
        10'b0101111101: data <= 15'h7f88; 
        10'b0101111110: data <= 15'h7fc5; 
        10'b0101111111: data <= 15'h7fb1; 
        10'b0110000000: data <= 15'h7fc4; 
        10'b0110000001: data <= 15'h001a; 
        10'b0110000010: data <= 15'h0064; 
        10'b0110000011: data <= 15'h009d; 
        10'b0110000100: data <= 15'h0059; 
        10'b0110000101: data <= 15'h000e; 
        10'b0110000110: data <= 15'h0000; 
        10'b0110000111: data <= 15'h0009; 
        10'b0110001000: data <= 15'h7ffd; 
        10'b0110001001: data <= 15'h0007; 
        10'b0110001010: data <= 15'h7fef; 
        10'b0110001011: data <= 15'h7ff3; 
        10'b0110001100: data <= 15'h7fe5; 
        10'b0110001101: data <= 15'h0049; 
        10'b0110001110: data <= 15'h005f; 
        10'b0110001111: data <= 15'h0074; 
        10'b0110010000: data <= 15'h0038; 
        10'b0110010001: data <= 15'h0043; 
        10'b0110010010: data <= 15'h0062; 
        10'b0110010011: data <= 15'h0038; 
        10'b0110010100: data <= 15'h000e; 
        10'b0110010101: data <= 15'h7f85; 
        10'b0110010110: data <= 15'h7eee; 
        10'b0110010111: data <= 15'h7ed8; 
        10'b0110011000: data <= 15'h7f15; 
        10'b0110011001: data <= 15'h7f7f; 
        10'b0110011010: data <= 15'h7fc7; 
        10'b0110011011: data <= 15'h7fbb; 
        10'b0110011100: data <= 15'h0006; 
        10'b0110011101: data <= 15'h0038; 
        10'b0110011110: data <= 15'h0043; 
        10'b0110011111: data <= 15'h009e; 
        10'b0110100000: data <= 15'h0052; 
        10'b0110100001: data <= 15'h7fef; 
        10'b0110100010: data <= 15'h7ff8; 
        10'b0110100011: data <= 15'h7fee; 
        10'b0110100100: data <= 15'h0009; 
        10'b0110100101: data <= 15'h0005; 
        10'b0110100110: data <= 15'h7ff1; 
        10'b0110100111: data <= 15'h7ffd; 
        10'b0110101000: data <= 15'h7fff; 
        10'b0110101001: data <= 15'h0068; 
        10'b0110101010: data <= 15'h004b; 
        10'b0110101011: data <= 15'h0067; 
        10'b0110101100: data <= 15'h0047; 
        10'b0110101101: data <= 15'h005f; 
        10'b0110101110: data <= 15'h0078; 
        10'b0110101111: data <= 15'h0021; 
        10'b0110110000: data <= 15'h7fa6; 
        10'b0110110001: data <= 15'h7f1a; 
        10'b0110110010: data <= 15'h7ecd; 
        10'b0110110011: data <= 15'h7edc; 
        10'b0110110100: data <= 15'h7f3b; 
        10'b0110110101: data <= 15'h7fa0; 
        10'b0110110110: data <= 15'h7fdc; 
        10'b0110110111: data <= 15'h7fdd; 
        10'b0110111000: data <= 15'h001e; 
        10'b0110111001: data <= 15'h001a; 
        10'b0110111010: data <= 15'h0065; 
        10'b0110111011: data <= 15'h0076; 
        10'b0110111100: data <= 15'h003d; 
        10'b0110111101: data <= 15'h7ffa; 
        10'b0110111110: data <= 15'h0002; 
        10'b0110111111: data <= 15'h7ff0; 
        10'b0111000000: data <= 15'h0003; 
        10'b0111000001: data <= 15'h000c; 
        10'b0111000010: data <= 15'h7fe9; 
        10'b0111000011: data <= 15'h7ff3; 
        10'b0111000100: data <= 15'h0011; 
        10'b0111000101: data <= 15'h005e; 
        10'b0111000110: data <= 15'h0075; 
        10'b0111000111: data <= 15'h005a; 
        10'b0111001000: data <= 15'h003f; 
        10'b0111001001: data <= 15'h003f; 
        10'b0111001010: data <= 15'h006b; 
        10'b0111001011: data <= 15'h7ff2; 
        10'b0111001100: data <= 15'h7f51; 
        10'b0111001101: data <= 15'h7ecf; 
        10'b0111001110: data <= 15'h7ed7; 
        10'b0111001111: data <= 15'h7f15; 
        10'b0111010000: data <= 15'h7f82; 
        10'b0111010001: data <= 15'h7fc5; 
        10'b0111010010: data <= 15'h7fff; 
        10'b0111010011: data <= 15'h0013; 
        10'b0111010100: data <= 15'h002c; 
        10'b0111010101: data <= 15'h0042; 
        10'b0111010110: data <= 15'h005b; 
        10'b0111010111: data <= 15'h0057; 
        10'b0111011000: data <= 15'h0021; 
        10'b0111011001: data <= 15'h0002; 
        10'b0111011010: data <= 15'h7ff5; 
        10'b0111011011: data <= 15'h7ff2; 
        10'b0111011100: data <= 15'h7ff8; 
        10'b0111011101: data <= 15'h0003; 
        10'b0111011110: data <= 15'h7fec; 
        10'b0111011111: data <= 15'h7fd9; 
        10'b0111100000: data <= 15'h0003; 
        10'b0111100001: data <= 15'h0043; 
        10'b0111100010: data <= 15'h0054; 
        10'b0111100011: data <= 15'h0051; 
        10'b0111100100: data <= 15'h0019; 
        10'b0111100101: data <= 15'h0041; 
        10'b0111100110: data <= 15'h0067; 
        10'b0111100111: data <= 15'h7ff0; 
        10'b0111101000: data <= 15'h7f2e; 
        10'b0111101001: data <= 15'h7ed4; 
        10'b0111101010: data <= 15'h7ef8; 
        10'b0111101011: data <= 15'h7f62; 
        10'b0111101100: data <= 15'h7feb; 
        10'b0111101101: data <= 15'h0028; 
        10'b0111101110: data <= 15'h003a; 
        10'b0111101111: data <= 15'h0035; 
        10'b0111110000: data <= 15'h0044; 
        10'b0111110001: data <= 15'h0034; 
        10'b0111110010: data <= 15'h0029; 
        10'b0111110011: data <= 15'h002f; 
        10'b0111110100: data <= 15'h7ffd; 
        10'b0111110101: data <= 15'h7ff9; 
        10'b0111110110: data <= 15'h0004; 
        10'b0111110111: data <= 15'h7ff0; 
        10'b0111111000: data <= 15'h7ff5; 
        10'b0111111001: data <= 15'h0004; 
        10'b0111111010: data <= 15'h7ff8; 
        10'b0111111011: data <= 15'h7ff1; 
        10'b0111111100: data <= 15'h7ff8; 
        10'b0111111101: data <= 15'h002b; 
        10'b0111111110: data <= 15'h0057; 
        10'b0111111111: data <= 15'h0032; 
        10'b1000000000: data <= 15'h001f; 
        10'b1000000001: data <= 15'h0056; 
        10'b1000000010: data <= 15'h00a6; 
        10'b1000000011: data <= 15'h0007; 
        10'b1000000100: data <= 15'h7f7a; 
        10'b1000000101: data <= 15'h7f28; 
        10'b1000000110: data <= 15'h7f6a; 
        10'b1000000111: data <= 15'h7fd2; 
        10'b1000001000: data <= 15'h0031; 
        10'b1000001001: data <= 15'h0034; 
        10'b1000001010: data <= 15'h0036; 
        10'b1000001011: data <= 15'h001c; 
        10'b1000001100: data <= 15'h000e; 
        10'b1000001101: data <= 15'h0017; 
        10'b1000001110: data <= 15'h002d; 
        10'b1000001111: data <= 15'h001c; 
        10'b1000010000: data <= 15'h7ffd; 
        10'b1000010001: data <= 15'h7ff2; 
        10'b1000010010: data <= 15'h0002; 
        10'b1000010011: data <= 15'h7ff8; 
        10'b1000010100: data <= 15'h7ff9; 
        10'b1000010101: data <= 15'h7ff6; 
        10'b1000010110: data <= 15'h7ff7; 
        10'b1000010111: data <= 15'h7fda; 
        10'b1000011000: data <= 15'h0010; 
        10'b1000011001: data <= 15'h002f; 
        10'b1000011010: data <= 15'h0070; 
        10'b1000011011: data <= 15'h0065; 
        10'b1000011100: data <= 15'h004f; 
        10'b1000011101: data <= 15'h0069; 
        10'b1000011110: data <= 15'h00a6; 
        10'b1000011111: data <= 15'h0075; 
        10'b1000100000: data <= 15'h0019; 
        10'b1000100001: data <= 15'h7fca; 
        10'b1000100010: data <= 15'h7fe9; 
        10'b1000100011: data <= 15'h7ff1; 
        10'b1000100100: data <= 15'h0019; 
        10'b1000100101: data <= 15'h7ff4; 
        10'b1000100110: data <= 15'h7fea; 
        10'b1000100111: data <= 15'h7ff3; 
        10'b1000101000: data <= 15'h001a; 
        10'b1000101001: data <= 15'h0018; 
        10'b1000101010: data <= 15'h002f; 
        10'b1000101011: data <= 15'h7ffa; 
        10'b1000101100: data <= 15'h0007; 
        10'b1000101101: data <= 15'h7ff6; 
        10'b1000101110: data <= 15'h7fe8; 
        10'b1000101111: data <= 15'h0008; 
        10'b1000110000: data <= 15'h0008; 
        10'b1000110001: data <= 15'h000b; 
        10'b1000110010: data <= 15'h7ff8; 
        10'b1000110011: data <= 15'h7fee; 
        10'b1000110100: data <= 15'h7ff5; 
        10'b1000110101: data <= 15'h0030; 
        10'b1000110110: data <= 15'h005a; 
        10'b1000110111: data <= 15'h0042; 
        10'b1000111000: data <= 15'h0052; 
        10'b1000111001: data <= 15'h0065; 
        10'b1000111010: data <= 15'h009d; 
        10'b1000111011: data <= 15'h009d; 
        10'b1000111100: data <= 15'h004e; 
        10'b1000111101: data <= 15'h0018; 
        10'b1000111110: data <= 15'h7ff0; 
        10'b1000111111: data <= 15'h000b; 
        10'b1001000000: data <= 15'h000b; 
        10'b1001000001: data <= 15'h7fe9; 
        10'b1001000010: data <= 15'h7fef; 
        10'b1001000011: data <= 15'h7fe8; 
        10'b1001000100: data <= 15'h000d; 
        10'b1001000101: data <= 15'h0010; 
        10'b1001000110: data <= 15'h0019; 
        10'b1001000111: data <= 15'h0009; 
        10'b1001001000: data <= 15'h7ff2; 
        10'b1001001001: data <= 15'h7ffd; 
        10'b1001001010: data <= 15'h7fed; 
        10'b1001001011: data <= 15'h7ff6; 
        10'b1001001100: data <= 15'h7ff2; 
        10'b1001001101: data <= 15'h7feb; 
        10'b1001001110: data <= 15'h7ff8; 
        10'b1001001111: data <= 15'h7ff2; 
        10'b1001010000: data <= 15'h7ff7; 
        10'b1001010001: data <= 15'h000c; 
        10'b1001010010: data <= 15'h0037; 
        10'b1001010011: data <= 15'h005a; 
        10'b1001010100: data <= 15'h003f; 
        10'b1001010101: data <= 15'h0045; 
        10'b1001010110: data <= 15'h0086; 
        10'b1001010111: data <= 15'h0098; 
        10'b1001011000: data <= 15'h0065; 
        10'b1001011001: data <= 15'h0026; 
        10'b1001011010: data <= 15'h000e; 
        10'b1001011011: data <= 15'h0003; 
        10'b1001011100: data <= 15'h7ffe; 
        10'b1001011101: data <= 15'h7fd6; 
        10'b1001011110: data <= 15'h7fe0; 
        10'b1001011111: data <= 15'h7fee; 
        10'b1001100000: data <= 15'h0010; 
        10'b1001100001: data <= 15'h7fff; 
        10'b1001100010: data <= 15'h7fed; 
        10'b1001100011: data <= 15'h7fe2; 
        10'b1001100100: data <= 15'h7ff9; 
        10'b1001100101: data <= 15'h7ff6; 
        10'b1001100110: data <= 15'h7ff1; 
        10'b1001100111: data <= 15'h7ff3; 
        10'b1001101000: data <= 15'h7fee; 
        10'b1001101001: data <= 15'h0001; 
        10'b1001101010: data <= 15'h0002; 
        10'b1001101011: data <= 15'h7ff5; 
        10'b1001101100: data <= 15'h7fed; 
        10'b1001101101: data <= 15'h0007; 
        10'b1001101110: data <= 15'h0028; 
        10'b1001101111: data <= 15'h0023; 
        10'b1001110000: data <= 15'h0065; 
        10'b1001110001: data <= 15'h0052; 
        10'b1001110010: data <= 15'h005b; 
        10'b1001110011: data <= 15'h006c; 
        10'b1001110100: data <= 15'h005c; 
        10'b1001110101: data <= 15'h0076; 
        10'b1001110110: data <= 15'h0033; 
        10'b1001110111: data <= 15'h0034; 
        10'b1001111000: data <= 15'h001d; 
        10'b1001111001: data <= 15'h7fe8; 
        10'b1001111010: data <= 15'h7fed; 
        10'b1001111011: data <= 15'h7fff; 
        10'b1001111100: data <= 15'h7fe5; 
        10'b1001111101: data <= 15'h7fe3; 
        10'b1001111110: data <= 15'h7ff2; 
        10'b1001111111: data <= 15'h7ff1; 
        10'b1010000000: data <= 15'h7ffb; 
        10'b1010000001: data <= 15'h7ff7; 
        10'b1010000010: data <= 15'h7ff4; 
        10'b1010000011: data <= 15'h7ffa; 
        10'b1010000100: data <= 15'h7fee; 
        10'b1010000101: data <= 15'h7ffb; 
        10'b1010000110: data <= 15'h0000; 
        10'b1010000111: data <= 15'h7fea; 
        10'b1010001000: data <= 15'h7fea; 
        10'b1010001001: data <= 15'h7ffa; 
        10'b1010001010: data <= 15'h7ffd; 
        10'b1010001011: data <= 15'h001c; 
        10'b1010001100: data <= 15'h0028; 
        10'b1010001101: data <= 15'h005e; 
        10'b1010001110: data <= 15'h0070; 
        10'b1010001111: data <= 15'h0089; 
        10'b1010010000: data <= 15'h0088; 
        10'b1010010001: data <= 15'h0051; 
        10'b1010010010: data <= 15'h0042; 
        10'b1010010011: data <= 15'h0025; 
        10'b1010010100: data <= 15'h000f; 
        10'b1010010101: data <= 15'h7ffe; 
        10'b1010010110: data <= 15'h7fcc; 
        10'b1010010111: data <= 15'h7fbf; 
        10'b1010011000: data <= 15'h7fce; 
        10'b1010011001: data <= 15'h7fe7; 
        10'b1010011010: data <= 15'h7fec; 
        10'b1010011011: data <= 15'h7ffd; 
        10'b1010011100: data <= 15'h7ff8; 
        10'b1010011101: data <= 15'h0006; 
        10'b1010011110: data <= 15'h7ff5; 
        10'b1010011111: data <= 15'h7fe9; 
        10'b1010100000: data <= 15'h7ff6; 
        10'b1010100001: data <= 15'h7ffc; 
        10'b1010100010: data <= 15'h7fea; 
        10'b1010100011: data <= 15'h7fff; 
        10'b1010100100: data <= 15'h7ffa; 
        10'b1010100101: data <= 15'h7ffa; 
        10'b1010100110: data <= 15'h7fe5; 
        10'b1010100111: data <= 15'h7fdc; 
        10'b1010101000: data <= 15'h7fec; 
        10'b1010101001: data <= 15'h7fee; 
        10'b1010101010: data <= 15'h0015; 
        10'b1010101011: data <= 15'h0010; 
        10'b1010101100: data <= 15'h0026; 
        10'b1010101101: data <= 15'h0037; 
        10'b1010101110: data <= 15'h001d; 
        10'b1010101111: data <= 15'h7fea; 
        10'b1010110000: data <= 15'h7fdd; 
        10'b1010110001: data <= 15'h7fd7; 
        10'b1010110010: data <= 15'h7fdd; 
        10'b1010110011: data <= 15'h7fcf; 
        10'b1010110100: data <= 15'h7fd1; 
        10'b1010110101: data <= 15'h7fd4; 
        10'b1010110110: data <= 15'h7ff7; 
        10'b1010110111: data <= 15'h7ff4; 
        10'b1010111000: data <= 15'h7fed; 
        10'b1010111001: data <= 15'h7ff2; 
        10'b1010111010: data <= 15'h0001; 
        10'b1010111011: data <= 15'h7ff0; 
        10'b1010111100: data <= 15'h7ff2; 
        10'b1010111101: data <= 15'h000d; 
        10'b1010111110: data <= 15'h7ff9; 
        10'b1010111111: data <= 15'h000b; 
        10'b1011000000: data <= 15'h000c; 
        10'b1011000001: data <= 15'h7fff; 
        10'b1011000010: data <= 15'h7fe8; 
        10'b1011000011: data <= 15'h7ff5; 
        10'b1011000100: data <= 15'h7fd1; 
        10'b1011000101: data <= 15'h7fd4; 
        10'b1011000110: data <= 15'h7fc9; 
        10'b1011000111: data <= 15'h7fb8; 
        10'b1011001000: data <= 15'h7fae; 
        10'b1011001001: data <= 15'h7fb5; 
        10'b1011001010: data <= 15'h7fa9; 
        10'b1011001011: data <= 15'h7fb2; 
        10'b1011001100: data <= 15'h7fb6; 
        10'b1011001101: data <= 15'h7fd3; 
        10'b1011001110: data <= 15'h7fdb; 
        10'b1011001111: data <= 15'h7fe1; 
        10'b1011010000: data <= 15'h7fdd; 
        10'b1011010001: data <= 15'h7fe0; 
        10'b1011010010: data <= 15'h7ff5; 
        10'b1011010011: data <= 15'h000c; 
        10'b1011010100: data <= 15'h0006; 
        10'b1011010101: data <= 15'h7ff7; 
        10'b1011010110: data <= 15'h7ff5; 
        10'b1011010111: data <= 15'h7ffc; 
        10'b1011011000: data <= 15'h000a; 
        10'b1011011001: data <= 15'h0009; 
        10'b1011011010: data <= 15'h7ff7; 
        10'b1011011011: data <= 15'h0001; 
        10'b1011011100: data <= 15'h7ff3; 
        10'b1011011101: data <= 15'h7ff6; 
        10'b1011011110: data <= 15'h7fea; 
        10'b1011011111: data <= 15'h0004; 
        10'b1011100000: data <= 15'h7ff4; 
        10'b1011100001: data <= 15'h7fd9; 
        10'b1011100010: data <= 15'h7fd9; 
        10'b1011100011: data <= 15'h7fdc; 
        10'b1011100100: data <= 15'h7ff2; 
        10'b1011100101: data <= 15'h7fdc; 
        10'b1011100110: data <= 15'h7fde; 
        10'b1011100111: data <= 15'h7ff3; 
        10'b1011101000: data <= 15'h7fdc; 
        10'b1011101001: data <= 15'h7fe3; 
        10'b1011101010: data <= 15'h7fea; 
        10'b1011101011: data <= 15'h7fe5; 
        10'b1011101100: data <= 15'h7ff2; 
        10'b1011101101: data <= 15'h7fdf; 
        10'b1011101110: data <= 15'h7fe4; 
        10'b1011101111: data <= 15'h000b; 
        10'b1011110000: data <= 15'h7fef; 
        10'b1011110001: data <= 15'h0003; 
        10'b1011110010: data <= 15'h0009; 
        10'b1011110011: data <= 15'h7ffe; 
        10'b1011110100: data <= 15'h7fed; 
        10'b1011110101: data <= 15'h0007; 
        10'b1011110110: data <= 15'h7ffd; 
        10'b1011110111: data <= 15'h7ff6; 
        10'b1011111000: data <= 15'h000a; 
        10'b1011111001: data <= 15'h0002; 
        10'b1011111010: data <= 15'h0003; 
        10'b1011111011: data <= 15'h7fe9; 
        10'b1011111100: data <= 15'h000b; 
        10'b1011111101: data <= 15'h000b; 
        10'b1011111110: data <= 15'h0004; 
        10'b1011111111: data <= 15'h0008; 
        10'b1100000000: data <= 15'h7ffb; 
        10'b1100000001: data <= 15'h7ff3; 
        10'b1100000010: data <= 15'h0007; 
        10'b1100000011: data <= 15'h7fec; 
        10'b1100000100: data <= 15'h7ff9; 
        10'b1100000101: data <= 15'h7ff2; 
        10'b1100000110: data <= 15'h7ffd; 
        10'b1100000111: data <= 15'h7ff4; 
        10'b1100001000: data <= 15'h7fe9; 
        10'b1100001001: data <= 15'h7feb; 
        10'b1100001010: data <= 15'h7fe2; 
        10'b1100001011: data <= 15'h7ff9; 
        10'b1100001100: data <= 15'h0005; 
        10'b1100001101: data <= 15'h7fed; 
        10'b1100001110: data <= 15'h7fe8; 
        10'b1100001111: data <= 15'h0006; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 10) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 16'hffdf; 
        10'b0000000001: data <= 16'h0013; 
        10'b0000000010: data <= 16'hfff6; 
        10'b0000000011: data <= 16'hfffb; 
        10'b0000000100: data <= 16'h0016; 
        10'b0000000101: data <= 16'hfffe; 
        10'b0000000110: data <= 16'hffeb; 
        10'b0000000111: data <= 16'hffea; 
        10'b0000001000: data <= 16'hfffb; 
        10'b0000001001: data <= 16'hfff5; 
        10'b0000001010: data <= 16'h0019; 
        10'b0000001011: data <= 16'hfffe; 
        10'b0000001100: data <= 16'h000b; 
        10'b0000001101: data <= 16'hffe0; 
        10'b0000001110: data <= 16'hfffe; 
        10'b0000001111: data <= 16'hffd4; 
        10'b0000010000: data <= 16'hffdb; 
        10'b0000010001: data <= 16'hfff6; 
        10'b0000010010: data <= 16'hffda; 
        10'b0000010011: data <= 16'h0019; 
        10'b0000010100: data <= 16'hffdb; 
        10'b0000010101: data <= 16'hfff4; 
        10'b0000010110: data <= 16'hffd8; 
        10'b0000010111: data <= 16'hfffc; 
        10'b0000011000: data <= 16'h000c; 
        10'b0000011001: data <= 16'hfff7; 
        10'b0000011010: data <= 16'hfffe; 
        10'b0000011011: data <= 16'hffff; 
        10'b0000011100: data <= 16'h000e; 
        10'b0000011101: data <= 16'h0011; 
        10'b0000011110: data <= 16'h0006; 
        10'b0000011111: data <= 16'hffd9; 
        10'b0000100000: data <= 16'hffd7; 
        10'b0000100001: data <= 16'h0002; 
        10'b0000100010: data <= 16'hffe0; 
        10'b0000100011: data <= 16'hfff7; 
        10'b0000100100: data <= 16'hffe7; 
        10'b0000100101: data <= 16'hffd2; 
        10'b0000100110: data <= 16'hffe3; 
        10'b0000100111: data <= 16'h0002; 
        10'b0000101000: data <= 16'h001c; 
        10'b0000101001: data <= 16'hffda; 
        10'b0000101010: data <= 16'hffeb; 
        10'b0000101011: data <= 16'h000c; 
        10'b0000101100: data <= 16'hffe0; 
        10'b0000101101: data <= 16'hffd5; 
        10'b0000101110: data <= 16'h0008; 
        10'b0000101111: data <= 16'h0013; 
        10'b0000110000: data <= 16'hffdf; 
        10'b0000110001: data <= 16'h0009; 
        10'b0000110010: data <= 16'hffe4; 
        10'b0000110011: data <= 16'hffdc; 
        10'b0000110100: data <= 16'hfff9; 
        10'b0000110101: data <= 16'h0002; 
        10'b0000110110: data <= 16'hfff5; 
        10'b0000110111: data <= 16'h0018; 
        10'b0000111000: data <= 16'hffd7; 
        10'b0000111001: data <= 16'hffe7; 
        10'b0000111010: data <= 16'hffe4; 
        10'b0000111011: data <= 16'h000c; 
        10'b0000111100: data <= 16'h0003; 
        10'b0000111101: data <= 16'hffd5; 
        10'b0000111110: data <= 16'hfff6; 
        10'b0000111111: data <= 16'h0017; 
        10'b0001000000: data <= 16'hfff2; 
        10'b0001000001: data <= 16'hffe1; 
        10'b0001000010: data <= 16'hffe2; 
        10'b0001000011: data <= 16'hffcd; 
        10'b0001000100: data <= 16'hffca; 
        10'b0001000101: data <= 16'hffed; 
        10'b0001000110: data <= 16'hffc8; 
        10'b0001000111: data <= 16'hffb8; 
        10'b0001001000: data <= 16'hffcc; 
        10'b0001001001: data <= 16'hfff2; 
        10'b0001001010: data <= 16'hffd4; 
        10'b0001001011: data <= 16'hffc7; 
        10'b0001001100: data <= 16'hfff6; 
        10'b0001001101: data <= 16'h0011; 
        10'b0001001110: data <= 16'h0003; 
        10'b0001001111: data <= 16'hffe0; 
        10'b0001010000: data <= 16'h0016; 
        10'b0001010001: data <= 16'hffd2; 
        10'b0001010010: data <= 16'hfff5; 
        10'b0001010011: data <= 16'h000a; 
        10'b0001010100: data <= 16'hffd5; 
        10'b0001010101: data <= 16'hfff6; 
        10'b0001010110: data <= 16'h0018; 
        10'b0001010111: data <= 16'hffd7; 
        10'b0001011000: data <= 16'hffe2; 
        10'b0001011001: data <= 16'h0013; 
        10'b0001011010: data <= 16'h0008; 
        10'b0001011011: data <= 16'h0001; 
        10'b0001011100: data <= 16'h0003; 
        10'b0001011101: data <= 16'hfff5; 
        10'b0001011110: data <= 16'hfff2; 
        10'b0001011111: data <= 16'hffc8; 
        10'b0001100000: data <= 16'hffb3; 
        10'b0001100001: data <= 16'hffd4; 
        10'b0001100010: data <= 16'hffc4; 
        10'b0001100011: data <= 16'hffbc; 
        10'b0001100100: data <= 16'h000b; 
        10'b0001100101: data <= 16'h0005; 
        10'b0001100110: data <= 16'hffb4; 
        10'b0001100111: data <= 16'hffbf; 
        10'b0001101000: data <= 16'hffa3; 
        10'b0001101001: data <= 16'hffbe; 
        10'b0001101010: data <= 16'hffb0; 
        10'b0001101011: data <= 16'hffc8; 
        10'b0001101100: data <= 16'hffd9; 
        10'b0001101101: data <= 16'h000f; 
        10'b0001101110: data <= 16'h000e; 
        10'b0001101111: data <= 16'hffea; 
        10'b0001110000: data <= 16'h0006; 
        10'b0001110001: data <= 16'hffd5; 
        10'b0001110010: data <= 16'hffe2; 
        10'b0001110011: data <= 16'hffd6; 
        10'b0001110100: data <= 16'hffd0; 
        10'b0001110101: data <= 16'hfffa; 
        10'b0001110110: data <= 16'hfff3; 
        10'b0001110111: data <= 16'hffd5; 
        10'b0001111000: data <= 16'hfff2; 
        10'b0001111001: data <= 16'hfff7; 
        10'b0001111010: data <= 16'hffbb; 
        10'b0001111011: data <= 16'hffbc; 
        10'b0001111100: data <= 16'hffbd; 
        10'b0001111101: data <= 16'hffc0; 
        10'b0001111110: data <= 16'hffee; 
        10'b0001111111: data <= 16'hfff9; 
        10'b0010000000: data <= 16'hffcb; 
        10'b0010000001: data <= 16'hffce; 
        10'b0010000010: data <= 16'hffcd; 
        10'b0010000011: data <= 16'hffb8; 
        10'b0010000100: data <= 16'hffe3; 
        10'b0010000101: data <= 16'hffa4; 
        10'b0010000110: data <= 16'hffdc; 
        10'b0010000111: data <= 16'hfffb; 
        10'b0010001000: data <= 16'hffd8; 
        10'b0010001001: data <= 16'hffee; 
        10'b0010001010: data <= 16'hffe8; 
        10'b0010001011: data <= 16'hfffc; 
        10'b0010001100: data <= 16'h000b; 
        10'b0010001101: data <= 16'hffec; 
        10'b0010001110: data <= 16'hffff; 
        10'b0010001111: data <= 16'hffda; 
        10'b0010010000: data <= 16'hfff6; 
        10'b0010010001: data <= 16'hffee; 
        10'b0010010010: data <= 16'hfff2; 
        10'b0010010011: data <= 16'hffe3; 
        10'b0010010100: data <= 16'hfff3; 
        10'b0010010101: data <= 16'hffcc; 
        10'b0010010110: data <= 16'hffe9; 
        10'b0010010111: data <= 16'h000f; 
        10'b0010011000: data <= 16'h003c; 
        10'b0010011001: data <= 16'h0083; 
        10'b0010011010: data <= 16'h009e; 
        10'b0010011011: data <= 16'h009c; 
        10'b0010011100: data <= 16'h00b0; 
        10'b0010011101: data <= 16'h00bd; 
        10'b0010011110: data <= 16'h00c8; 
        10'b0010011111: data <= 16'h0046; 
        10'b0010100000: data <= 16'h000d; 
        10'b0010100001: data <= 16'h0021; 
        10'b0010100010: data <= 16'hfff0; 
        10'b0010100011: data <= 16'hfffe; 
        10'b0010100100: data <= 16'hffab; 
        10'b0010100101: data <= 16'hffc2; 
        10'b0010100110: data <= 16'hfffc; 
        10'b0010100111: data <= 16'hffdf; 
        10'b0010101000: data <= 16'hffef; 
        10'b0010101001: data <= 16'hfff8; 
        10'b0010101010: data <= 16'h0005; 
        10'b0010101011: data <= 16'hfff2; 
        10'b0010101100: data <= 16'h0001; 
        10'b0010101101: data <= 16'h0002; 
        10'b0010101110: data <= 16'h0005; 
        10'b0010101111: data <= 16'hfffe; 
        10'b0010110000: data <= 16'hffd5; 
        10'b0010110001: data <= 16'hffb7; 
        10'b0010110010: data <= 16'h0028; 
        10'b0010110011: data <= 16'hfffa; 
        10'b0010110100: data <= 16'h006c; 
        10'b0010110101: data <= 16'h0060; 
        10'b0010110110: data <= 16'h005b; 
        10'b0010110111: data <= 16'h0088; 
        10'b0010111000: data <= 16'h00a6; 
        10'b0010111001: data <= 16'h00eb; 
        10'b0010111010: data <= 16'h00da; 
        10'b0010111011: data <= 16'h00ba; 
        10'b0010111100: data <= 16'h00b3; 
        10'b0010111101: data <= 16'h00cd; 
        10'b0010111110: data <= 16'h0074; 
        10'b0010111111: data <= 16'h002a; 
        10'b0011000000: data <= 16'hffa7; 
        10'b0011000001: data <= 16'hffa3; 
        10'b0011000010: data <= 16'hffc1; 
        10'b0011000011: data <= 16'h0009; 
        10'b0011000100: data <= 16'h0015; 
        10'b0011000101: data <= 16'h0003; 
        10'b0011000110: data <= 16'hfffc; 
        10'b0011000111: data <= 16'hffc9; 
        10'b0011001000: data <= 16'hffab; 
        10'b0011001001: data <= 16'hfff9; 
        10'b0011001010: data <= 16'hffde; 
        10'b0011001011: data <= 16'h0001; 
        10'b0011001100: data <= 16'hffd8; 
        10'b0011001101: data <= 16'hfff4; 
        10'b0011001110: data <= 16'h0008; 
        10'b0011001111: data <= 16'h004d; 
        10'b0011010000: data <= 16'h00a1; 
        10'b0011010001: data <= 16'h0094; 
        10'b0011010010: data <= 16'h003d; 
        10'b0011010011: data <= 16'h005f; 
        10'b0011010100: data <= 16'h0087; 
        10'b0011010101: data <= 16'h00fc; 
        10'b0011010110: data <= 16'h00b9; 
        10'b0011010111: data <= 16'h00a2; 
        10'b0011011000: data <= 16'h0042; 
        10'b0011011001: data <= 16'h007f; 
        10'b0011011010: data <= 16'h008c; 
        10'b0011011011: data <= 16'h0048; 
        10'b0011011100: data <= 16'hffca; 
        10'b0011011101: data <= 16'hffa7; 
        10'b0011011110: data <= 16'hffb0; 
        10'b0011011111: data <= 16'hfffb; 
        10'b0011100000: data <= 16'h0018; 
        10'b0011100001: data <= 16'h0009; 
        10'b0011100010: data <= 16'hfff6; 
        10'b0011100011: data <= 16'h0000; 
        10'b0011100100: data <= 16'hffc2; 
        10'b0011100101: data <= 16'hffd0; 
        10'b0011100110: data <= 16'hffd8; 
        10'b0011100111: data <= 16'hffcf; 
        10'b0011101000: data <= 16'hffe6; 
        10'b0011101001: data <= 16'hffe5; 
        10'b0011101010: data <= 16'h004c; 
        10'b0011101011: data <= 16'h0050; 
        10'b0011101100: data <= 16'h0029; 
        10'b0011101101: data <= 16'h0011; 
        10'b0011101110: data <= 16'h001d; 
        10'b0011101111: data <= 16'h0071; 
        10'b0011110000: data <= 16'h014a; 
        10'b0011110001: data <= 16'h0107; 
        10'b0011110010: data <= 16'h00f4; 
        10'b0011110011: data <= 16'h004d; 
        10'b0011110100: data <= 16'h0041; 
        10'b0011110101: data <= 16'h003b; 
        10'b0011110110: data <= 16'h0091; 
        10'b0011110111: data <= 16'h00fc; 
        10'b0011111000: data <= 16'hffe4; 
        10'b0011111001: data <= 16'hffac; 
        10'b0011111010: data <= 16'hfff8; 
        10'b0011111011: data <= 16'hffd4; 
        10'b0011111100: data <= 16'hfff9; 
        10'b0011111101: data <= 16'hfffc; 
        10'b0011111110: data <= 16'h0007; 
        10'b0011111111: data <= 16'h0006; 
        10'b0100000000: data <= 16'hffb2; 
        10'b0100000001: data <= 16'hffc8; 
        10'b0100000010: data <= 16'hffb0; 
        10'b0100000011: data <= 16'hffd2; 
        10'b0100000100: data <= 16'hffd3; 
        10'b0100000101: data <= 16'hffe9; 
        10'b0100000110: data <= 16'h0037; 
        10'b0100000111: data <= 16'hffd1; 
        10'b0100001000: data <= 16'h001b; 
        10'b0100001001: data <= 16'h0053; 
        10'b0100001010: data <= 16'h004a; 
        10'b0100001011: data <= 16'h003f; 
        10'b0100001100: data <= 16'h00b5; 
        10'b0100001101: data <= 16'h00f1; 
        10'b0100001110: data <= 16'h0115; 
        10'b0100001111: data <= 16'h00a0; 
        10'b0100010000: data <= 16'h0031; 
        10'b0100010001: data <= 16'hfff7; 
        10'b0100010010: data <= 16'h0077; 
        10'b0100010011: data <= 16'h0101; 
        10'b0100010100: data <= 16'h004b; 
        10'b0100010101: data <= 16'hffc1; 
        10'b0100010110: data <= 16'h0001; 
        10'b0100010111: data <= 16'hfff8; 
        10'b0100011000: data <= 16'hffd7; 
        10'b0100011001: data <= 16'h0014; 
        10'b0100011010: data <= 16'hffde; 
        10'b0100011011: data <= 16'hffc2; 
        10'b0100011100: data <= 16'hffc7; 
        10'b0100011101: data <= 16'hffd3; 
        10'b0100011110: data <= 16'hffda; 
        10'b0100011111: data <= 16'h0005; 
        10'b0100100000: data <= 16'h001a; 
        10'b0100100001: data <= 16'hfffa; 
        10'b0100100010: data <= 16'hffd4; 
        10'b0100100011: data <= 16'h000e; 
        10'b0100100100: data <= 16'h0012; 
        10'b0100100101: data <= 16'hfff6; 
        10'b0100100110: data <= 16'hffa9; 
        10'b0100100111: data <= 16'hff6a; 
        10'b0100101000: data <= 16'hffa6; 
        10'b0100101001: data <= 16'h0057; 
        10'b0100101010: data <= 16'h00dd; 
        10'b0100101011: data <= 16'h00e5; 
        10'b0100101100: data <= 16'h00ca; 
        10'b0100101101: data <= 16'h0093; 
        10'b0100101110: data <= 16'h00d9; 
        10'b0100101111: data <= 16'h0129; 
        10'b0100110000: data <= 16'h008d; 
        10'b0100110001: data <= 16'hffc6; 
        10'b0100110010: data <= 16'hffc5; 
        10'b0100110011: data <= 16'hffd3; 
        10'b0100110100: data <= 16'hffe2; 
        10'b0100110101: data <= 16'hffd7; 
        10'b0100110110: data <= 16'h0011; 
        10'b0100110111: data <= 16'hfff3; 
        10'b0100111000: data <= 16'hff91; 
        10'b0100111001: data <= 16'hffe8; 
        10'b0100111010: data <= 16'h0011; 
        10'b0100111011: data <= 16'h0054; 
        10'b0100111100: data <= 16'h003f; 
        10'b0100111101: data <= 16'hffe8; 
        10'b0100111110: data <= 16'h0016; 
        10'b0100111111: data <= 16'h0002; 
        10'b0101000000: data <= 16'h002b; 
        10'b0101000001: data <= 16'hffe2; 
        10'b0101000010: data <= 16'hff14; 
        10'b0101000011: data <= 16'hfe4a; 
        10'b0101000100: data <= 16'hfe64; 
        10'b0101000101: data <= 16'hff5f; 
        10'b0101000110: data <= 16'hffeb; 
        10'b0101000111: data <= 16'h0074; 
        10'b0101001000: data <= 16'h00ba; 
        10'b0101001001: data <= 16'h00ac; 
        10'b0101001010: data <= 16'h00eb; 
        10'b0101001011: data <= 16'h010a; 
        10'b0101001100: data <= 16'h00c0; 
        10'b0101001101: data <= 16'hffdb; 
        10'b0101001110: data <= 16'hfffe; 
        10'b0101001111: data <= 16'hffd1; 
        10'b0101010000: data <= 16'hffe0; 
        10'b0101010001: data <= 16'hfff6; 
        10'b0101010010: data <= 16'hfff1; 
        10'b0101010011: data <= 16'hfff4; 
        10'b0101010100: data <= 16'hffc1; 
        10'b0101010101: data <= 16'h000a; 
        10'b0101010110: data <= 16'h005c; 
        10'b0101010111: data <= 16'h0060; 
        10'b0101011000: data <= 16'h002e; 
        10'b0101011001: data <= 16'hfff3; 
        10'b0101011010: data <= 16'h0042; 
        10'b0101011011: data <= 16'h002f; 
        10'b0101011100: data <= 16'h0056; 
        10'b0101011101: data <= 16'hffb9; 
        10'b0101011110: data <= 16'hfe30; 
        10'b0101011111: data <= 16'hfdc2; 
        10'b0101100000: data <= 16'hfdc4; 
        10'b0101100001: data <= 16'hfec7; 
        10'b0101100010: data <= 16'hffc9; 
        10'b0101100011: data <= 16'hffe9; 
        10'b0101100100: data <= 16'h001c; 
        10'b0101100101: data <= 16'h0050; 
        10'b0101100110: data <= 16'h0131; 
        10'b0101100111: data <= 16'h0117; 
        10'b0101101000: data <= 16'h00c2; 
        10'b0101101001: data <= 16'h0007; 
        10'b0101101010: data <= 16'hffe2; 
        10'b0101101011: data <= 16'hffe1; 
        10'b0101101100: data <= 16'hffd3; 
        10'b0101101101: data <= 16'hffff; 
        10'b0101101110: data <= 16'h0010; 
        10'b0101101111: data <= 16'hffd5; 
        10'b0101110000: data <= 16'hffef; 
        10'b0101110001: data <= 16'h0039; 
        10'b0101110010: data <= 16'h006f; 
        10'b0101110011: data <= 16'h008f; 
        10'b0101110100: data <= 16'h006c; 
        10'b0101110101: data <= 16'h004c; 
        10'b0101110110: data <= 16'h0068; 
        10'b0101110111: data <= 16'h0051; 
        10'b0101111000: data <= 16'h003a; 
        10'b0101111001: data <= 16'hfee6; 
        10'b0101111010: data <= 16'hfe30; 
        10'b0101111011: data <= 16'hfdb2; 
        10'b0101111100: data <= 16'hfe1b; 
        10'b0101111101: data <= 16'hff0f; 
        10'b0101111110: data <= 16'hff8a; 
        10'b0101111111: data <= 16'hff62; 
        10'b0110000000: data <= 16'hff87; 
        10'b0110000001: data <= 16'h0035; 
        10'b0110000010: data <= 16'h00c8; 
        10'b0110000011: data <= 16'h013a; 
        10'b0110000100: data <= 16'h00b2; 
        10'b0110000101: data <= 16'h001d; 
        10'b0110000110: data <= 16'h0000; 
        10'b0110000111: data <= 16'h0011; 
        10'b0110001000: data <= 16'hfffa; 
        10'b0110001001: data <= 16'h000e; 
        10'b0110001010: data <= 16'hffdd; 
        10'b0110001011: data <= 16'hffe7; 
        10'b0110001100: data <= 16'hffca; 
        10'b0110001101: data <= 16'h0093; 
        10'b0110001110: data <= 16'h00bf; 
        10'b0110001111: data <= 16'h00e7; 
        10'b0110010000: data <= 16'h006f; 
        10'b0110010001: data <= 16'h0085; 
        10'b0110010010: data <= 16'h00c4; 
        10'b0110010011: data <= 16'h0071; 
        10'b0110010100: data <= 16'h001c; 
        10'b0110010101: data <= 16'hff0a; 
        10'b0110010110: data <= 16'hfddc; 
        10'b0110010111: data <= 16'hfdb0; 
        10'b0110011000: data <= 16'hfe29; 
        10'b0110011001: data <= 16'hfefe; 
        10'b0110011010: data <= 16'hff8f; 
        10'b0110011011: data <= 16'hff77; 
        10'b0110011100: data <= 16'h000c; 
        10'b0110011101: data <= 16'h0070; 
        10'b0110011110: data <= 16'h0085; 
        10'b0110011111: data <= 16'h013d; 
        10'b0110100000: data <= 16'h00a5; 
        10'b0110100001: data <= 16'hffdf; 
        10'b0110100010: data <= 16'hffef; 
        10'b0110100011: data <= 16'hffdc; 
        10'b0110100100: data <= 16'h0012; 
        10'b0110100101: data <= 16'h000a; 
        10'b0110100110: data <= 16'hffe2; 
        10'b0110100111: data <= 16'hfff9; 
        10'b0110101000: data <= 16'hfffe; 
        10'b0110101001: data <= 16'h00cf; 
        10'b0110101010: data <= 16'h0096; 
        10'b0110101011: data <= 16'h00cf; 
        10'b0110101100: data <= 16'h008f; 
        10'b0110101101: data <= 16'h00bd; 
        10'b0110101110: data <= 16'h00ef; 
        10'b0110101111: data <= 16'h0042; 
        10'b0110110000: data <= 16'hff4c; 
        10'b0110110001: data <= 16'hfe34; 
        10'b0110110010: data <= 16'hfd9a; 
        10'b0110110011: data <= 16'hfdb8; 
        10'b0110110100: data <= 16'hfe75; 
        10'b0110110101: data <= 16'hff3f; 
        10'b0110110110: data <= 16'hffb8; 
        10'b0110110111: data <= 16'hffba; 
        10'b0110111000: data <= 16'h003c; 
        10'b0110111001: data <= 16'h0035; 
        10'b0110111010: data <= 16'h00c9; 
        10'b0110111011: data <= 16'h00ed; 
        10'b0110111100: data <= 16'h007b; 
        10'b0110111101: data <= 16'hfff4; 
        10'b0110111110: data <= 16'h0003; 
        10'b0110111111: data <= 16'hffe0; 
        10'b0111000000: data <= 16'h0005; 
        10'b0111000001: data <= 16'h0017; 
        10'b0111000010: data <= 16'hffd1; 
        10'b0111000011: data <= 16'hffe7; 
        10'b0111000100: data <= 16'h0023; 
        10'b0111000101: data <= 16'h00bc; 
        10'b0111000110: data <= 16'h00ea; 
        10'b0111000111: data <= 16'h00b5; 
        10'b0111001000: data <= 16'h007d; 
        10'b0111001001: data <= 16'h007e; 
        10'b0111001010: data <= 16'h00d5; 
        10'b0111001011: data <= 16'hffe4; 
        10'b0111001100: data <= 16'hfea2; 
        10'b0111001101: data <= 16'hfd9f; 
        10'b0111001110: data <= 16'hfdaf; 
        10'b0111001111: data <= 16'hfe29; 
        10'b0111010000: data <= 16'hff04; 
        10'b0111010001: data <= 16'hff8a; 
        10'b0111010010: data <= 16'hfffe; 
        10'b0111010011: data <= 16'h0027; 
        10'b0111010100: data <= 16'h0059; 
        10'b0111010101: data <= 16'h0084; 
        10'b0111010110: data <= 16'h00b5; 
        10'b0111010111: data <= 16'h00ad; 
        10'b0111011000: data <= 16'h0042; 
        10'b0111011001: data <= 16'h0003; 
        10'b0111011010: data <= 16'hffeb; 
        10'b0111011011: data <= 16'hffe3; 
        10'b0111011100: data <= 16'hffef; 
        10'b0111011101: data <= 16'h0006; 
        10'b0111011110: data <= 16'hffd8; 
        10'b0111011111: data <= 16'hffb3; 
        10'b0111100000: data <= 16'h0007; 
        10'b0111100001: data <= 16'h0086; 
        10'b0111100010: data <= 16'h00a8; 
        10'b0111100011: data <= 16'h00a3; 
        10'b0111100100: data <= 16'h0033; 
        10'b0111100101: data <= 16'h0083; 
        10'b0111100110: data <= 16'h00cf; 
        10'b0111100111: data <= 16'hffe0; 
        10'b0111101000: data <= 16'hfe5c; 
        10'b0111101001: data <= 16'hfda7; 
        10'b0111101010: data <= 16'hfdef; 
        10'b0111101011: data <= 16'hfec5; 
        10'b0111101100: data <= 16'hffd7; 
        10'b0111101101: data <= 16'h0050; 
        10'b0111101110: data <= 16'h0074; 
        10'b0111101111: data <= 16'h006b; 
        10'b0111110000: data <= 16'h0088; 
        10'b0111110001: data <= 16'h0068; 
        10'b0111110010: data <= 16'h0052; 
        10'b0111110011: data <= 16'h005d; 
        10'b0111110100: data <= 16'hfffb; 
        10'b0111110101: data <= 16'hfff2; 
        10'b0111110110: data <= 16'h0007; 
        10'b0111110111: data <= 16'hffdf; 
        10'b0111111000: data <= 16'hffea; 
        10'b0111111001: data <= 16'h0007; 
        10'b0111111010: data <= 16'hfff0; 
        10'b0111111011: data <= 16'hffe3; 
        10'b0111111100: data <= 16'hfff0; 
        10'b0111111101: data <= 16'h0055; 
        10'b0111111110: data <= 16'h00ae; 
        10'b0111111111: data <= 16'h0064; 
        10'b1000000000: data <= 16'h003e; 
        10'b1000000001: data <= 16'h00ad; 
        10'b1000000010: data <= 16'h014b; 
        10'b1000000011: data <= 16'h000d; 
        10'b1000000100: data <= 16'hfef5; 
        10'b1000000101: data <= 16'hfe51; 
        10'b1000000110: data <= 16'hfed3; 
        10'b1000000111: data <= 16'hffa4; 
        10'b1000001000: data <= 16'h0061; 
        10'b1000001001: data <= 16'h0068; 
        10'b1000001010: data <= 16'h006c; 
        10'b1000001011: data <= 16'h0038; 
        10'b1000001100: data <= 16'h001c; 
        10'b1000001101: data <= 16'h002f; 
        10'b1000001110: data <= 16'h005a; 
        10'b1000001111: data <= 16'h0038; 
        10'b1000010000: data <= 16'hfff9; 
        10'b1000010001: data <= 16'hffe4; 
        10'b1000010010: data <= 16'h0003; 
        10'b1000010011: data <= 16'hfff0; 
        10'b1000010100: data <= 16'hfff2; 
        10'b1000010101: data <= 16'hffed; 
        10'b1000010110: data <= 16'hffef; 
        10'b1000010111: data <= 16'hffb5; 
        10'b1000011000: data <= 16'h0020; 
        10'b1000011001: data <= 16'h005d; 
        10'b1000011010: data <= 16'h00df; 
        10'b1000011011: data <= 16'h00cb; 
        10'b1000011100: data <= 16'h009f; 
        10'b1000011101: data <= 16'h00d2; 
        10'b1000011110: data <= 16'h014c; 
        10'b1000011111: data <= 16'h00e9; 
        10'b1000100000: data <= 16'h0031; 
        10'b1000100001: data <= 16'hff95; 
        10'b1000100010: data <= 16'hffd1; 
        10'b1000100011: data <= 16'hffe2; 
        10'b1000100100: data <= 16'h0033; 
        10'b1000100101: data <= 16'hffe9; 
        10'b1000100110: data <= 16'hffd5; 
        10'b1000100111: data <= 16'hffe6; 
        10'b1000101000: data <= 16'h0034; 
        10'b1000101001: data <= 16'h0030; 
        10'b1000101010: data <= 16'h005d; 
        10'b1000101011: data <= 16'hfff4; 
        10'b1000101100: data <= 16'h000d; 
        10'b1000101101: data <= 16'hffec; 
        10'b1000101110: data <= 16'hffd0; 
        10'b1000101111: data <= 16'h0011; 
        10'b1000110000: data <= 16'h0010; 
        10'b1000110001: data <= 16'h0016; 
        10'b1000110010: data <= 16'hfff0; 
        10'b1000110011: data <= 16'hffdc; 
        10'b1000110100: data <= 16'hffeb; 
        10'b1000110101: data <= 16'h0060; 
        10'b1000110110: data <= 16'h00b3; 
        10'b1000110111: data <= 16'h0084; 
        10'b1000111000: data <= 16'h00a4; 
        10'b1000111001: data <= 16'h00c9; 
        10'b1000111010: data <= 16'h0139; 
        10'b1000111011: data <= 16'h0139; 
        10'b1000111100: data <= 16'h009d; 
        10'b1000111101: data <= 16'h0030; 
        10'b1000111110: data <= 16'hffdf; 
        10'b1000111111: data <= 16'h0017; 
        10'b1001000000: data <= 16'h0015; 
        10'b1001000001: data <= 16'hffd2; 
        10'b1001000010: data <= 16'hffdd; 
        10'b1001000011: data <= 16'hffcf; 
        10'b1001000100: data <= 16'h001a; 
        10'b1001000101: data <= 16'h0020; 
        10'b1001000110: data <= 16'h0031; 
        10'b1001000111: data <= 16'h0011; 
        10'b1001001000: data <= 16'hffe4; 
        10'b1001001001: data <= 16'hfffa; 
        10'b1001001010: data <= 16'hffd9; 
        10'b1001001011: data <= 16'hffec; 
        10'b1001001100: data <= 16'hffe3; 
        10'b1001001101: data <= 16'hffd5; 
        10'b1001001110: data <= 16'hfff1; 
        10'b1001001111: data <= 16'hffe4; 
        10'b1001010000: data <= 16'hffee; 
        10'b1001010001: data <= 16'h0019; 
        10'b1001010010: data <= 16'h006f; 
        10'b1001010011: data <= 16'h00b4; 
        10'b1001010100: data <= 16'h007e; 
        10'b1001010101: data <= 16'h0089; 
        10'b1001010110: data <= 16'h010c; 
        10'b1001010111: data <= 16'h012f; 
        10'b1001011000: data <= 16'h00c9; 
        10'b1001011001: data <= 16'h004c; 
        10'b1001011010: data <= 16'h001c; 
        10'b1001011011: data <= 16'h0006; 
        10'b1001011100: data <= 16'hfffb; 
        10'b1001011101: data <= 16'hffad; 
        10'b1001011110: data <= 16'hffc1; 
        10'b1001011111: data <= 16'hffdc; 
        10'b1001100000: data <= 16'h0020; 
        10'b1001100001: data <= 16'hfffe; 
        10'b1001100010: data <= 16'hffda; 
        10'b1001100011: data <= 16'hffc4; 
        10'b1001100100: data <= 16'hfff1; 
        10'b1001100101: data <= 16'hffec; 
        10'b1001100110: data <= 16'hffe3; 
        10'b1001100111: data <= 16'hffe7; 
        10'b1001101000: data <= 16'hffdc; 
        10'b1001101001: data <= 16'h0002; 
        10'b1001101010: data <= 16'h0003; 
        10'b1001101011: data <= 16'hffeb; 
        10'b1001101100: data <= 16'hffda; 
        10'b1001101101: data <= 16'h000e; 
        10'b1001101110: data <= 16'h0051; 
        10'b1001101111: data <= 16'h0046; 
        10'b1001110000: data <= 16'h00ca; 
        10'b1001110001: data <= 16'h00a4; 
        10'b1001110010: data <= 16'h00b5; 
        10'b1001110011: data <= 16'h00d8; 
        10'b1001110100: data <= 16'h00b8; 
        10'b1001110101: data <= 16'h00ec; 
        10'b1001110110: data <= 16'h0066; 
        10'b1001110111: data <= 16'h0069; 
        10'b1001111000: data <= 16'h0039; 
        10'b1001111001: data <= 16'hffcf; 
        10'b1001111010: data <= 16'hffd9; 
        10'b1001111011: data <= 16'hfffd; 
        10'b1001111100: data <= 16'hffc9; 
        10'b1001111101: data <= 16'hffc7; 
        10'b1001111110: data <= 16'hffe4; 
        10'b1001111111: data <= 16'hffe2; 
        10'b1010000000: data <= 16'hfff5; 
        10'b1010000001: data <= 16'hffee; 
        10'b1010000010: data <= 16'hffe8; 
        10'b1010000011: data <= 16'hfff3; 
        10'b1010000100: data <= 16'hffdc; 
        10'b1010000101: data <= 16'hfff6; 
        10'b1010000110: data <= 16'hffff; 
        10'b1010000111: data <= 16'hffd5; 
        10'b1010001000: data <= 16'hffd4; 
        10'b1010001001: data <= 16'hfff3; 
        10'b1010001010: data <= 16'hfffb; 
        10'b1010001011: data <= 16'h0038; 
        10'b1010001100: data <= 16'h004f; 
        10'b1010001101: data <= 16'h00bb; 
        10'b1010001110: data <= 16'h00e0; 
        10'b1010001111: data <= 16'h0112; 
        10'b1010010000: data <= 16'h0110; 
        10'b1010010001: data <= 16'h00a3; 
        10'b1010010010: data <= 16'h0085; 
        10'b1010010011: data <= 16'h0049; 
        10'b1010010100: data <= 16'h001f; 
        10'b1010010101: data <= 16'hfffd; 
        10'b1010010110: data <= 16'hff99; 
        10'b1010010111: data <= 16'hff7e; 
        10'b1010011000: data <= 16'hff9c; 
        10'b1010011001: data <= 16'hffce; 
        10'b1010011010: data <= 16'hffd8; 
        10'b1010011011: data <= 16'hfffb; 
        10'b1010011100: data <= 16'hfff1; 
        10'b1010011101: data <= 16'h000d; 
        10'b1010011110: data <= 16'hffea; 
        10'b1010011111: data <= 16'hffd3; 
        10'b1010100000: data <= 16'hffec; 
        10'b1010100001: data <= 16'hfff7; 
        10'b1010100010: data <= 16'hffd4; 
        10'b1010100011: data <= 16'hfffe; 
        10'b1010100100: data <= 16'hfff4; 
        10'b1010100101: data <= 16'hfff4; 
        10'b1010100110: data <= 16'hffcb; 
        10'b1010100111: data <= 16'hffb9; 
        10'b1010101000: data <= 16'hffd8; 
        10'b1010101001: data <= 16'hffdc; 
        10'b1010101010: data <= 16'h0029; 
        10'b1010101011: data <= 16'h001f; 
        10'b1010101100: data <= 16'h004c; 
        10'b1010101101: data <= 16'h006f; 
        10'b1010101110: data <= 16'h003b; 
        10'b1010101111: data <= 16'hffd3; 
        10'b1010110000: data <= 16'hffbb; 
        10'b1010110001: data <= 16'hffad; 
        10'b1010110010: data <= 16'hffba; 
        10'b1010110011: data <= 16'hff9d; 
        10'b1010110100: data <= 16'hffa2; 
        10'b1010110101: data <= 16'hffa7; 
        10'b1010110110: data <= 16'hffef; 
        10'b1010110111: data <= 16'hffe9; 
        10'b1010111000: data <= 16'hffdb; 
        10'b1010111001: data <= 16'hffe4; 
        10'b1010111010: data <= 16'h0002; 
        10'b1010111011: data <= 16'hffe0; 
        10'b1010111100: data <= 16'hffe5; 
        10'b1010111101: data <= 16'h0019; 
        10'b1010111110: data <= 16'hfff2; 
        10'b1010111111: data <= 16'h0015; 
        10'b1011000000: data <= 16'h0018; 
        10'b1011000001: data <= 16'hffff; 
        10'b1011000010: data <= 16'hffd0; 
        10'b1011000011: data <= 16'hffeb; 
        10'b1011000100: data <= 16'hffa2; 
        10'b1011000101: data <= 16'hffa7; 
        10'b1011000110: data <= 16'hff92; 
        10'b1011000111: data <= 16'hff71; 
        10'b1011001000: data <= 16'hff5c; 
        10'b1011001001: data <= 16'hff6b; 
        10'b1011001010: data <= 16'hff52; 
        10'b1011001011: data <= 16'hff63; 
        10'b1011001100: data <= 16'hff6c; 
        10'b1011001101: data <= 16'hffa7; 
        10'b1011001110: data <= 16'hffb6; 
        10'b1011001111: data <= 16'hffc2; 
        10'b1011010000: data <= 16'hffbb; 
        10'b1011010001: data <= 16'hffc0; 
        10'b1011010010: data <= 16'hffeb; 
        10'b1011010011: data <= 16'h0018; 
        10'b1011010100: data <= 16'h000c; 
        10'b1011010101: data <= 16'hffef; 
        10'b1011010110: data <= 16'hffe9; 
        10'b1011010111: data <= 16'hfff7; 
        10'b1011011000: data <= 16'h0014; 
        10'b1011011001: data <= 16'h0012; 
        10'b1011011010: data <= 16'hffee; 
        10'b1011011011: data <= 16'h0001; 
        10'b1011011100: data <= 16'hffe7; 
        10'b1011011101: data <= 16'hffec; 
        10'b1011011110: data <= 16'hffd5; 
        10'b1011011111: data <= 16'h0009; 
        10'b1011100000: data <= 16'hffe9; 
        10'b1011100001: data <= 16'hffb1; 
        10'b1011100010: data <= 16'hffb1; 
        10'b1011100011: data <= 16'hffb9; 
        10'b1011100100: data <= 16'hffe3; 
        10'b1011100101: data <= 16'hffb9; 
        10'b1011100110: data <= 16'hffbc; 
        10'b1011100111: data <= 16'hffe7; 
        10'b1011101000: data <= 16'hffb8; 
        10'b1011101001: data <= 16'hffc6; 
        10'b1011101010: data <= 16'hffd4; 
        10'b1011101011: data <= 16'hffc9; 
        10'b1011101100: data <= 16'hffe5; 
        10'b1011101101: data <= 16'hffbe; 
        10'b1011101110: data <= 16'hffc8; 
        10'b1011101111: data <= 16'h0016; 
        10'b1011110000: data <= 16'hffde; 
        10'b1011110001: data <= 16'h0006; 
        10'b1011110010: data <= 16'h0012; 
        10'b1011110011: data <= 16'hfffc; 
        10'b1011110100: data <= 16'hffdb; 
        10'b1011110101: data <= 16'h000f; 
        10'b1011110110: data <= 16'hfffa; 
        10'b1011110111: data <= 16'hffec; 
        10'b1011111000: data <= 16'h0013; 
        10'b1011111001: data <= 16'h0004; 
        10'b1011111010: data <= 16'h0007; 
        10'b1011111011: data <= 16'hffd3; 
        10'b1011111100: data <= 16'h0016; 
        10'b1011111101: data <= 16'h0016; 
        10'b1011111110: data <= 16'h0008; 
        10'b1011111111: data <= 16'h0010; 
        10'b1100000000: data <= 16'hfff5; 
        10'b1100000001: data <= 16'hffe5; 
        10'b1100000010: data <= 16'h000f; 
        10'b1100000011: data <= 16'hffd9; 
        10'b1100000100: data <= 16'hfff2; 
        10'b1100000101: data <= 16'hffe5; 
        10'b1100000110: data <= 16'hfff9; 
        10'b1100000111: data <= 16'hffe8; 
        10'b1100001000: data <= 16'hffd2; 
        10'b1100001001: data <= 16'hffd6; 
        10'b1100001010: data <= 16'hffc5; 
        10'b1100001011: data <= 16'hfff2; 
        10'b1100001100: data <= 16'h000a; 
        10'b1100001101: data <= 16'hffda; 
        10'b1100001110: data <= 16'hffd1; 
        10'b1100001111: data <= 16'h000c; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 11) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 17'h1ffbe; 
        10'b0000000001: data <= 17'h00026; 
        10'b0000000010: data <= 17'h1ffeb; 
        10'b0000000011: data <= 17'h1fff6; 
        10'b0000000100: data <= 17'h0002d; 
        10'b0000000101: data <= 17'h1fffb; 
        10'b0000000110: data <= 17'h1ffd6; 
        10'b0000000111: data <= 17'h1ffd3; 
        10'b0000001000: data <= 17'h1fff6; 
        10'b0000001001: data <= 17'h1ffea; 
        10'b0000001010: data <= 17'h00032; 
        10'b0000001011: data <= 17'h1fffc; 
        10'b0000001100: data <= 17'h00017; 
        10'b0000001101: data <= 17'h1ffbf; 
        10'b0000001110: data <= 17'h1fffc; 
        10'b0000001111: data <= 17'h1ffa7; 
        10'b0000010000: data <= 17'h1ffb6; 
        10'b0000010001: data <= 17'h1ffec; 
        10'b0000010010: data <= 17'h1ffb4; 
        10'b0000010011: data <= 17'h00031; 
        10'b0000010100: data <= 17'h1ffb6; 
        10'b0000010101: data <= 17'h1ffe8; 
        10'b0000010110: data <= 17'h1ffb0; 
        10'b0000010111: data <= 17'h1fff8; 
        10'b0000011000: data <= 17'h00019; 
        10'b0000011001: data <= 17'h1ffee; 
        10'b0000011010: data <= 17'h1fffc; 
        10'b0000011011: data <= 17'h1fffd; 
        10'b0000011100: data <= 17'h0001c; 
        10'b0000011101: data <= 17'h00023; 
        10'b0000011110: data <= 17'h0000b; 
        10'b0000011111: data <= 17'h1ffb2; 
        10'b0000100000: data <= 17'h1ffae; 
        10'b0000100001: data <= 17'h00004; 
        10'b0000100010: data <= 17'h1ffbf; 
        10'b0000100011: data <= 17'h1ffee; 
        10'b0000100100: data <= 17'h1ffce; 
        10'b0000100101: data <= 17'h1ffa5; 
        10'b0000100110: data <= 17'h1ffc6; 
        10'b0000100111: data <= 17'h00005; 
        10'b0000101000: data <= 17'h00038; 
        10'b0000101001: data <= 17'h1ffb4; 
        10'b0000101010: data <= 17'h1ffd7; 
        10'b0000101011: data <= 17'h00018; 
        10'b0000101100: data <= 17'h1ffc1; 
        10'b0000101101: data <= 17'h1ffaa; 
        10'b0000101110: data <= 17'h00010; 
        10'b0000101111: data <= 17'h00027; 
        10'b0000110000: data <= 17'h1ffbe; 
        10'b0000110001: data <= 17'h00012; 
        10'b0000110010: data <= 17'h1ffc8; 
        10'b0000110011: data <= 17'h1ffb9; 
        10'b0000110100: data <= 17'h1fff2; 
        10'b0000110101: data <= 17'h00005; 
        10'b0000110110: data <= 17'h1ffe9; 
        10'b0000110111: data <= 17'h00030; 
        10'b0000111000: data <= 17'h1ffad; 
        10'b0000111001: data <= 17'h1ffcd; 
        10'b0000111010: data <= 17'h1ffc8; 
        10'b0000111011: data <= 17'h00018; 
        10'b0000111100: data <= 17'h00006; 
        10'b0000111101: data <= 17'h1ffaa; 
        10'b0000111110: data <= 17'h1ffec; 
        10'b0000111111: data <= 17'h0002e; 
        10'b0001000000: data <= 17'h1ffe4; 
        10'b0001000001: data <= 17'h1ffc3; 
        10'b0001000010: data <= 17'h1ffc5; 
        10'b0001000011: data <= 17'h1ff9b; 
        10'b0001000100: data <= 17'h1ff94; 
        10'b0001000101: data <= 17'h1ffdb; 
        10'b0001000110: data <= 17'h1ff90; 
        10'b0001000111: data <= 17'h1ff71; 
        10'b0001001000: data <= 17'h1ff98; 
        10'b0001001001: data <= 17'h1ffe5; 
        10'b0001001010: data <= 17'h1ffa7; 
        10'b0001001011: data <= 17'h1ff8e; 
        10'b0001001100: data <= 17'h1ffec; 
        10'b0001001101: data <= 17'h00022; 
        10'b0001001110: data <= 17'h00006; 
        10'b0001001111: data <= 17'h1ffc1; 
        10'b0001010000: data <= 17'h0002b; 
        10'b0001010001: data <= 17'h1ffa5; 
        10'b0001010010: data <= 17'h1ffea; 
        10'b0001010011: data <= 17'h00015; 
        10'b0001010100: data <= 17'h1ffab; 
        10'b0001010101: data <= 17'h1ffec; 
        10'b0001010110: data <= 17'h00030; 
        10'b0001010111: data <= 17'h1ffad; 
        10'b0001011000: data <= 17'h1ffc5; 
        10'b0001011001: data <= 17'h00027; 
        10'b0001011010: data <= 17'h00010; 
        10'b0001011011: data <= 17'h00002; 
        10'b0001011100: data <= 17'h00006; 
        10'b0001011101: data <= 17'h1ffea; 
        10'b0001011110: data <= 17'h1ffe3; 
        10'b0001011111: data <= 17'h1ff8f; 
        10'b0001100000: data <= 17'h1ff66; 
        10'b0001100001: data <= 17'h1ffa9; 
        10'b0001100010: data <= 17'h1ff87; 
        10'b0001100011: data <= 17'h1ff77; 
        10'b0001100100: data <= 17'h00017; 
        10'b0001100101: data <= 17'h0000b; 
        10'b0001100110: data <= 17'h1ff68; 
        10'b0001100111: data <= 17'h1ff7e; 
        10'b0001101000: data <= 17'h1ff45; 
        10'b0001101001: data <= 17'h1ff7b; 
        10'b0001101010: data <= 17'h1ff60; 
        10'b0001101011: data <= 17'h1ff91; 
        10'b0001101100: data <= 17'h1ffb3; 
        10'b0001101101: data <= 17'h0001d; 
        10'b0001101110: data <= 17'h0001c; 
        10'b0001101111: data <= 17'h1ffd4; 
        10'b0001110000: data <= 17'h0000b; 
        10'b0001110001: data <= 17'h1ffaa; 
        10'b0001110010: data <= 17'h1ffc3; 
        10'b0001110011: data <= 17'h1ffac; 
        10'b0001110100: data <= 17'h1ffa1; 
        10'b0001110101: data <= 17'h1fff4; 
        10'b0001110110: data <= 17'h1ffe6; 
        10'b0001110111: data <= 17'h1ffaa; 
        10'b0001111000: data <= 17'h1ffe3; 
        10'b0001111001: data <= 17'h1ffed; 
        10'b0001111010: data <= 17'h1ff75; 
        10'b0001111011: data <= 17'h1ff77; 
        10'b0001111100: data <= 17'h1ff79; 
        10'b0001111101: data <= 17'h1ff7f; 
        10'b0001111110: data <= 17'h1ffdd; 
        10'b0001111111: data <= 17'h1fff2; 
        10'b0010000000: data <= 17'h1ff96; 
        10'b0010000001: data <= 17'h1ff9c; 
        10'b0010000010: data <= 17'h1ff99; 
        10'b0010000011: data <= 17'h1ff71; 
        10'b0010000100: data <= 17'h1ffc6; 
        10'b0010000101: data <= 17'h1ff48; 
        10'b0010000110: data <= 17'h1ffb8; 
        10'b0010000111: data <= 17'h1fff6; 
        10'b0010001000: data <= 17'h1ffb0; 
        10'b0010001001: data <= 17'h1ffdc; 
        10'b0010001010: data <= 17'h1ffd1; 
        10'b0010001011: data <= 17'h1fff8; 
        10'b0010001100: data <= 17'h00017; 
        10'b0010001101: data <= 17'h1ffd7; 
        10'b0010001110: data <= 17'h1fffe; 
        10'b0010001111: data <= 17'h1ffb4; 
        10'b0010010000: data <= 17'h1ffeb; 
        10'b0010010001: data <= 17'h1ffdb; 
        10'b0010010010: data <= 17'h1ffe5; 
        10'b0010010011: data <= 17'h1ffc7; 
        10'b0010010100: data <= 17'h1ffe6; 
        10'b0010010101: data <= 17'h1ff99; 
        10'b0010010110: data <= 17'h1ffd1; 
        10'b0010010111: data <= 17'h0001e; 
        10'b0010011000: data <= 17'h00079; 
        10'b0010011001: data <= 17'h00105; 
        10'b0010011010: data <= 17'h0013c; 
        10'b0010011011: data <= 17'h00138; 
        10'b0010011100: data <= 17'h0015f; 
        10'b0010011101: data <= 17'h0017a; 
        10'b0010011110: data <= 17'h00190; 
        10'b0010011111: data <= 17'h0008d; 
        10'b0010100000: data <= 17'h00019; 
        10'b0010100001: data <= 17'h00041; 
        10'b0010100010: data <= 17'h1ffe0; 
        10'b0010100011: data <= 17'h1fffb; 
        10'b0010100100: data <= 17'h1ff55; 
        10'b0010100101: data <= 17'h1ff84; 
        10'b0010100110: data <= 17'h1fff7; 
        10'b0010100111: data <= 17'h1ffbe; 
        10'b0010101000: data <= 17'h1ffde; 
        10'b0010101001: data <= 17'h1fff0; 
        10'b0010101010: data <= 17'h00009; 
        10'b0010101011: data <= 17'h1ffe4; 
        10'b0010101100: data <= 17'h00001; 
        10'b0010101101: data <= 17'h00004; 
        10'b0010101110: data <= 17'h0000a; 
        10'b0010101111: data <= 17'h1fffc; 
        10'b0010110000: data <= 17'h1ffaa; 
        10'b0010110001: data <= 17'h1ff6e; 
        10'b0010110010: data <= 17'h00050; 
        10'b0010110011: data <= 17'h1fff3; 
        10'b0010110100: data <= 17'h000d9; 
        10'b0010110101: data <= 17'h000c0; 
        10'b0010110110: data <= 17'h000b7; 
        10'b0010110111: data <= 17'h00110; 
        10'b0010111000: data <= 17'h0014b; 
        10'b0010111001: data <= 17'h001d5; 
        10'b0010111010: data <= 17'h001b4; 
        10'b0010111011: data <= 17'h00174; 
        10'b0010111100: data <= 17'h00167; 
        10'b0010111101: data <= 17'h0019a; 
        10'b0010111110: data <= 17'h000e8; 
        10'b0010111111: data <= 17'h00053; 
        10'b0011000000: data <= 17'h1ff4e; 
        10'b0011000001: data <= 17'h1ff47; 
        10'b0011000010: data <= 17'h1ff83; 
        10'b0011000011: data <= 17'h00013; 
        10'b0011000100: data <= 17'h0002b; 
        10'b0011000101: data <= 17'h00007; 
        10'b0011000110: data <= 17'h1fff7; 
        10'b0011000111: data <= 17'h1ff93; 
        10'b0011001000: data <= 17'h1ff57; 
        10'b0011001001: data <= 17'h1fff1; 
        10'b0011001010: data <= 17'h1ffbc; 
        10'b0011001011: data <= 17'h00001; 
        10'b0011001100: data <= 17'h1ffb1; 
        10'b0011001101: data <= 17'h1ffe9; 
        10'b0011001110: data <= 17'h0000f; 
        10'b0011001111: data <= 17'h0009b; 
        10'b0011010000: data <= 17'h00142; 
        10'b0011010001: data <= 17'h00128; 
        10'b0011010010: data <= 17'h00079; 
        10'b0011010011: data <= 17'h000bd; 
        10'b0011010100: data <= 17'h0010e; 
        10'b0011010101: data <= 17'h001f8; 
        10'b0011010110: data <= 17'h00173; 
        10'b0011010111: data <= 17'h00144; 
        10'b0011011000: data <= 17'h00085; 
        10'b0011011001: data <= 17'h000ff; 
        10'b0011011010: data <= 17'h00118; 
        10'b0011011011: data <= 17'h0008f; 
        10'b0011011100: data <= 17'h1ff93; 
        10'b0011011101: data <= 17'h1ff4e; 
        10'b0011011110: data <= 17'h1ff60; 
        10'b0011011111: data <= 17'h1fff6; 
        10'b0011100000: data <= 17'h00030; 
        10'b0011100001: data <= 17'h00012; 
        10'b0011100010: data <= 17'h1ffeb; 
        10'b0011100011: data <= 17'h1ffff; 
        10'b0011100100: data <= 17'h1ff84; 
        10'b0011100101: data <= 17'h1ffa0; 
        10'b0011100110: data <= 17'h1ffb1; 
        10'b0011100111: data <= 17'h1ff9f; 
        10'b0011101000: data <= 17'h1ffcd; 
        10'b0011101001: data <= 17'h1ffca; 
        10'b0011101010: data <= 17'h00099; 
        10'b0011101011: data <= 17'h000a1; 
        10'b0011101100: data <= 17'h00052; 
        10'b0011101101: data <= 17'h00023; 
        10'b0011101110: data <= 17'h00039; 
        10'b0011101111: data <= 17'h000e3; 
        10'b0011110000: data <= 17'h00295; 
        10'b0011110001: data <= 17'h0020e; 
        10'b0011110010: data <= 17'h001e8; 
        10'b0011110011: data <= 17'h0009a; 
        10'b0011110100: data <= 17'h00081; 
        10'b0011110101: data <= 17'h00076; 
        10'b0011110110: data <= 17'h00122; 
        10'b0011110111: data <= 17'h001f9; 
        10'b0011111000: data <= 17'h1ffc8; 
        10'b0011111001: data <= 17'h1ff58; 
        10'b0011111010: data <= 17'h1ffef; 
        10'b0011111011: data <= 17'h1ffa8; 
        10'b0011111100: data <= 17'h1fff2; 
        10'b0011111101: data <= 17'h1fff8; 
        10'b0011111110: data <= 17'h0000f; 
        10'b0011111111: data <= 17'h0000b; 
        10'b0100000000: data <= 17'h1ff64; 
        10'b0100000001: data <= 17'h1ff91; 
        10'b0100000010: data <= 17'h1ff61; 
        10'b0100000011: data <= 17'h1ffa5; 
        10'b0100000100: data <= 17'h1ffa6; 
        10'b0100000101: data <= 17'h1ffd2; 
        10'b0100000110: data <= 17'h0006e; 
        10'b0100000111: data <= 17'h1ffa2; 
        10'b0100001000: data <= 17'h00037; 
        10'b0100001001: data <= 17'h000a5; 
        10'b0100001010: data <= 17'h00093; 
        10'b0100001011: data <= 17'h0007d; 
        10'b0100001100: data <= 17'h0016a; 
        10'b0100001101: data <= 17'h001e2; 
        10'b0100001110: data <= 17'h0022a; 
        10'b0100001111: data <= 17'h00141; 
        10'b0100010000: data <= 17'h00062; 
        10'b0100010001: data <= 17'h1ffee; 
        10'b0100010010: data <= 17'h000ee; 
        10'b0100010011: data <= 17'h00201; 
        10'b0100010100: data <= 17'h00096; 
        10'b0100010101: data <= 17'h1ff82; 
        10'b0100010110: data <= 17'h00002; 
        10'b0100010111: data <= 17'h1fff0; 
        10'b0100011000: data <= 17'h1ffaf; 
        10'b0100011001: data <= 17'h00028; 
        10'b0100011010: data <= 17'h1ffbc; 
        10'b0100011011: data <= 17'h1ff84; 
        10'b0100011100: data <= 17'h1ff8e; 
        10'b0100011101: data <= 17'h1ffa6; 
        10'b0100011110: data <= 17'h1ffb4; 
        10'b0100011111: data <= 17'h0000a; 
        10'b0100100000: data <= 17'h00034; 
        10'b0100100001: data <= 17'h1fff4; 
        10'b0100100010: data <= 17'h1ffa9; 
        10'b0100100011: data <= 17'h0001c; 
        10'b0100100100: data <= 17'h00024; 
        10'b0100100101: data <= 17'h1ffeb; 
        10'b0100100110: data <= 17'h1ff52; 
        10'b0100100111: data <= 17'h1fed5; 
        10'b0100101000: data <= 17'h1ff4c; 
        10'b0100101001: data <= 17'h000ae; 
        10'b0100101010: data <= 17'h001b9; 
        10'b0100101011: data <= 17'h001c9; 
        10'b0100101100: data <= 17'h00194; 
        10'b0100101101: data <= 17'h00125; 
        10'b0100101110: data <= 17'h001b2; 
        10'b0100101111: data <= 17'h00252; 
        10'b0100110000: data <= 17'h0011b; 
        10'b0100110001: data <= 17'h1ff8b; 
        10'b0100110010: data <= 17'h1ff8b; 
        10'b0100110011: data <= 17'h1ffa7; 
        10'b0100110100: data <= 17'h1ffc3; 
        10'b0100110101: data <= 17'h1ffaf; 
        10'b0100110110: data <= 17'h00022; 
        10'b0100110111: data <= 17'h1ffe7; 
        10'b0100111000: data <= 17'h1ff21; 
        10'b0100111001: data <= 17'h1ffd0; 
        10'b0100111010: data <= 17'h00023; 
        10'b0100111011: data <= 17'h000a8; 
        10'b0100111100: data <= 17'h0007e; 
        10'b0100111101: data <= 17'h1ffd0; 
        10'b0100111110: data <= 17'h0002c; 
        10'b0100111111: data <= 17'h00004; 
        10'b0101000000: data <= 17'h00057; 
        10'b0101000001: data <= 17'h1ffc5; 
        10'b0101000010: data <= 17'h1fe27; 
        10'b0101000011: data <= 17'h1fc95; 
        10'b0101000100: data <= 17'h1fcc8; 
        10'b0101000101: data <= 17'h1febe; 
        10'b0101000110: data <= 17'h1ffd5; 
        10'b0101000111: data <= 17'h000e8; 
        10'b0101001000: data <= 17'h00174; 
        10'b0101001001: data <= 17'h00158; 
        10'b0101001010: data <= 17'h001d6; 
        10'b0101001011: data <= 17'h00215; 
        10'b0101001100: data <= 17'h0017f; 
        10'b0101001101: data <= 17'h1ffb6; 
        10'b0101001110: data <= 17'h1fffb; 
        10'b0101001111: data <= 17'h1ffa1; 
        10'b0101010000: data <= 17'h1ffc0; 
        10'b0101010001: data <= 17'h1ffec; 
        10'b0101010010: data <= 17'h1ffe3; 
        10'b0101010011: data <= 17'h1ffe8; 
        10'b0101010100: data <= 17'h1ff82; 
        10'b0101010101: data <= 17'h00014; 
        10'b0101010110: data <= 17'h000b7; 
        10'b0101010111: data <= 17'h000c0; 
        10'b0101011000: data <= 17'h0005d; 
        10'b0101011001: data <= 17'h1ffe6; 
        10'b0101011010: data <= 17'h00083; 
        10'b0101011011: data <= 17'h0005d; 
        10'b0101011100: data <= 17'h000ac; 
        10'b0101011101: data <= 17'h1ff73; 
        10'b0101011110: data <= 17'h1fc61; 
        10'b0101011111: data <= 17'h1fb83; 
        10'b0101100000: data <= 17'h1fb88; 
        10'b0101100001: data <= 17'h1fd8f; 
        10'b0101100010: data <= 17'h1ff91; 
        10'b0101100011: data <= 17'h1ffd2; 
        10'b0101100100: data <= 17'h00038; 
        10'b0101100101: data <= 17'h000a0; 
        10'b0101100110: data <= 17'h00261; 
        10'b0101100111: data <= 17'h0022d; 
        10'b0101101000: data <= 17'h00183; 
        10'b0101101001: data <= 17'h0000e; 
        10'b0101101010: data <= 17'h1ffc3; 
        10'b0101101011: data <= 17'h1ffc2; 
        10'b0101101100: data <= 17'h1ffa5; 
        10'b0101101101: data <= 17'h1fffe; 
        10'b0101101110: data <= 17'h00020; 
        10'b0101101111: data <= 17'h1ffa9; 
        10'b0101110000: data <= 17'h1ffdf; 
        10'b0101110001: data <= 17'h00072; 
        10'b0101110010: data <= 17'h000de; 
        10'b0101110011: data <= 17'h0011f; 
        10'b0101110100: data <= 17'h000d9; 
        10'b0101110101: data <= 17'h00098; 
        10'b0101110110: data <= 17'h000cf; 
        10'b0101110111: data <= 17'h000a1; 
        10'b0101111000: data <= 17'h00074; 
        10'b0101111001: data <= 17'h1fdcb; 
        10'b0101111010: data <= 17'h1fc5f; 
        10'b0101111011: data <= 17'h1fb64; 
        10'b0101111100: data <= 17'h1fc37; 
        10'b0101111101: data <= 17'h1fe1f; 
        10'b0101111110: data <= 17'h1ff15; 
        10'b0101111111: data <= 17'h1fec4; 
        10'b0110000000: data <= 17'h1ff0f; 
        10'b0110000001: data <= 17'h0006a; 
        10'b0110000010: data <= 17'h00190; 
        10'b0110000011: data <= 17'h00273; 
        10'b0110000100: data <= 17'h00164; 
        10'b0110000101: data <= 17'h00039; 
        10'b0110000110: data <= 17'h00000; 
        10'b0110000111: data <= 17'h00023; 
        10'b0110001000: data <= 17'h1fff3; 
        10'b0110001001: data <= 17'h0001b; 
        10'b0110001010: data <= 17'h1ffba; 
        10'b0110001011: data <= 17'h1ffce; 
        10'b0110001100: data <= 17'h1ff94; 
        10'b0110001101: data <= 17'h00125; 
        10'b0110001110: data <= 17'h0017d; 
        10'b0110001111: data <= 17'h001cf; 
        10'b0110010000: data <= 17'h000de; 
        10'b0110010001: data <= 17'h0010b; 
        10'b0110010010: data <= 17'h00188; 
        10'b0110010011: data <= 17'h000e1; 
        10'b0110010100: data <= 17'h00037; 
        10'b0110010101: data <= 17'h1fe15; 
        10'b0110010110: data <= 17'h1fbb9; 
        10'b0110010111: data <= 17'h1fb60; 
        10'b0110011000: data <= 17'h1fc52; 
        10'b0110011001: data <= 17'h1fdfd; 
        10'b0110011010: data <= 17'h1ff1d; 
        10'b0110011011: data <= 17'h1feee; 
        10'b0110011100: data <= 17'h00019; 
        10'b0110011101: data <= 17'h000df; 
        10'b0110011110: data <= 17'h0010a; 
        10'b0110011111: data <= 17'h0027a; 
        10'b0110100000: data <= 17'h0014a; 
        10'b0110100001: data <= 17'h1ffbd; 
        10'b0110100010: data <= 17'h1ffdf; 
        10'b0110100011: data <= 17'h1ffb9; 
        10'b0110100100: data <= 17'h00025; 
        10'b0110100101: data <= 17'h00014; 
        10'b0110100110: data <= 17'h1ffc4; 
        10'b0110100111: data <= 17'h1fff2; 
        10'b0110101000: data <= 17'h1fffb; 
        10'b0110101001: data <= 17'h0019e; 
        10'b0110101010: data <= 17'h0012d; 
        10'b0110101011: data <= 17'h0019e; 
        10'b0110101100: data <= 17'h0011e; 
        10'b0110101101: data <= 17'h0017b; 
        10'b0110101110: data <= 17'h001df; 
        10'b0110101111: data <= 17'h00084; 
        10'b0110110000: data <= 17'h1fe97; 
        10'b0110110001: data <= 17'h1fc69; 
        10'b0110110010: data <= 17'h1fb35; 
        10'b0110110011: data <= 17'h1fb6f; 
        10'b0110110100: data <= 17'h1fceb; 
        10'b0110110101: data <= 17'h1fe7f; 
        10'b0110110110: data <= 17'h1ff70; 
        10'b0110110111: data <= 17'h1ff75; 
        10'b0110111000: data <= 17'h00078; 
        10'b0110111001: data <= 17'h00069; 
        10'b0110111010: data <= 17'h00193; 
        10'b0110111011: data <= 17'h001d9; 
        10'b0110111100: data <= 17'h000f5; 
        10'b0110111101: data <= 17'h1ffe8; 
        10'b0110111110: data <= 17'h00007; 
        10'b0110111111: data <= 17'h1ffbf; 
        10'b0111000000: data <= 17'h0000b; 
        10'b0111000001: data <= 17'h0002e; 
        10'b0111000010: data <= 17'h1ffa2; 
        10'b0111000011: data <= 17'h1ffcd; 
        10'b0111000100: data <= 17'h00046; 
        10'b0111000101: data <= 17'h00178; 
        10'b0111000110: data <= 17'h001d3; 
        10'b0111000111: data <= 17'h00169; 
        10'b0111001000: data <= 17'h000fb; 
        10'b0111001001: data <= 17'h000fd; 
        10'b0111001010: data <= 17'h001ab; 
        10'b0111001011: data <= 17'h1ffc8; 
        10'b0111001100: data <= 17'h1fd44; 
        10'b0111001101: data <= 17'h1fb3e; 
        10'b0111001110: data <= 17'h1fb5e; 
        10'b0111001111: data <= 17'h1fc53; 
        10'b0111010000: data <= 17'h1fe08; 
        10'b0111010001: data <= 17'h1ff15; 
        10'b0111010010: data <= 17'h1fffd; 
        10'b0111010011: data <= 17'h0004d; 
        10'b0111010100: data <= 17'h000b1; 
        10'b0111010101: data <= 17'h00108; 
        10'b0111010110: data <= 17'h0016b; 
        10'b0111010111: data <= 17'h0015a; 
        10'b0111011000: data <= 17'h00084; 
        10'b0111011001: data <= 17'h00006; 
        10'b0111011010: data <= 17'h1ffd5; 
        10'b0111011011: data <= 17'h1ffc6; 
        10'b0111011100: data <= 17'h1ffde; 
        10'b0111011101: data <= 17'h0000b; 
        10'b0111011110: data <= 17'h1ffb1; 
        10'b0111011111: data <= 17'h1ff66; 
        10'b0111100000: data <= 17'h0000d; 
        10'b0111100001: data <= 17'h0010b; 
        10'b0111100010: data <= 17'h0014f; 
        10'b0111100011: data <= 17'h00146; 
        10'b0111100100: data <= 17'h00066; 
        10'b0111100101: data <= 17'h00105; 
        10'b0111100110: data <= 17'h0019d; 
        10'b0111100111: data <= 17'h1ffc1; 
        10'b0111101000: data <= 17'h1fcb9; 
        10'b0111101001: data <= 17'h1fb4e; 
        10'b0111101010: data <= 17'h1fbde; 
        10'b0111101011: data <= 17'h1fd89; 
        10'b0111101100: data <= 17'h1ffad; 
        10'b0111101101: data <= 17'h000a1; 
        10'b0111101110: data <= 17'h000e8; 
        10'b0111101111: data <= 17'h000d6; 
        10'b0111110000: data <= 17'h00110; 
        10'b0111110001: data <= 17'h000d0; 
        10'b0111110010: data <= 17'h000a4; 
        10'b0111110011: data <= 17'h000ba; 
        10'b0111110100: data <= 17'h1fff6; 
        10'b0111110101: data <= 17'h1ffe4; 
        10'b0111110110: data <= 17'h0000e; 
        10'b0111110111: data <= 17'h1ffbf; 
        10'b0111111000: data <= 17'h1ffd3; 
        10'b0111111001: data <= 17'h0000f; 
        10'b0111111010: data <= 17'h1ffe1; 
        10'b0111111011: data <= 17'h1ffc5; 
        10'b0111111100: data <= 17'h1ffe0; 
        10'b0111111101: data <= 17'h000aa; 
        10'b0111111110: data <= 17'h0015b; 
        10'b0111111111: data <= 17'h000c9; 
        10'b1000000000: data <= 17'h0007b; 
        10'b1000000001: data <= 17'h00159; 
        10'b1000000010: data <= 17'h00296; 
        10'b1000000011: data <= 17'h0001a; 
        10'b1000000100: data <= 17'h1fde9; 
        10'b1000000101: data <= 17'h1fca1; 
        10'b1000000110: data <= 17'h1fda7; 
        10'b1000000111: data <= 17'h1ff49; 
        10'b1000001000: data <= 17'h000c2; 
        10'b1000001001: data <= 17'h000cf; 
        10'b1000001010: data <= 17'h000d9; 
        10'b1000001011: data <= 17'h00071; 
        10'b1000001100: data <= 17'h00038; 
        10'b1000001101: data <= 17'h0005e; 
        10'b1000001110: data <= 17'h000b5; 
        10'b1000001111: data <= 17'h00071; 
        10'b1000010000: data <= 17'h1fff2; 
        10'b1000010001: data <= 17'h1ffc9; 
        10'b1000010010: data <= 17'h00007; 
        10'b1000010011: data <= 17'h1ffe1; 
        10'b1000010100: data <= 17'h1ffe4; 
        10'b1000010101: data <= 17'h1ffd9; 
        10'b1000010110: data <= 17'h1ffdd; 
        10'b1000010111: data <= 17'h1ff6a; 
        10'b1000011000: data <= 17'h00040; 
        10'b1000011001: data <= 17'h000bb; 
        10'b1000011010: data <= 17'h001be; 
        10'b1000011011: data <= 17'h00195; 
        10'b1000011100: data <= 17'h0013d; 
        10'b1000011101: data <= 17'h001a5; 
        10'b1000011110: data <= 17'h00298; 
        10'b1000011111: data <= 17'h001d3; 
        10'b1000100000: data <= 17'h00063; 
        10'b1000100001: data <= 17'h1ff29; 
        10'b1000100010: data <= 17'h1ffa2; 
        10'b1000100011: data <= 17'h1ffc4; 
        10'b1000100100: data <= 17'h00065; 
        10'b1000100101: data <= 17'h1ffd1; 
        10'b1000100110: data <= 17'h1ffaa; 
        10'b1000100111: data <= 17'h1ffcc; 
        10'b1000101000: data <= 17'h00068; 
        10'b1000101001: data <= 17'h0005f; 
        10'b1000101010: data <= 17'h000ba; 
        10'b1000101011: data <= 17'h1ffe7; 
        10'b1000101100: data <= 17'h0001b; 
        10'b1000101101: data <= 17'h1ffd7; 
        10'b1000101110: data <= 17'h1ffa0; 
        10'b1000101111: data <= 17'h00021; 
        10'b1000110000: data <= 17'h00021; 
        10'b1000110001: data <= 17'h0002b; 
        10'b1000110010: data <= 17'h1ffe1; 
        10'b1000110011: data <= 17'h1ffb9; 
        10'b1000110100: data <= 17'h1ffd6; 
        10'b1000110101: data <= 17'h000bf; 
        10'b1000110110: data <= 17'h00167; 
        10'b1000110111: data <= 17'h00108; 
        10'b1000111000: data <= 17'h00147; 
        10'b1000111001: data <= 17'h00192; 
        10'b1000111010: data <= 17'h00273; 
        10'b1000111011: data <= 17'h00272; 
        10'b1000111100: data <= 17'h0013a; 
        10'b1000111101: data <= 17'h00060; 
        10'b1000111110: data <= 17'h1ffbf; 
        10'b1000111111: data <= 17'h0002d; 
        10'b1001000000: data <= 17'h0002b; 
        10'b1001000001: data <= 17'h1ffa5; 
        10'b1001000010: data <= 17'h1ffbb; 
        10'b1001000011: data <= 17'h1ff9f; 
        10'b1001000100: data <= 17'h00034; 
        10'b1001000101: data <= 17'h00040; 
        10'b1001000110: data <= 17'h00063; 
        10'b1001000111: data <= 17'h00022; 
        10'b1001001000: data <= 17'h1ffc9; 
        10'b1001001001: data <= 17'h1fff3; 
        10'b1001001010: data <= 17'h1ffb2; 
        10'b1001001011: data <= 17'h1ffd8; 
        10'b1001001100: data <= 17'h1ffc6; 
        10'b1001001101: data <= 17'h1ffab; 
        10'b1001001110: data <= 17'h1ffe2; 
        10'b1001001111: data <= 17'h1ffc8; 
        10'b1001010000: data <= 17'h1ffdc; 
        10'b1001010001: data <= 17'h00032; 
        10'b1001010010: data <= 17'h000de; 
        10'b1001010011: data <= 17'h00168; 
        10'b1001010100: data <= 17'h000fd; 
        10'b1001010101: data <= 17'h00112; 
        10'b1001010110: data <= 17'h00219; 
        10'b1001010111: data <= 17'h0025f; 
        10'b1001011000: data <= 17'h00192; 
        10'b1001011001: data <= 17'h00098; 
        10'b1001011010: data <= 17'h00039; 
        10'b1001011011: data <= 17'h0000c; 
        10'b1001011100: data <= 17'h1fff6; 
        10'b1001011101: data <= 17'h1ff5a; 
        10'b1001011110: data <= 17'h1ff81; 
        10'b1001011111: data <= 17'h1ffb7; 
        10'b1001100000: data <= 17'h0003f; 
        10'b1001100001: data <= 17'h1fffb; 
        10'b1001100010: data <= 17'h1ffb5; 
        10'b1001100011: data <= 17'h1ff88; 
        10'b1001100100: data <= 17'h1ffe2; 
        10'b1001100101: data <= 17'h1ffd8; 
        10'b1001100110: data <= 17'h1ffc6; 
        10'b1001100111: data <= 17'h1ffce; 
        10'b1001101000: data <= 17'h1ffb8; 
        10'b1001101001: data <= 17'h00004; 
        10'b1001101010: data <= 17'h00007; 
        10'b1001101011: data <= 17'h1ffd6; 
        10'b1001101100: data <= 17'h1ffb4; 
        10'b1001101101: data <= 17'h0001c; 
        10'b1001101110: data <= 17'h000a1; 
        10'b1001101111: data <= 17'h0008c; 
        10'b1001110000: data <= 17'h00194; 
        10'b1001110001: data <= 17'h00149; 
        10'b1001110010: data <= 17'h0016a; 
        10'b1001110011: data <= 17'h001af; 
        10'b1001110100: data <= 17'h00170; 
        10'b1001110101: data <= 17'h001d9; 
        10'b1001110110: data <= 17'h000cd; 
        10'b1001110111: data <= 17'h000d1; 
        10'b1001111000: data <= 17'h00073; 
        10'b1001111001: data <= 17'h1ff9f; 
        10'b1001111010: data <= 17'h1ffb3; 
        10'b1001111011: data <= 17'h1fffa; 
        10'b1001111100: data <= 17'h1ff93; 
        10'b1001111101: data <= 17'h1ff8d; 
        10'b1001111110: data <= 17'h1ffc9; 
        10'b1001111111: data <= 17'h1ffc4; 
        10'b1010000000: data <= 17'h1ffeb; 
        10'b1010000001: data <= 17'h1ffdb; 
        10'b1010000010: data <= 17'h1ffd0; 
        10'b1010000011: data <= 17'h1ffe7; 
        10'b1010000100: data <= 17'h1ffb8; 
        10'b1010000101: data <= 17'h1ffed; 
        10'b1010000110: data <= 17'h1fffe; 
        10'b1010000111: data <= 17'h1ffa9; 
        10'b1010001000: data <= 17'h1ffa7; 
        10'b1010001001: data <= 17'h1ffe6; 
        10'b1010001010: data <= 17'h1fff5; 
        10'b1010001011: data <= 17'h00070; 
        10'b1010001100: data <= 17'h0009e; 
        10'b1010001101: data <= 17'h00177; 
        10'b1010001110: data <= 17'h001c1; 
        10'b1010001111: data <= 17'h00225; 
        10'b1010010000: data <= 17'h0021f; 
        10'b1010010001: data <= 17'h00146; 
        10'b1010010010: data <= 17'h00109; 
        10'b1010010011: data <= 17'h00093; 
        10'b1010010100: data <= 17'h0003e; 
        10'b1010010101: data <= 17'h1fffa; 
        10'b1010010110: data <= 17'h1ff31; 
        10'b1010010111: data <= 17'h1fefd; 
        10'b1010011000: data <= 17'h1ff37; 
        10'b1010011001: data <= 17'h1ff9d; 
        10'b1010011010: data <= 17'h1ffaf; 
        10'b1010011011: data <= 17'h1fff6; 
        10'b1010011100: data <= 17'h1ffe1; 
        10'b1010011101: data <= 17'h00019; 
        10'b1010011110: data <= 17'h1ffd5; 
        10'b1010011111: data <= 17'h1ffa6; 
        10'b1010100000: data <= 17'h1ffd8; 
        10'b1010100001: data <= 17'h1ffee; 
        10'b1010100010: data <= 17'h1ffa7; 
        10'b1010100011: data <= 17'h1fffc; 
        10'b1010100100: data <= 17'h1ffe8; 
        10'b1010100101: data <= 17'h1ffe9; 
        10'b1010100110: data <= 17'h1ff95; 
        10'b1010100111: data <= 17'h1ff71; 
        10'b1010101000: data <= 17'h1ffb1; 
        10'b1010101001: data <= 17'h1ffb9; 
        10'b1010101010: data <= 17'h00053; 
        10'b1010101011: data <= 17'h0003f; 
        10'b1010101100: data <= 17'h00098; 
        10'b1010101101: data <= 17'h000de; 
        10'b1010101110: data <= 17'h00075; 
        10'b1010101111: data <= 17'h1ffa7; 
        10'b1010110000: data <= 17'h1ff76; 
        10'b1010110001: data <= 17'h1ff5b; 
        10'b1010110010: data <= 17'h1ff73; 
        10'b1010110011: data <= 17'h1ff3a; 
        10'b1010110100: data <= 17'h1ff44; 
        10'b1010110101: data <= 17'h1ff4e; 
        10'b1010110110: data <= 17'h1ffdd; 
        10'b1010110111: data <= 17'h1ffd1; 
        10'b1010111000: data <= 17'h1ffb5; 
        10'b1010111001: data <= 17'h1ffc9; 
        10'b1010111010: data <= 17'h00004; 
        10'b1010111011: data <= 17'h1ffbf; 
        10'b1010111100: data <= 17'h1ffca; 
        10'b1010111101: data <= 17'h00033; 
        10'b1010111110: data <= 17'h1ffe5; 
        10'b1010111111: data <= 17'h0002a; 
        10'b1011000000: data <= 17'h00030; 
        10'b1011000001: data <= 17'h1fffe; 
        10'b1011000010: data <= 17'h1ffa0; 
        10'b1011000011: data <= 17'h1ffd6; 
        10'b1011000100: data <= 17'h1ff45; 
        10'b1011000101: data <= 17'h1ff4f; 
        10'b1011000110: data <= 17'h1ff23; 
        10'b1011000111: data <= 17'h1fee2; 
        10'b1011001000: data <= 17'h1feb9; 
        10'b1011001001: data <= 17'h1fed6; 
        10'b1011001010: data <= 17'h1fea5; 
        10'b1011001011: data <= 17'h1fec7; 
        10'b1011001100: data <= 17'h1fed8; 
        10'b1011001101: data <= 17'h1ff4e; 
        10'b1011001110: data <= 17'h1ff6c; 
        10'b1011001111: data <= 17'h1ff83; 
        10'b1011010000: data <= 17'h1ff76; 
        10'b1011010001: data <= 17'h1ff80; 
        10'b1011010010: data <= 17'h1ffd5; 
        10'b1011010011: data <= 17'h00030; 
        10'b1011010100: data <= 17'h00017; 
        10'b1011010101: data <= 17'h1ffde; 
        10'b1011010110: data <= 17'h1ffd2; 
        10'b1011010111: data <= 17'h1ffef; 
        10'b1011011000: data <= 17'h00028; 
        10'b1011011001: data <= 17'h00024; 
        10'b1011011010: data <= 17'h1ffdb; 
        10'b1011011011: data <= 17'h00002; 
        10'b1011011100: data <= 17'h1ffce; 
        10'b1011011101: data <= 17'h1ffd8; 
        10'b1011011110: data <= 17'h1ffa9; 
        10'b1011011111: data <= 17'h00011; 
        10'b1011100000: data <= 17'h1ffd2; 
        10'b1011100001: data <= 17'h1ff63; 
        10'b1011100010: data <= 17'h1ff62; 
        10'b1011100011: data <= 17'h1ff71; 
        10'b1011100100: data <= 17'h1ffc7; 
        10'b1011100101: data <= 17'h1ff72; 
        10'b1011100110: data <= 17'h1ff79; 
        10'b1011100111: data <= 17'h1ffce; 
        10'b1011101000: data <= 17'h1ff70; 
        10'b1011101001: data <= 17'h1ff8b; 
        10'b1011101010: data <= 17'h1ffa9; 
        10'b1011101011: data <= 17'h1ff92; 
        10'b1011101100: data <= 17'h1ffc9; 
        10'b1011101101: data <= 17'h1ff7c; 
        10'b1011101110: data <= 17'h1ff91; 
        10'b1011101111: data <= 17'h0002b; 
        10'b1011110000: data <= 17'h1ffbc; 
        10'b1011110001: data <= 17'h0000d; 
        10'b1011110010: data <= 17'h00024; 
        10'b1011110011: data <= 17'h1fff8; 
        10'b1011110100: data <= 17'h1ffb6; 
        10'b1011110101: data <= 17'h0001e; 
        10'b1011110110: data <= 17'h1fff3; 
        10'b1011110111: data <= 17'h1ffd8; 
        10'b1011111000: data <= 17'h00026; 
        10'b1011111001: data <= 17'h00007; 
        10'b1011111010: data <= 17'h0000d; 
        10'b1011111011: data <= 17'h1ffa5; 
        10'b1011111100: data <= 17'h0002d; 
        10'b1011111101: data <= 17'h0002b; 
        10'b1011111110: data <= 17'h0000f; 
        10'b1011111111: data <= 17'h0001f; 
        10'b1100000000: data <= 17'h1ffea; 
        10'b1100000001: data <= 17'h1ffca; 
        10'b1100000010: data <= 17'h0001e; 
        10'b1100000011: data <= 17'h1ffb2; 
        10'b1100000100: data <= 17'h1ffe3; 
        10'b1100000101: data <= 17'h1ffc9; 
        10'b1100000110: data <= 17'h1fff3; 
        10'b1100000111: data <= 17'h1ffcf; 
        10'b1100001000: data <= 17'h1ffa3; 
        10'b1100001001: data <= 17'h1ffad; 
        10'b1100001010: data <= 17'h1ff8a; 
        10'b1100001011: data <= 17'h1ffe5; 
        10'b1100001100: data <= 17'h00013; 
        10'b1100001101: data <= 17'h1ffb5; 
        10'b1100001110: data <= 17'h1ffa1; 
        10'b1100001111: data <= 17'h00019; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 12) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 18'h3ff7b; 
        10'b0000000001: data <= 18'h0004c; 
        10'b0000000010: data <= 18'h3ffd7; 
        10'b0000000011: data <= 18'h3ffed; 
        10'b0000000100: data <= 18'h00059; 
        10'b0000000101: data <= 18'h3fff7; 
        10'b0000000110: data <= 18'h3ffac; 
        10'b0000000111: data <= 18'h3ffa6; 
        10'b0000001000: data <= 18'h3ffeb; 
        10'b0000001001: data <= 18'h3ffd4; 
        10'b0000001010: data <= 18'h00063; 
        10'b0000001011: data <= 18'h3fff8; 
        10'b0000001100: data <= 18'h0002e; 
        10'b0000001101: data <= 18'h3ff7f; 
        10'b0000001110: data <= 18'h3fff9; 
        10'b0000001111: data <= 18'h3ff4f; 
        10'b0000010000: data <= 18'h3ff6c; 
        10'b0000010001: data <= 18'h3ffd9; 
        10'b0000010010: data <= 18'h3ff68; 
        10'b0000010011: data <= 18'h00063; 
        10'b0000010100: data <= 18'h3ff6b; 
        10'b0000010101: data <= 18'h3ffd1; 
        10'b0000010110: data <= 18'h3ff60; 
        10'b0000010111: data <= 18'h3fff0; 
        10'b0000011000: data <= 18'h00031; 
        10'b0000011001: data <= 18'h3ffdd; 
        10'b0000011010: data <= 18'h3fff9; 
        10'b0000011011: data <= 18'h3fffb; 
        10'b0000011100: data <= 18'h00038; 
        10'b0000011101: data <= 18'h00045; 
        10'b0000011110: data <= 18'h00017; 
        10'b0000011111: data <= 18'h3ff64; 
        10'b0000100000: data <= 18'h3ff5d; 
        10'b0000100001: data <= 18'h00008; 
        10'b0000100010: data <= 18'h3ff7f; 
        10'b0000100011: data <= 18'h3ffdc; 
        10'b0000100100: data <= 18'h3ff9c; 
        10'b0000100101: data <= 18'h3ff49; 
        10'b0000100110: data <= 18'h3ff8b; 
        10'b0000100111: data <= 18'h0000a; 
        10'b0000101000: data <= 18'h0006f; 
        10'b0000101001: data <= 18'h3ff68; 
        10'b0000101010: data <= 18'h3ffad; 
        10'b0000101011: data <= 18'h00030; 
        10'b0000101100: data <= 18'h3ff82; 
        10'b0000101101: data <= 18'h3ff54; 
        10'b0000101110: data <= 18'h00020; 
        10'b0000101111: data <= 18'h0004d; 
        10'b0000110000: data <= 18'h3ff7b; 
        10'b0000110001: data <= 18'h00024; 
        10'b0000110010: data <= 18'h3ff90; 
        10'b0000110011: data <= 18'h3ff71; 
        10'b0000110100: data <= 18'h3ffe4; 
        10'b0000110101: data <= 18'h00009; 
        10'b0000110110: data <= 18'h3ffd3; 
        10'b0000110111: data <= 18'h00060; 
        10'b0000111000: data <= 18'h3ff5a; 
        10'b0000111001: data <= 18'h3ff9a; 
        10'b0000111010: data <= 18'h3ff91; 
        10'b0000111011: data <= 18'h0002f; 
        10'b0000111100: data <= 18'h0000d; 
        10'b0000111101: data <= 18'h3ff55; 
        10'b0000111110: data <= 18'h3ffd7; 
        10'b0000111111: data <= 18'h0005b; 
        10'b0001000000: data <= 18'h3ffc9; 
        10'b0001000001: data <= 18'h3ff85; 
        10'b0001000010: data <= 18'h3ff8a; 
        10'b0001000011: data <= 18'h3ff36; 
        10'b0001000100: data <= 18'h3ff29; 
        10'b0001000101: data <= 18'h3ffb6; 
        10'b0001000110: data <= 18'h3ff21; 
        10'b0001000111: data <= 18'h3fee2; 
        10'b0001001000: data <= 18'h3ff2f; 
        10'b0001001001: data <= 18'h3ffc9; 
        10'b0001001010: data <= 18'h3ff4f; 
        10'b0001001011: data <= 18'h3ff1b; 
        10'b0001001100: data <= 18'h3ffd9; 
        10'b0001001101: data <= 18'h00045; 
        10'b0001001110: data <= 18'h0000d; 
        10'b0001001111: data <= 18'h3ff82; 
        10'b0001010000: data <= 18'h00056; 
        10'b0001010001: data <= 18'h3ff4a; 
        10'b0001010010: data <= 18'h3ffd4; 
        10'b0001010011: data <= 18'h0002a; 
        10'b0001010100: data <= 18'h3ff56; 
        10'b0001010101: data <= 18'h3ffd8; 
        10'b0001010110: data <= 18'h00060; 
        10'b0001010111: data <= 18'h3ff5a; 
        10'b0001011000: data <= 18'h3ff89; 
        10'b0001011001: data <= 18'h0004e; 
        10'b0001011010: data <= 18'h0001f; 
        10'b0001011011: data <= 18'h00004; 
        10'b0001011100: data <= 18'h0000c; 
        10'b0001011101: data <= 18'h3ffd4; 
        10'b0001011110: data <= 18'h3ffc6; 
        10'b0001011111: data <= 18'h3ff1e; 
        10'b0001100000: data <= 18'h3fecb; 
        10'b0001100001: data <= 18'h3ff51; 
        10'b0001100010: data <= 18'h3ff0e; 
        10'b0001100011: data <= 18'h3feee; 
        10'b0001100100: data <= 18'h0002e; 
        10'b0001100101: data <= 18'h00016; 
        10'b0001100110: data <= 18'h3fecf; 
        10'b0001100111: data <= 18'h3fefb; 
        10'b0001101000: data <= 18'h3fe8b; 
        10'b0001101001: data <= 18'h3fef7; 
        10'b0001101010: data <= 18'h3fec0; 
        10'b0001101011: data <= 18'h3ff22; 
        10'b0001101100: data <= 18'h3ff66; 
        10'b0001101101: data <= 18'h0003a; 
        10'b0001101110: data <= 18'h00039; 
        10'b0001101111: data <= 18'h3ffa8; 
        10'b0001110000: data <= 18'h00016; 
        10'b0001110001: data <= 18'h3ff53; 
        10'b0001110010: data <= 18'h3ff86; 
        10'b0001110011: data <= 18'h3ff57; 
        10'b0001110100: data <= 18'h3ff41; 
        10'b0001110101: data <= 18'h3ffe7; 
        10'b0001110110: data <= 18'h3ffcc; 
        10'b0001110111: data <= 18'h3ff55; 
        10'b0001111000: data <= 18'h3ffc6; 
        10'b0001111001: data <= 18'h3ffdb; 
        10'b0001111010: data <= 18'h3feeb; 
        10'b0001111011: data <= 18'h3feee; 
        10'b0001111100: data <= 18'h3fef2; 
        10'b0001111101: data <= 18'h3feff; 
        10'b0001111110: data <= 18'h3ffba; 
        10'b0001111111: data <= 18'h3ffe5; 
        10'b0010000000: data <= 18'h3ff2c; 
        10'b0010000001: data <= 18'h3ff39; 
        10'b0010000010: data <= 18'h3ff33; 
        10'b0010000011: data <= 18'h3fee1; 
        10'b0010000100: data <= 18'h3ff8b; 
        10'b0010000101: data <= 18'h3fe8f; 
        10'b0010000110: data <= 18'h3ff70; 
        10'b0010000111: data <= 18'h3ffec; 
        10'b0010001000: data <= 18'h3ff5f; 
        10'b0010001001: data <= 18'h3ffb8; 
        10'b0010001010: data <= 18'h3ffa2; 
        10'b0010001011: data <= 18'h3fff0; 
        10'b0010001100: data <= 18'h0002d; 
        10'b0010001101: data <= 18'h3ffaf; 
        10'b0010001110: data <= 18'h3fffc; 
        10'b0010001111: data <= 18'h3ff68; 
        10'b0010010000: data <= 18'h3ffd7; 
        10'b0010010001: data <= 18'h3ffb6; 
        10'b0010010010: data <= 18'h3ffca; 
        10'b0010010011: data <= 18'h3ff8d; 
        10'b0010010100: data <= 18'h3ffcc; 
        10'b0010010101: data <= 18'h3ff31; 
        10'b0010010110: data <= 18'h3ffa3; 
        10'b0010010111: data <= 18'h0003d; 
        10'b0010011000: data <= 18'h000f2; 
        10'b0010011001: data <= 18'h0020b; 
        10'b0010011010: data <= 18'h00277; 
        10'b0010011011: data <= 18'h00270; 
        10'b0010011100: data <= 18'h002be; 
        10'b0010011101: data <= 18'h002f4; 
        10'b0010011110: data <= 18'h00320; 
        10'b0010011111: data <= 18'h0011a; 
        10'b0010100000: data <= 18'h00032; 
        10'b0010100001: data <= 18'h00082; 
        10'b0010100010: data <= 18'h3ffbf; 
        10'b0010100011: data <= 18'h3fff7; 
        10'b0010100100: data <= 18'h3feab; 
        10'b0010100101: data <= 18'h3ff08; 
        10'b0010100110: data <= 18'h3ffee; 
        10'b0010100111: data <= 18'h3ff7c; 
        10'b0010101000: data <= 18'h3ffbb; 
        10'b0010101001: data <= 18'h3ffe0; 
        10'b0010101010: data <= 18'h00012; 
        10'b0010101011: data <= 18'h3ffc7; 
        10'b0010101100: data <= 18'h00003; 
        10'b0010101101: data <= 18'h00009; 
        10'b0010101110: data <= 18'h00014; 
        10'b0010101111: data <= 18'h3fff8; 
        10'b0010110000: data <= 18'h3ff55; 
        10'b0010110001: data <= 18'h3fedd; 
        10'b0010110010: data <= 18'h0009f; 
        10'b0010110011: data <= 18'h3ffe7; 
        10'b0010110100: data <= 18'h001b1; 
        10'b0010110101: data <= 18'h0017f; 
        10'b0010110110: data <= 18'h0016e; 
        10'b0010110111: data <= 18'h0021f; 
        10'b0010111000: data <= 18'h00296; 
        10'b0010111001: data <= 18'h003aa; 
        10'b0010111010: data <= 18'h00369; 
        10'b0010111011: data <= 18'h002e8; 
        10'b0010111100: data <= 18'h002ce; 
        10'b0010111101: data <= 18'h00333; 
        10'b0010111110: data <= 18'h001d0; 
        10'b0010111111: data <= 18'h000a6; 
        10'b0011000000: data <= 18'h3fe9c; 
        10'b0011000001: data <= 18'h3fe8e; 
        10'b0011000010: data <= 18'h3ff05; 
        10'b0011000011: data <= 18'h00025; 
        10'b0011000100: data <= 18'h00056; 
        10'b0011000101: data <= 18'h0000e; 
        10'b0011000110: data <= 18'h3ffee; 
        10'b0011000111: data <= 18'h3ff26; 
        10'b0011001000: data <= 18'h3feae; 
        10'b0011001001: data <= 18'h3ffe2; 
        10'b0011001010: data <= 18'h3ff78; 
        10'b0011001011: data <= 18'h00002; 
        10'b0011001100: data <= 18'h3ff61; 
        10'b0011001101: data <= 18'h3ffd1; 
        10'b0011001110: data <= 18'h0001e; 
        10'b0011001111: data <= 18'h00135; 
        10'b0011010000: data <= 18'h00284; 
        10'b0011010001: data <= 18'h00251; 
        10'b0011010010: data <= 18'h000f3; 
        10'b0011010011: data <= 18'h0017a; 
        10'b0011010100: data <= 18'h0021c; 
        10'b0011010101: data <= 18'h003ef; 
        10'b0011010110: data <= 18'h002e5; 
        10'b0011010111: data <= 18'h00289; 
        10'b0011011000: data <= 18'h00109; 
        10'b0011011001: data <= 18'h001fd; 
        10'b0011011010: data <= 18'h0022f; 
        10'b0011011011: data <= 18'h0011e; 
        10'b0011011100: data <= 18'h3ff27; 
        10'b0011011101: data <= 18'h3fe9c; 
        10'b0011011110: data <= 18'h3fec0; 
        10'b0011011111: data <= 18'h3ffec; 
        10'b0011100000: data <= 18'h00061; 
        10'b0011100001: data <= 18'h00023; 
        10'b0011100010: data <= 18'h3ffd7; 
        10'b0011100011: data <= 18'h3fffe; 
        10'b0011100100: data <= 18'h3ff08; 
        10'b0011100101: data <= 18'h3ff3f; 
        10'b0011100110: data <= 18'h3ff62; 
        10'b0011100111: data <= 18'h3ff3d; 
        10'b0011101000: data <= 18'h3ff99; 
        10'b0011101001: data <= 18'h3ff94; 
        10'b0011101010: data <= 18'h00131; 
        10'b0011101011: data <= 18'h00141; 
        10'b0011101100: data <= 18'h000a5; 
        10'b0011101101: data <= 18'h00045; 
        10'b0011101110: data <= 18'h00072; 
        10'b0011101111: data <= 18'h001c5; 
        10'b0011110000: data <= 18'h0052a; 
        10'b0011110001: data <= 18'h0041c; 
        10'b0011110010: data <= 18'h003d1; 
        10'b0011110011: data <= 18'h00133; 
        10'b0011110100: data <= 18'h00102; 
        10'b0011110101: data <= 18'h000ec; 
        10'b0011110110: data <= 18'h00243; 
        10'b0011110111: data <= 18'h003f1; 
        10'b0011111000: data <= 18'h3ff91; 
        10'b0011111001: data <= 18'h3feb0; 
        10'b0011111010: data <= 18'h3ffdf; 
        10'b0011111011: data <= 18'h3ff50; 
        10'b0011111100: data <= 18'h3ffe5; 
        10'b0011111101: data <= 18'h3ffef; 
        10'b0011111110: data <= 18'h0001e; 
        10'b0011111111: data <= 18'h00016; 
        10'b0100000000: data <= 18'h3fec8; 
        10'b0100000001: data <= 18'h3ff22; 
        10'b0100000010: data <= 18'h3fec1; 
        10'b0100000011: data <= 18'h3ff49; 
        10'b0100000100: data <= 18'h3ff4c; 
        10'b0100000101: data <= 18'h3ffa4; 
        10'b0100000110: data <= 18'h000dc; 
        10'b0100000111: data <= 18'h3ff44; 
        10'b0100001000: data <= 18'h0006d; 
        10'b0100001001: data <= 18'h0014b; 
        10'b0100001010: data <= 18'h00126; 
        10'b0100001011: data <= 18'h000fb; 
        10'b0100001100: data <= 18'h002d4; 
        10'b0100001101: data <= 18'h003c5; 
        10'b0100001110: data <= 18'h00455; 
        10'b0100001111: data <= 18'h00282; 
        10'b0100010000: data <= 18'h000c3; 
        10'b0100010001: data <= 18'h3ffdc; 
        10'b0100010010: data <= 18'h001dc; 
        10'b0100010011: data <= 18'h00403; 
        10'b0100010100: data <= 18'h0012b; 
        10'b0100010101: data <= 18'h3ff03; 
        10'b0100010110: data <= 18'h00004; 
        10'b0100010111: data <= 18'h3ffe1; 
        10'b0100011000: data <= 18'h3ff5e; 
        10'b0100011001: data <= 18'h0004f; 
        10'b0100011010: data <= 18'h3ff77; 
        10'b0100011011: data <= 18'h3ff08; 
        10'b0100011100: data <= 18'h3ff1c; 
        10'b0100011101: data <= 18'h3ff4c; 
        10'b0100011110: data <= 18'h3ff67; 
        10'b0100011111: data <= 18'h00014; 
        10'b0100100000: data <= 18'h00069; 
        10'b0100100001: data <= 18'h3ffe8; 
        10'b0100100010: data <= 18'h3ff52; 
        10'b0100100011: data <= 18'h00039; 
        10'b0100100100: data <= 18'h00047; 
        10'b0100100101: data <= 18'h3ffd7; 
        10'b0100100110: data <= 18'h3fea4; 
        10'b0100100111: data <= 18'h3fda9; 
        10'b0100101000: data <= 18'h3fe98; 
        10'b0100101001: data <= 18'h0015b; 
        10'b0100101010: data <= 18'h00372; 
        10'b0100101011: data <= 18'h00392; 
        10'b0100101100: data <= 18'h00329; 
        10'b0100101101: data <= 18'h0024a; 
        10'b0100101110: data <= 18'h00365; 
        10'b0100101111: data <= 18'h004a4; 
        10'b0100110000: data <= 18'h00236; 
        10'b0100110001: data <= 18'h3ff17; 
        10'b0100110010: data <= 18'h3ff16; 
        10'b0100110011: data <= 18'h3ff4d; 
        10'b0100110100: data <= 18'h3ff87; 
        10'b0100110101: data <= 18'h3ff5e; 
        10'b0100110110: data <= 18'h00044; 
        10'b0100110111: data <= 18'h3ffce; 
        10'b0100111000: data <= 18'h3fe42; 
        10'b0100111001: data <= 18'h3ffa1; 
        10'b0100111010: data <= 18'h00046; 
        10'b0100111011: data <= 18'h00150; 
        10'b0100111100: data <= 18'h000fd; 
        10'b0100111101: data <= 18'h3ff9f; 
        10'b0100111110: data <= 18'h00058; 
        10'b0100111111: data <= 18'h00009; 
        10'b0101000000: data <= 18'h000ae; 
        10'b0101000001: data <= 18'h3ff8a; 
        10'b0101000010: data <= 18'h3fc4f; 
        10'b0101000011: data <= 18'h3f929; 
        10'b0101000100: data <= 18'h3f991; 
        10'b0101000101: data <= 18'h3fd7c; 
        10'b0101000110: data <= 18'h3ffaa; 
        10'b0101000111: data <= 18'h001d1; 
        10'b0101001000: data <= 18'h002e8; 
        10'b0101001001: data <= 18'h002b1; 
        10'b0101001010: data <= 18'h003ab; 
        10'b0101001011: data <= 18'h0042a; 
        10'b0101001100: data <= 18'h002fe; 
        10'b0101001101: data <= 18'h3ff6d; 
        10'b0101001110: data <= 18'h3fff6; 
        10'b0101001111: data <= 18'h3ff42; 
        10'b0101010000: data <= 18'h3ff80; 
        10'b0101010001: data <= 18'h3ffd7; 
        10'b0101010010: data <= 18'h3ffc6; 
        10'b0101010011: data <= 18'h3ffcf; 
        10'b0101010100: data <= 18'h3ff05; 
        10'b0101010101: data <= 18'h00028; 
        10'b0101010110: data <= 18'h0016f; 
        10'b0101010111: data <= 18'h0017f; 
        10'b0101011000: data <= 18'h000b9; 
        10'b0101011001: data <= 18'h3ffcd; 
        10'b0101011010: data <= 18'h00107; 
        10'b0101011011: data <= 18'h000ba; 
        10'b0101011100: data <= 18'h00158; 
        10'b0101011101: data <= 18'h3fee5; 
        10'b0101011110: data <= 18'h3f8c2; 
        10'b0101011111: data <= 18'h3f707; 
        10'b0101100000: data <= 18'h3f711; 
        10'b0101100001: data <= 18'h3fb1e; 
        10'b0101100010: data <= 18'h3ff23; 
        10'b0101100011: data <= 18'h3ffa4; 
        10'b0101100100: data <= 18'h00070; 
        10'b0101100101: data <= 18'h00140; 
        10'b0101100110: data <= 18'h004c2; 
        10'b0101100111: data <= 18'h0045a; 
        10'b0101101000: data <= 18'h00306; 
        10'b0101101001: data <= 18'h0001c; 
        10'b0101101010: data <= 18'h3ff86; 
        10'b0101101011: data <= 18'h3ff85; 
        10'b0101101100: data <= 18'h3ff4a; 
        10'b0101101101: data <= 18'h3fffc; 
        10'b0101101110: data <= 18'h00040; 
        10'b0101101111: data <= 18'h3ff52; 
        10'b0101110000: data <= 18'h3ffbd; 
        10'b0101110001: data <= 18'h000e3; 
        10'b0101110010: data <= 18'h001bc; 
        10'b0101110011: data <= 18'h0023e; 
        10'b0101110100: data <= 18'h001b2; 
        10'b0101110101: data <= 18'h00130; 
        10'b0101110110: data <= 18'h0019f; 
        10'b0101110111: data <= 18'h00142; 
        10'b0101111000: data <= 18'h000e8; 
        10'b0101111001: data <= 18'h3fb97; 
        10'b0101111010: data <= 18'h3f8be; 
        10'b0101111011: data <= 18'h3f6c7; 
        10'b0101111100: data <= 18'h3f86e; 
        10'b0101111101: data <= 18'h3fc3e; 
        10'b0101111110: data <= 18'h3fe2a; 
        10'b0101111111: data <= 18'h3fd89; 
        10'b0110000000: data <= 18'h3fe1d; 
        10'b0110000001: data <= 18'h000d4; 
        10'b0110000010: data <= 18'h0031f; 
        10'b0110000011: data <= 18'h004e7; 
        10'b0110000100: data <= 18'h002c8; 
        10'b0110000101: data <= 18'h00073; 
        10'b0110000110: data <= 18'h00001; 
        10'b0110000111: data <= 18'h00045; 
        10'b0110001000: data <= 18'h3ffe6; 
        10'b0110001001: data <= 18'h00037; 
        10'b0110001010: data <= 18'h3ff75; 
        10'b0110001011: data <= 18'h3ff9b; 
        10'b0110001100: data <= 18'h3ff28; 
        10'b0110001101: data <= 18'h0024b; 
        10'b0110001110: data <= 18'h002fa; 
        10'b0110001111: data <= 18'h0039e; 
        10'b0110010000: data <= 18'h001bc; 
        10'b0110010001: data <= 18'h00216; 
        10'b0110010010: data <= 18'h00311; 
        10'b0110010011: data <= 18'h001c3; 
        10'b0110010100: data <= 18'h0006e; 
        10'b0110010101: data <= 18'h3fc29; 
        10'b0110010110: data <= 18'h3f771; 
        10'b0110010111: data <= 18'h3f6c1; 
        10'b0110011000: data <= 18'h3f8a5; 
        10'b0110011001: data <= 18'h3fbfa; 
        10'b0110011010: data <= 18'h3fe3a; 
        10'b0110011011: data <= 18'h3fddc; 
        10'b0110011100: data <= 18'h00031; 
        10'b0110011101: data <= 18'h001be; 
        10'b0110011110: data <= 18'h00215; 
        10'b0110011111: data <= 18'h004f4; 
        10'b0110100000: data <= 18'h00294; 
        10'b0110100001: data <= 18'h3ff7b; 
        10'b0110100010: data <= 18'h3ffbe; 
        10'b0110100011: data <= 18'h3ff72; 
        10'b0110100100: data <= 18'h0004a; 
        10'b0110100101: data <= 18'h00029; 
        10'b0110100110: data <= 18'h3ff87; 
        10'b0110100111: data <= 18'h3ffe4; 
        10'b0110101000: data <= 18'h3fff6; 
        10'b0110101001: data <= 18'h0033d; 
        10'b0110101010: data <= 18'h00259; 
        10'b0110101011: data <= 18'h0033c; 
        10'b0110101100: data <= 18'h0023b; 
        10'b0110101101: data <= 18'h002f6; 
        10'b0110101110: data <= 18'h003be; 
        10'b0110101111: data <= 18'h00108; 
        10'b0110110000: data <= 18'h3fd2f; 
        10'b0110110001: data <= 18'h3f8d2; 
        10'b0110110010: data <= 18'h3f669; 
        10'b0110110011: data <= 18'h3f6df; 
        10'b0110110100: data <= 18'h3f9d5; 
        10'b0110110101: data <= 18'h3fcfd; 
        10'b0110110110: data <= 18'h3fee0; 
        10'b0110110111: data <= 18'h3feea; 
        10'b0110111000: data <= 18'h000f0; 
        10'b0110111001: data <= 18'h000d2; 
        10'b0110111010: data <= 18'h00325; 
        10'b0110111011: data <= 18'h003b2; 
        10'b0110111100: data <= 18'h001ea; 
        10'b0110111101: data <= 18'h3ffd0; 
        10'b0110111110: data <= 18'h0000e; 
        10'b0110111111: data <= 18'h3ff7f; 
        10'b0111000000: data <= 18'h00015; 
        10'b0111000001: data <= 18'h0005d; 
        10'b0111000010: data <= 18'h3ff44; 
        10'b0111000011: data <= 18'h3ff9b; 
        10'b0111000100: data <= 18'h0008c; 
        10'b0111000101: data <= 18'h002f0; 
        10'b0111000110: data <= 18'h003a6; 
        10'b0111000111: data <= 18'h002d3; 
        10'b0111001000: data <= 18'h001f6; 
        10'b0111001001: data <= 18'h001fa; 
        10'b0111001010: data <= 18'h00355; 
        10'b0111001011: data <= 18'h3ff90; 
        10'b0111001100: data <= 18'h3fa87; 
        10'b0111001101: data <= 18'h3f67c; 
        10'b0111001110: data <= 18'h3f6bb; 
        10'b0111001111: data <= 18'h3f8a6; 
        10'b0111010000: data <= 18'h3fc10; 
        10'b0111010001: data <= 18'h3fe29; 
        10'b0111010010: data <= 18'h3fffa; 
        10'b0111010011: data <= 18'h0009a; 
        10'b0111010100: data <= 18'h00163; 
        10'b0111010101: data <= 18'h0020f; 
        10'b0111010110: data <= 18'h002d5; 
        10'b0111010111: data <= 18'h002b4; 
        10'b0111011000: data <= 18'h00107; 
        10'b0111011001: data <= 18'h0000d; 
        10'b0111011010: data <= 18'h3ffaa; 
        10'b0111011011: data <= 18'h3ff8c; 
        10'b0111011100: data <= 18'h3ffbd; 
        10'b0111011101: data <= 18'h00017; 
        10'b0111011110: data <= 18'h3ff61; 
        10'b0111011111: data <= 18'h3fecc; 
        10'b0111100000: data <= 18'h0001a; 
        10'b0111100001: data <= 18'h00216; 
        10'b0111100010: data <= 18'h0029e; 
        10'b0111100011: data <= 18'h0028b; 
        10'b0111100100: data <= 18'h000cb; 
        10'b0111100101: data <= 18'h0020b; 
        10'b0111100110: data <= 18'h0033b; 
        10'b0111100111: data <= 18'h3ff81; 
        10'b0111101000: data <= 18'h3f972; 
        10'b0111101001: data <= 18'h3f69d; 
        10'b0111101010: data <= 18'h3f7bc; 
        10'b0111101011: data <= 18'h3fb13; 
        10'b0111101100: data <= 18'h3ff5a; 
        10'b0111101101: data <= 18'h00142; 
        10'b0111101110: data <= 18'h001cf; 
        10'b0111101111: data <= 18'h001ab; 
        10'b0111110000: data <= 18'h00221; 
        10'b0111110001: data <= 18'h0019f; 
        10'b0111110010: data <= 18'h00148; 
        10'b0111110011: data <= 18'h00175; 
        10'b0111110100: data <= 18'h3ffec; 
        10'b0111110101: data <= 18'h3ffc9; 
        10'b0111110110: data <= 18'h0001d; 
        10'b0111110111: data <= 18'h3ff7e; 
        10'b0111111000: data <= 18'h3ffa6; 
        10'b0111111001: data <= 18'h0001d; 
        10'b0111111010: data <= 18'h3ffc1; 
        10'b0111111011: data <= 18'h3ff8a; 
        10'b0111111100: data <= 18'h3ffbf; 
        10'b0111111101: data <= 18'h00155; 
        10'b0111111110: data <= 18'h002b7; 
        10'b0111111111: data <= 18'h00191; 
        10'b1000000000: data <= 18'h000f6; 
        10'b1000000001: data <= 18'h002b3; 
        10'b1000000010: data <= 18'h0052d; 
        10'b1000000011: data <= 18'h00034; 
        10'b1000000100: data <= 18'h3fbd3; 
        10'b1000000101: data <= 18'h3f943; 
        10'b1000000110: data <= 18'h3fb4d; 
        10'b1000000111: data <= 18'h3fe91; 
        10'b1000001000: data <= 18'h00184; 
        10'b1000001001: data <= 18'h0019e; 
        10'b1000001010: data <= 18'h001b2; 
        10'b1000001011: data <= 18'h000e2; 
        10'b1000001100: data <= 18'h00070; 
        10'b1000001101: data <= 18'h000bc; 
        10'b1000001110: data <= 18'h00169; 
        10'b1000001111: data <= 18'h000e1; 
        10'b1000010000: data <= 18'h3ffe4; 
        10'b1000010001: data <= 18'h3ff91; 
        10'b1000010010: data <= 18'h0000d; 
        10'b1000010011: data <= 18'h3ffc2; 
        10'b1000010100: data <= 18'h3ffc9; 
        10'b1000010101: data <= 18'h3ffb3; 
        10'b1000010110: data <= 18'h3ffbb; 
        10'b1000010111: data <= 18'h3fed4; 
        10'b1000011000: data <= 18'h00081; 
        10'b1000011001: data <= 18'h00176; 
        10'b1000011010: data <= 18'h0037c; 
        10'b1000011011: data <= 18'h0032b; 
        10'b1000011100: data <= 18'h0027a; 
        10'b1000011101: data <= 18'h0034a; 
        10'b1000011110: data <= 18'h00530; 
        10'b1000011111: data <= 18'h003a6; 
        10'b1000100000: data <= 18'h000c5; 
        10'b1000100001: data <= 18'h3fe53; 
        10'b1000100010: data <= 18'h3ff44; 
        10'b1000100011: data <= 18'h3ff88; 
        10'b1000100100: data <= 18'h000cb; 
        10'b1000100101: data <= 18'h3ffa3; 
        10'b1000100110: data <= 18'h3ff54; 
        10'b1000100111: data <= 18'h3ff97; 
        10'b1000101000: data <= 18'h000d1; 
        10'b1000101001: data <= 18'h000be; 
        10'b1000101010: data <= 18'h00175; 
        10'b1000101011: data <= 18'h3ffcf; 
        10'b1000101100: data <= 18'h00035; 
        10'b1000101101: data <= 18'h3ffae; 
        10'b1000101110: data <= 18'h3ff40; 
        10'b1000101111: data <= 18'h00043; 
        10'b1000110000: data <= 18'h00041; 
        10'b1000110001: data <= 18'h00057; 
        10'b1000110010: data <= 18'h3ffc2; 
        10'b1000110011: data <= 18'h3ff71; 
        10'b1000110100: data <= 18'h3ffab; 
        10'b1000110101: data <= 18'h0017f; 
        10'b1000110110: data <= 18'h002cd; 
        10'b1000110111: data <= 18'h00210; 
        10'b1000111000: data <= 18'h0028f; 
        10'b1000111001: data <= 18'h00324; 
        10'b1000111010: data <= 18'h004e6; 
        10'b1000111011: data <= 18'h004e4; 
        10'b1000111100: data <= 18'h00273; 
        10'b1000111101: data <= 18'h000bf; 
        10'b1000111110: data <= 18'h3ff7e; 
        10'b1000111111: data <= 18'h0005a; 
        10'b1001000000: data <= 18'h00055; 
        10'b1001000001: data <= 18'h3ff49; 
        10'b1001000010: data <= 18'h3ff75; 
        10'b1001000011: data <= 18'h3ff3d; 
        10'b1001000100: data <= 18'h00068; 
        10'b1001000101: data <= 18'h00080; 
        10'b1001000110: data <= 18'h000c5; 
        10'b1001000111: data <= 18'h00044; 
        10'b1001001000: data <= 18'h3ff92; 
        10'b1001001001: data <= 18'h3ffe7; 
        10'b1001001010: data <= 18'h3ff65; 
        10'b1001001011: data <= 18'h3ffaf; 
        10'b1001001100: data <= 18'h3ff8d; 
        10'b1001001101: data <= 18'h3ff56; 
        10'b1001001110: data <= 18'h3ffc3; 
        10'b1001001111: data <= 18'h3ff90; 
        10'b1001010000: data <= 18'h3ffb8; 
        10'b1001010001: data <= 18'h00063; 
        10'b1001010010: data <= 18'h001bb; 
        10'b1001010011: data <= 18'h002d1; 
        10'b1001010100: data <= 18'h001fa; 
        10'b1001010101: data <= 18'h00225; 
        10'b1001010110: data <= 18'h00431; 
        10'b1001010111: data <= 18'h004bd; 
        10'b1001011000: data <= 18'h00325; 
        10'b1001011001: data <= 18'h00130; 
        10'b1001011010: data <= 18'h00071; 
        10'b1001011011: data <= 18'h00018; 
        10'b1001011100: data <= 18'h3ffec; 
        10'b1001011101: data <= 18'h3feb4; 
        10'b1001011110: data <= 18'h3ff03; 
        10'b1001011111: data <= 18'h3ff6e; 
        10'b1001100000: data <= 18'h0007f; 
        10'b1001100001: data <= 18'h3fff7; 
        10'b1001100010: data <= 18'h3ff6a; 
        10'b1001100011: data <= 18'h3ff0f; 
        10'b1001100100: data <= 18'h3ffc5; 
        10'b1001100101: data <= 18'h3ffb1; 
        10'b1001100110: data <= 18'h3ff8b; 
        10'b1001100111: data <= 18'h3ff9c; 
        10'b1001101000: data <= 18'h3ff71; 
        10'b1001101001: data <= 18'h00009; 
        10'b1001101010: data <= 18'h0000d; 
        10'b1001101011: data <= 18'h3ffab; 
        10'b1001101100: data <= 18'h3ff69; 
        10'b1001101101: data <= 18'h00038; 
        10'b1001101110: data <= 18'h00142; 
        10'b1001101111: data <= 18'h00118; 
        10'b1001110000: data <= 18'h00329; 
        10'b1001110001: data <= 18'h00292; 
        10'b1001110010: data <= 18'h002d5; 
        10'b1001110011: data <= 18'h0035e; 
        10'b1001110100: data <= 18'h002df; 
        10'b1001110101: data <= 18'h003b1; 
        10'b1001110110: data <= 18'h00199; 
        10'b1001110111: data <= 18'h001a3; 
        10'b1001111000: data <= 18'h000e5; 
        10'b1001111001: data <= 18'h3ff3d; 
        10'b1001111010: data <= 18'h3ff65; 
        10'b1001111011: data <= 18'h3fff5; 
        10'b1001111100: data <= 18'h3ff25; 
        10'b1001111101: data <= 18'h3ff1b; 
        10'b1001111110: data <= 18'h3ff92; 
        10'b1001111111: data <= 18'h3ff89; 
        10'b1010000000: data <= 18'h3ffd5; 
        10'b1010000001: data <= 18'h3ffb6; 
        10'b1010000010: data <= 18'h3ffa1; 
        10'b1010000011: data <= 18'h3ffce; 
        10'b1010000100: data <= 18'h3ff70; 
        10'b1010000101: data <= 18'h3ffd9; 
        10'b1010000110: data <= 18'h3fffc; 
        10'b1010000111: data <= 18'h3ff52; 
        10'b1010001000: data <= 18'h3ff4e; 
        10'b1010001001: data <= 18'h3ffcd; 
        10'b1010001010: data <= 18'h3ffeb; 
        10'b1010001011: data <= 18'h000e0; 
        10'b1010001100: data <= 18'h0013c; 
        10'b1010001101: data <= 18'h002ee; 
        10'b1010001110: data <= 18'h00381; 
        10'b1010001111: data <= 18'h00449; 
        10'b1010010000: data <= 18'h0043e; 
        10'b1010010001: data <= 18'h0028b; 
        10'b1010010010: data <= 18'h00212; 
        10'b1010010011: data <= 18'h00125; 
        10'b1010010100: data <= 18'h0007c; 
        10'b1010010101: data <= 18'h3fff4; 
        10'b1010010110: data <= 18'h3fe63; 
        10'b1010010111: data <= 18'h3fdfa; 
        10'b1010011000: data <= 18'h3fe6e; 
        10'b1010011001: data <= 18'h3ff3a; 
        10'b1010011010: data <= 18'h3ff5f; 
        10'b1010011011: data <= 18'h3ffeb; 
        10'b1010011100: data <= 18'h3ffc3; 
        10'b1010011101: data <= 18'h00032; 
        10'b1010011110: data <= 18'h3ffaa; 
        10'b1010011111: data <= 18'h3ff4b; 
        10'b1010100000: data <= 18'h3ffb0; 
        10'b1010100001: data <= 18'h3ffdd; 
        10'b1010100010: data <= 18'h3ff4e; 
        10'b1010100011: data <= 18'h3fff9; 
        10'b1010100100: data <= 18'h3ffcf; 
        10'b1010100101: data <= 18'h3ffd2; 
        10'b1010100110: data <= 18'h3ff2a; 
        10'b1010100111: data <= 18'h3fee3; 
        10'b1010101000: data <= 18'h3ff61; 
        10'b1010101001: data <= 18'h3ff72; 
        10'b1010101010: data <= 18'h000a6; 
        10'b1010101011: data <= 18'h0007d; 
        10'b1010101100: data <= 18'h0012f; 
        10'b1010101101: data <= 18'h001bc; 
        10'b1010101110: data <= 18'h000ea; 
        10'b1010101111: data <= 18'h3ff4e; 
        10'b1010110000: data <= 18'h3feeb; 
        10'b1010110001: data <= 18'h3feb5; 
        10'b1010110010: data <= 18'h3fee6; 
        10'b1010110011: data <= 18'h3fe75; 
        10'b1010110100: data <= 18'h3fe87; 
        10'b1010110101: data <= 18'h3fe9c; 
        10'b1010110110: data <= 18'h3ffba; 
        10'b1010110111: data <= 18'h3ffa3; 
        10'b1010111000: data <= 18'h3ff6a; 
        10'b1010111001: data <= 18'h3ff92; 
        10'b1010111010: data <= 18'h00009; 
        10'b1010111011: data <= 18'h3ff7e; 
        10'b1010111100: data <= 18'h3ff93; 
        10'b1010111101: data <= 18'h00066; 
        10'b1010111110: data <= 18'h3ffca; 
        10'b1010111111: data <= 18'h00055; 
        10'b1011000000: data <= 18'h00060; 
        10'b1011000001: data <= 18'h3fffb; 
        10'b1011000010: data <= 18'h3ff40; 
        10'b1011000011: data <= 18'h3ffac; 
        10'b1011000100: data <= 18'h3fe89; 
        10'b1011000101: data <= 18'h3fe9d; 
        10'b1011000110: data <= 18'h3fe47; 
        10'b1011000111: data <= 18'h3fdc3; 
        10'b1011001000: data <= 18'h3fd71; 
        10'b1011001001: data <= 18'h3fdac; 
        10'b1011001010: data <= 18'h3fd4a; 
        10'b1011001011: data <= 18'h3fd8e; 
        10'b1011001100: data <= 18'h3fdb0; 
        10'b1011001101: data <= 18'h3fe9c; 
        10'b1011001110: data <= 18'h3fed9; 
        10'b1011001111: data <= 18'h3ff06; 
        10'b1011010000: data <= 18'h3feeb; 
        10'b1011010001: data <= 18'h3ff01; 
        10'b1011010010: data <= 18'h3ffab; 
        10'b1011010011: data <= 18'h00060; 
        10'b1011010100: data <= 18'h0002f; 
        10'b1011010101: data <= 18'h3ffbc; 
        10'b1011010110: data <= 18'h3ffa5; 
        10'b1011010111: data <= 18'h3ffdd; 
        10'b1011011000: data <= 18'h00051; 
        10'b1011011001: data <= 18'h00048; 
        10'b1011011010: data <= 18'h3ffb7; 
        10'b1011011011: data <= 18'h00005; 
        10'b1011011100: data <= 18'h3ff9c; 
        10'b1011011101: data <= 18'h3ffaf; 
        10'b1011011110: data <= 18'h3ff53; 
        10'b1011011111: data <= 18'h00022; 
        10'b1011100000: data <= 18'h3ffa4; 
        10'b1011100001: data <= 18'h3fec6; 
        10'b1011100010: data <= 18'h3fec5; 
        10'b1011100011: data <= 18'h3fee3; 
        10'b1011100100: data <= 18'h3ff8d; 
        10'b1011100101: data <= 18'h3fee3; 
        10'b1011100110: data <= 18'h3fef2; 
        10'b1011100111: data <= 18'h3ff9b; 
        10'b1011101000: data <= 18'h3fee0; 
        10'b1011101001: data <= 18'h3ff16; 
        10'b1011101010: data <= 18'h3ff52; 
        10'b1011101011: data <= 18'h3ff24; 
        10'b1011101100: data <= 18'h3ff93; 
        10'b1011101101: data <= 18'h3fef8; 
        10'b1011101110: data <= 18'h3ff21; 
        10'b1011101111: data <= 18'h00057; 
        10'b1011110000: data <= 18'h3ff78; 
        10'b1011110001: data <= 18'h00019; 
        10'b1011110010: data <= 18'h00048; 
        10'b1011110011: data <= 18'h3fff0; 
        10'b1011110100: data <= 18'h3ff6c; 
        10'b1011110101: data <= 18'h0003c; 
        10'b1011110110: data <= 18'h3ffe7; 
        10'b1011110111: data <= 18'h3ffb0; 
        10'b1011111000: data <= 18'h0004c; 
        10'b1011111001: data <= 18'h0000f; 
        10'b1011111010: data <= 18'h0001b; 
        10'b1011111011: data <= 18'h3ff4a; 
        10'b1011111100: data <= 18'h00059; 
        10'b1011111101: data <= 18'h00057; 
        10'b1011111110: data <= 18'h0001e; 
        10'b1011111111: data <= 18'h0003f; 
        10'b1100000000: data <= 18'h3ffd5; 
        10'b1100000001: data <= 18'h3ff94; 
        10'b1100000010: data <= 18'h0003b; 
        10'b1100000011: data <= 18'h3ff64; 
        10'b1100000100: data <= 18'h3ffc6; 
        10'b1100000101: data <= 18'h3ff92; 
        10'b1100000110: data <= 18'h3ffe5; 
        10'b1100000111: data <= 18'h3ff9f; 
        10'b1100001000: data <= 18'h3ff46; 
        10'b1100001001: data <= 18'h3ff5a; 
        10'b1100001010: data <= 18'h3ff13; 
        10'b1100001011: data <= 18'h3ffc9; 
        10'b1100001100: data <= 18'h00026; 
        10'b1100001101: data <= 18'h3ff6a; 
        10'b1100001110: data <= 18'h3ff43; 
        10'b1100001111: data <= 18'h00032; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 13) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 19'h7fef7; 
        10'b0000000001: data <= 19'h00098; 
        10'b0000000010: data <= 19'h7ffae; 
        10'b0000000011: data <= 19'h7ffd9; 
        10'b0000000100: data <= 19'h000b2; 
        10'b0000000101: data <= 19'h7ffee; 
        10'b0000000110: data <= 19'h7ff58; 
        10'b0000000111: data <= 19'h7ff4d; 
        10'b0000001000: data <= 19'h7ffd7; 
        10'b0000001001: data <= 19'h7ffa7; 
        10'b0000001010: data <= 19'h000c6; 
        10'b0000001011: data <= 19'h7fff0; 
        10'b0000001100: data <= 19'h0005b; 
        10'b0000001101: data <= 19'h7fefe; 
        10'b0000001110: data <= 19'h7fff2; 
        10'b0000001111: data <= 19'h7fe9d; 
        10'b0000010000: data <= 19'h7fed9; 
        10'b0000010001: data <= 19'h7ffb1; 
        10'b0000010010: data <= 19'h7fed0; 
        10'b0000010011: data <= 19'h000c5; 
        10'b0000010100: data <= 19'h7fed7; 
        10'b0000010101: data <= 19'h7ffa1; 
        10'b0000010110: data <= 19'h7fec0; 
        10'b0000010111: data <= 19'h7ffe0; 
        10'b0000011000: data <= 19'h00063; 
        10'b0000011001: data <= 19'h7ffb9; 
        10'b0000011010: data <= 19'h7fff1; 
        10'b0000011011: data <= 19'h7fff6; 
        10'b0000011100: data <= 19'h00070; 
        10'b0000011101: data <= 19'h0008a; 
        10'b0000011110: data <= 19'h0002d; 
        10'b0000011111: data <= 19'h7fec9; 
        10'b0000100000: data <= 19'h7feb9; 
        10'b0000100001: data <= 19'h00011; 
        10'b0000100010: data <= 19'h7fefd; 
        10'b0000100011: data <= 19'h7ffb8; 
        10'b0000100100: data <= 19'h7ff38; 
        10'b0000100101: data <= 19'h7fe92; 
        10'b0000100110: data <= 19'h7ff17; 
        10'b0000100111: data <= 19'h00013; 
        10'b0000101000: data <= 19'h000de; 
        10'b0000101001: data <= 19'h7fecf; 
        10'b0000101010: data <= 19'h7ff5b; 
        10'b0000101011: data <= 19'h00060; 
        10'b0000101100: data <= 19'h7ff03; 
        10'b0000101101: data <= 19'h7fea7; 
        10'b0000101110: data <= 19'h00041; 
        10'b0000101111: data <= 19'h0009a; 
        10'b0000110000: data <= 19'h7fef7; 
        10'b0000110001: data <= 19'h00048; 
        10'b0000110010: data <= 19'h7ff1f; 
        10'b0000110011: data <= 19'h7fee3; 
        10'b0000110100: data <= 19'h7ffc8; 
        10'b0000110101: data <= 19'h00013; 
        10'b0000110110: data <= 19'h7ffa6; 
        10'b0000110111: data <= 19'h000c0; 
        10'b0000111000: data <= 19'h7feb4; 
        10'b0000111001: data <= 19'h7ff34; 
        10'b0000111010: data <= 19'h7ff21; 
        10'b0000111011: data <= 19'h0005e; 
        10'b0000111100: data <= 19'h0001a; 
        10'b0000111101: data <= 19'h7feaa; 
        10'b0000111110: data <= 19'h7ffae; 
        10'b0000111111: data <= 19'h000b7; 
        10'b0001000000: data <= 19'h7ff91; 
        10'b0001000001: data <= 19'h7ff0a; 
        10'b0001000010: data <= 19'h7ff14; 
        10'b0001000011: data <= 19'h7fe6b; 
        10'b0001000100: data <= 19'h7fe51; 
        10'b0001000101: data <= 19'h7ff6b; 
        10'b0001000110: data <= 19'h7fe42; 
        10'b0001000111: data <= 19'h7fdc4; 
        10'b0001001000: data <= 19'h7fe5e; 
        10'b0001001001: data <= 19'h7ff93; 
        10'b0001001010: data <= 19'h7fe9d; 
        10'b0001001011: data <= 19'h7fe37; 
        10'b0001001100: data <= 19'h7ffb1; 
        10'b0001001101: data <= 19'h0008a; 
        10'b0001001110: data <= 19'h00019; 
        10'b0001001111: data <= 19'h7ff03; 
        10'b0001010000: data <= 19'h000ac; 
        10'b0001010001: data <= 19'h7fe94; 
        10'b0001010010: data <= 19'h7ffa8; 
        10'b0001010011: data <= 19'h00053; 
        10'b0001010100: data <= 19'h7feab; 
        10'b0001010101: data <= 19'h7ffb0; 
        10'b0001010110: data <= 19'h000c0; 
        10'b0001010111: data <= 19'h7feb5; 
        10'b0001011000: data <= 19'h7ff12; 
        10'b0001011001: data <= 19'h0009c; 
        10'b0001011010: data <= 19'h0003f; 
        10'b0001011011: data <= 19'h00007; 
        10'b0001011100: data <= 19'h00019; 
        10'b0001011101: data <= 19'h7ffa9; 
        10'b0001011110: data <= 19'h7ff8d; 
        10'b0001011111: data <= 19'h7fe3d; 
        10'b0001100000: data <= 19'h7fd96; 
        10'b0001100001: data <= 19'h7fea2; 
        10'b0001100010: data <= 19'h7fe1d; 
        10'b0001100011: data <= 19'h7fddd; 
        10'b0001100100: data <= 19'h0005b; 
        10'b0001100101: data <= 19'h0002c; 
        10'b0001100110: data <= 19'h7fd9e; 
        10'b0001100111: data <= 19'h7fdf6; 
        10'b0001101000: data <= 19'h7fd15; 
        10'b0001101001: data <= 19'h7fded; 
        10'b0001101010: data <= 19'h7fd80; 
        10'b0001101011: data <= 19'h7fe43; 
        10'b0001101100: data <= 19'h7fecc; 
        10'b0001101101: data <= 19'h00075; 
        10'b0001101110: data <= 19'h00071; 
        10'b0001101111: data <= 19'h7ff50; 
        10'b0001110000: data <= 19'h0002c; 
        10'b0001110001: data <= 19'h7fea6; 
        10'b0001110010: data <= 19'h7ff0d; 
        10'b0001110011: data <= 19'h7feae; 
        10'b0001110100: data <= 19'h7fe82; 
        10'b0001110101: data <= 19'h7ffce; 
        10'b0001110110: data <= 19'h7ff98; 
        10'b0001110111: data <= 19'h7feaa; 
        10'b0001111000: data <= 19'h7ff8d; 
        10'b0001111001: data <= 19'h7ffb6; 
        10'b0001111010: data <= 19'h7fdd6; 
        10'b0001111011: data <= 19'h7fddc; 
        10'b0001111100: data <= 19'h7fde5; 
        10'b0001111101: data <= 19'h7fdfd; 
        10'b0001111110: data <= 19'h7ff74; 
        10'b0001111111: data <= 19'h7ffc9; 
        10'b0010000000: data <= 19'h7fe58; 
        10'b0010000001: data <= 19'h7fe72; 
        10'b0010000010: data <= 19'h7fe65; 
        10'b0010000011: data <= 19'h7fdc3; 
        10'b0010000100: data <= 19'h7ff17; 
        10'b0010000101: data <= 19'h7fd1e; 
        10'b0010000110: data <= 19'h7fee1; 
        10'b0010000111: data <= 19'h7ffd8; 
        10'b0010001000: data <= 19'h7febf; 
        10'b0010001001: data <= 19'h7ff6f; 
        10'b0010001010: data <= 19'h7ff43; 
        10'b0010001011: data <= 19'h7ffe1; 
        10'b0010001100: data <= 19'h0005b; 
        10'b0010001101: data <= 19'h7ff5d; 
        10'b0010001110: data <= 19'h7fff8; 
        10'b0010001111: data <= 19'h7fed1; 
        10'b0010010000: data <= 19'h7ffae; 
        10'b0010010001: data <= 19'h7ff6c; 
        10'b0010010010: data <= 19'h7ff94; 
        10'b0010010011: data <= 19'h7ff1b; 
        10'b0010010100: data <= 19'h7ff98; 
        10'b0010010101: data <= 19'h7fe62; 
        10'b0010010110: data <= 19'h7ff46; 
        10'b0010010111: data <= 19'h0007a; 
        10'b0010011000: data <= 19'h001e4; 
        10'b0010011001: data <= 19'h00415; 
        10'b0010011010: data <= 19'h004ef; 
        10'b0010011011: data <= 19'h004e1; 
        10'b0010011100: data <= 19'h0057d; 
        10'b0010011101: data <= 19'h005e8; 
        10'b0010011110: data <= 19'h0063f; 
        10'b0010011111: data <= 19'h00234; 
        10'b0010100000: data <= 19'h00064; 
        10'b0010100001: data <= 19'h00104; 
        10'b0010100010: data <= 19'h7ff7f; 
        10'b0010100011: data <= 19'h7ffee; 
        10'b0010100100: data <= 19'h7fd55; 
        10'b0010100101: data <= 19'h7fe10; 
        10'b0010100110: data <= 19'h7ffdd; 
        10'b0010100111: data <= 19'h7fef8; 
        10'b0010101000: data <= 19'h7ff77; 
        10'b0010101001: data <= 19'h7ffc0; 
        10'b0010101010: data <= 19'h00025; 
        10'b0010101011: data <= 19'h7ff8f; 
        10'b0010101100: data <= 19'h00005; 
        10'b0010101101: data <= 19'h00011; 
        10'b0010101110: data <= 19'h00027; 
        10'b0010101111: data <= 19'h7fff1; 
        10'b0010110000: data <= 19'h7fea9; 
        10'b0010110001: data <= 19'h7fdba; 
        10'b0010110010: data <= 19'h0013f; 
        10'b0010110011: data <= 19'h7ffce; 
        10'b0010110100: data <= 19'h00362; 
        10'b0010110101: data <= 19'h002ff; 
        10'b0010110110: data <= 19'h002dc; 
        10'b0010110111: data <= 19'h0043e; 
        10'b0010111000: data <= 19'h0052c; 
        10'b0010111001: data <= 19'h00754; 
        10'b0010111010: data <= 19'h006d2; 
        10'b0010111011: data <= 19'h005d1; 
        10'b0010111100: data <= 19'h0059c; 
        10'b0010111101: data <= 19'h00667; 
        10'b0010111110: data <= 19'h003a1; 
        10'b0010111111: data <= 19'h0014c; 
        10'b0011000000: data <= 19'h7fd38; 
        10'b0011000001: data <= 19'h7fd1b; 
        10'b0011000010: data <= 19'h7fe0b; 
        10'b0011000011: data <= 19'h0004b; 
        10'b0011000100: data <= 19'h000ab; 
        10'b0011000101: data <= 19'h0001c; 
        10'b0011000110: data <= 19'h7ffdd; 
        10'b0011000111: data <= 19'h7fe4b; 
        10'b0011001000: data <= 19'h7fd5c; 
        10'b0011001001: data <= 19'h7ffc4; 
        10'b0011001010: data <= 19'h7fef0; 
        10'b0011001011: data <= 19'h00005; 
        10'b0011001100: data <= 19'h7fec3; 
        10'b0011001101: data <= 19'h7ffa3; 
        10'b0011001110: data <= 19'h0003d; 
        10'b0011001111: data <= 19'h0026b; 
        10'b0011010000: data <= 19'h00508; 
        10'b0011010001: data <= 19'h004a1; 
        10'b0011010010: data <= 19'h001e6; 
        10'b0011010011: data <= 19'h002f4; 
        10'b0011010100: data <= 19'h00437; 
        10'b0011010101: data <= 19'h007df; 
        10'b0011010110: data <= 19'h005cb; 
        10'b0011010111: data <= 19'h00512; 
        10'b0011011000: data <= 19'h00212; 
        10'b0011011001: data <= 19'h003fa; 
        10'b0011011010: data <= 19'h0045f; 
        10'b0011011011: data <= 19'h0023c; 
        10'b0011011100: data <= 19'h7fe4e; 
        10'b0011011101: data <= 19'h7fd37; 
        10'b0011011110: data <= 19'h7fd80; 
        10'b0011011111: data <= 19'h7ffd9; 
        10'b0011100000: data <= 19'h000c1; 
        10'b0011100001: data <= 19'h00047; 
        10'b0011100010: data <= 19'h7ffae; 
        10'b0011100011: data <= 19'h7fffd; 
        10'b0011100100: data <= 19'h7fe0f; 
        10'b0011100101: data <= 19'h7fe7f; 
        10'b0011100110: data <= 19'h7fec3; 
        10'b0011100111: data <= 19'h7fe7b; 
        10'b0011101000: data <= 19'h7ff32; 
        10'b0011101001: data <= 19'h7ff28; 
        10'b0011101010: data <= 19'h00263; 
        10'b0011101011: data <= 19'h00283; 
        10'b0011101100: data <= 19'h00149; 
        10'b0011101101: data <= 19'h0008a; 
        10'b0011101110: data <= 19'h000e4; 
        10'b0011101111: data <= 19'h0038a; 
        10'b0011110000: data <= 19'h00a53; 
        10'b0011110001: data <= 19'h00838; 
        10'b0011110010: data <= 19'h007a1; 
        10'b0011110011: data <= 19'h00266; 
        10'b0011110100: data <= 19'h00204; 
        10'b0011110101: data <= 19'h001d9; 
        10'b0011110110: data <= 19'h00487; 
        10'b0011110111: data <= 19'h007e3; 
        10'b0011111000: data <= 19'h7ff22; 
        10'b0011111001: data <= 19'h7fd60; 
        10'b0011111010: data <= 19'h7ffbd; 
        10'b0011111011: data <= 19'h7fe9f; 
        10'b0011111100: data <= 19'h7ffc9; 
        10'b0011111101: data <= 19'h7ffde; 
        10'b0011111110: data <= 19'h0003b; 
        10'b0011111111: data <= 19'h0002c; 
        10'b0100000000: data <= 19'h7fd90; 
        10'b0100000001: data <= 19'h7fe44; 
        10'b0100000010: data <= 19'h7fd83; 
        10'b0100000011: data <= 19'h7fe92; 
        10'b0100000100: data <= 19'h7fe97; 
        10'b0100000101: data <= 19'h7ff47; 
        10'b0100000110: data <= 19'h001b7; 
        10'b0100000111: data <= 19'h7fe89; 
        10'b0100001000: data <= 19'h000da; 
        10'b0100001001: data <= 19'h00296; 
        10'b0100001010: data <= 19'h0024c; 
        10'b0100001011: data <= 19'h001f6; 
        10'b0100001100: data <= 19'h005a8; 
        10'b0100001101: data <= 19'h00789; 
        10'b0100001110: data <= 19'h008aa; 
        10'b0100001111: data <= 19'h00503; 
        10'b0100010000: data <= 19'h00187; 
        10'b0100010001: data <= 19'h7ffb8; 
        10'b0100010010: data <= 19'h003b8; 
        10'b0100010011: data <= 19'h00806; 
        10'b0100010100: data <= 19'h00257; 
        10'b0100010101: data <= 19'h7fe06; 
        10'b0100010110: data <= 19'h00007; 
        10'b0100010111: data <= 19'h7ffc2; 
        10'b0100011000: data <= 19'h7febc; 
        10'b0100011001: data <= 19'h0009f; 
        10'b0100011010: data <= 19'h7feef; 
        10'b0100011011: data <= 19'h7fe10; 
        10'b0100011100: data <= 19'h7fe39; 
        10'b0100011101: data <= 19'h7fe98; 
        10'b0100011110: data <= 19'h7fecf; 
        10'b0100011111: data <= 19'h00028; 
        10'b0100100000: data <= 19'h000d2; 
        10'b0100100001: data <= 19'h7ffcf; 
        10'b0100100010: data <= 19'h7fea3; 
        10'b0100100011: data <= 19'h00071; 
        10'b0100100100: data <= 19'h0008e; 
        10'b0100100101: data <= 19'h7ffad; 
        10'b0100100110: data <= 19'h7fd47; 
        10'b0100100111: data <= 19'h7fb52; 
        10'b0100101000: data <= 19'h7fd31; 
        10'b0100101001: data <= 19'h002b7; 
        10'b0100101010: data <= 19'h006e4; 
        10'b0100101011: data <= 19'h00724; 
        10'b0100101100: data <= 19'h00652; 
        10'b0100101101: data <= 19'h00494; 
        10'b0100101110: data <= 19'h006ca; 
        10'b0100101111: data <= 19'h00949; 
        10'b0100110000: data <= 19'h0046b; 
        10'b0100110001: data <= 19'h7fe2d; 
        10'b0100110010: data <= 19'h7fe2c; 
        10'b0100110011: data <= 19'h7fe9a; 
        10'b0100110100: data <= 19'h7ff0e; 
        10'b0100110101: data <= 19'h7febc; 
        10'b0100110110: data <= 19'h00088; 
        10'b0100110111: data <= 19'h7ff9b; 
        10'b0100111000: data <= 19'h7fc84; 
        10'b0100111001: data <= 19'h7ff42; 
        10'b0100111010: data <= 19'h0008b; 
        10'b0100111011: data <= 19'h002a1; 
        10'b0100111100: data <= 19'h001fa; 
        10'b0100111101: data <= 19'h7ff3e; 
        10'b0100111110: data <= 19'h000b1; 
        10'b0100111111: data <= 19'h00012; 
        10'b0101000000: data <= 19'h0015c; 
        10'b0101000001: data <= 19'h7ff13; 
        10'b0101000010: data <= 19'h7f89e; 
        10'b0101000011: data <= 19'h7f252; 
        10'b0101000100: data <= 19'h7f322; 
        10'b0101000101: data <= 19'h7faf9; 
        10'b0101000110: data <= 19'h7ff54; 
        10'b0101000111: data <= 19'h003a2; 
        10'b0101001000: data <= 19'h005d0; 
        10'b0101001001: data <= 19'h00561; 
        10'b0101001010: data <= 19'h00756; 
        10'b0101001011: data <= 19'h00854; 
        10'b0101001100: data <= 19'h005fd; 
        10'b0101001101: data <= 19'h7fed9; 
        10'b0101001110: data <= 19'h7ffec; 
        10'b0101001111: data <= 19'h7fe85; 
        10'b0101010000: data <= 19'h7ff00; 
        10'b0101010001: data <= 19'h7ffaf; 
        10'b0101010010: data <= 19'h7ff8b; 
        10'b0101010011: data <= 19'h7ff9f; 
        10'b0101010100: data <= 19'h7fe09; 
        10'b0101010101: data <= 19'h00051; 
        10'b0101010110: data <= 19'h002dd; 
        10'b0101010111: data <= 19'h002fe; 
        10'b0101011000: data <= 19'h00173; 
        10'b0101011001: data <= 19'h7ff99; 
        10'b0101011010: data <= 19'h0020e; 
        10'b0101011011: data <= 19'h00175; 
        10'b0101011100: data <= 19'h002b0; 
        10'b0101011101: data <= 19'h7fdcb; 
        10'b0101011110: data <= 19'h7f183; 
        10'b0101011111: data <= 19'h7ee0e; 
        10'b0101100000: data <= 19'h7ee22; 
        10'b0101100001: data <= 19'h7f63b; 
        10'b0101100010: data <= 19'h7fe45; 
        10'b0101100011: data <= 19'h7ff48; 
        10'b0101100100: data <= 19'h000e1; 
        10'b0101100101: data <= 19'h00280; 
        10'b0101100110: data <= 19'h00984; 
        10'b0101100111: data <= 19'h008b4; 
        10'b0101101000: data <= 19'h0060c; 
        10'b0101101001: data <= 19'h00037; 
        10'b0101101010: data <= 19'h7ff0c; 
        10'b0101101011: data <= 19'h7ff09; 
        10'b0101101100: data <= 19'h7fe95; 
        10'b0101101101: data <= 19'h7fff8; 
        10'b0101101110: data <= 19'h00080; 
        10'b0101101111: data <= 19'h7fea4; 
        10'b0101110000: data <= 19'h7ff7b; 
        10'b0101110001: data <= 19'h001c7; 
        10'b0101110010: data <= 19'h00378; 
        10'b0101110011: data <= 19'h0047b; 
        10'b0101110100: data <= 19'h00364; 
        10'b0101110101: data <= 19'h00260; 
        10'b0101110110: data <= 19'h0033e; 
        10'b0101110111: data <= 19'h00285; 
        10'b0101111000: data <= 19'h001d1; 
        10'b0101111001: data <= 19'h7f72e; 
        10'b0101111010: data <= 19'h7f17d; 
        10'b0101111011: data <= 19'h7ed8f; 
        10'b0101111100: data <= 19'h7f0db; 
        10'b0101111101: data <= 19'h7f87b; 
        10'b0101111110: data <= 19'h7fc53; 
        10'b0101111111: data <= 19'h7fb11; 
        10'b0110000000: data <= 19'h7fc3b; 
        10'b0110000001: data <= 19'h001a8; 
        10'b0110000010: data <= 19'h0063e; 
        10'b0110000011: data <= 19'h009cd; 
        10'b0110000100: data <= 19'h00591; 
        10'b0110000101: data <= 19'h000e5; 
        10'b0110000110: data <= 19'h00002; 
        10'b0110000111: data <= 19'h0008a; 
        10'b0110001000: data <= 19'h7ffcc; 
        10'b0110001001: data <= 19'h0006d; 
        10'b0110001010: data <= 19'h7fee9; 
        10'b0110001011: data <= 19'h7ff36; 
        10'b0110001100: data <= 19'h7fe4f; 
        10'b0110001101: data <= 19'h00496; 
        10'b0110001110: data <= 19'h005f4; 
        10'b0110001111: data <= 19'h0073b; 
        10'b0110010000: data <= 19'h00378; 
        10'b0110010001: data <= 19'h0042b; 
        10'b0110010010: data <= 19'h00622; 
        10'b0110010011: data <= 19'h00386; 
        10'b0110010100: data <= 19'h000dc; 
        10'b0110010101: data <= 19'h7f852; 
        10'b0110010110: data <= 19'h7eee3; 
        10'b0110010111: data <= 19'h7ed81; 
        10'b0110011000: data <= 19'h7f149; 
        10'b0110011001: data <= 19'h7f7f3; 
        10'b0110011010: data <= 19'h7fc75; 
        10'b0110011011: data <= 19'h7fbb7; 
        10'b0110011100: data <= 19'h00062; 
        10'b0110011101: data <= 19'h0037d; 
        10'b0110011110: data <= 19'h0042a; 
        10'b0110011111: data <= 19'h009e7; 
        10'b0110100000: data <= 19'h00527; 
        10'b0110100001: data <= 19'h7fef5; 
        10'b0110100010: data <= 19'h7ff7b; 
        10'b0110100011: data <= 19'h7fee3; 
        10'b0110100100: data <= 19'h00094; 
        10'b0110100101: data <= 19'h00052; 
        10'b0110100110: data <= 19'h7ff0f; 
        10'b0110100111: data <= 19'h7ffc8; 
        10'b0110101000: data <= 19'h7ffec; 
        10'b0110101001: data <= 19'h0067a; 
        10'b0110101010: data <= 19'h004b3; 
        10'b0110101011: data <= 19'h00677; 
        10'b0110101100: data <= 19'h00477; 
        10'b0110101101: data <= 19'h005eb; 
        10'b0110101110: data <= 19'h0077c; 
        10'b0110101111: data <= 19'h00210; 
        10'b0110110000: data <= 19'h7fa5d; 
        10'b0110110001: data <= 19'h7f1a4; 
        10'b0110110010: data <= 19'h7ecd2; 
        10'b0110110011: data <= 19'h7edbd; 
        10'b0110110100: data <= 19'h7f3aa; 
        10'b0110110101: data <= 19'h7f9fb; 
        10'b0110110110: data <= 19'h7fdc1; 
        10'b0110110111: data <= 19'h7fdd3; 
        10'b0110111000: data <= 19'h001df; 
        10'b0110111001: data <= 19'h001a5; 
        10'b0110111010: data <= 19'h0064a; 
        10'b0110111011: data <= 19'h00765; 
        10'b0110111100: data <= 19'h003d4; 
        10'b0110111101: data <= 19'h7ff9f; 
        10'b0110111110: data <= 19'h0001c; 
        10'b0110111111: data <= 19'h7fefd; 
        10'b0111000000: data <= 19'h0002b; 
        10'b0111000001: data <= 19'h000b9; 
        10'b0111000010: data <= 19'h7fe89; 
        10'b0111000011: data <= 19'h7ff35; 
        10'b0111000100: data <= 19'h00118; 
        10'b0111000101: data <= 19'h005e0; 
        10'b0111000110: data <= 19'h0074d; 
        10'b0111000111: data <= 19'h005a5; 
        10'b0111001000: data <= 19'h003ec; 
        10'b0111001001: data <= 19'h003f4; 
        10'b0111001010: data <= 19'h006aa; 
        10'b0111001011: data <= 19'h7ff20; 
        10'b0111001100: data <= 19'h7f50e; 
        10'b0111001101: data <= 19'h7ecf7; 
        10'b0111001110: data <= 19'h7ed76; 
        10'b0111001111: data <= 19'h7f14b; 
        10'b0111010000: data <= 19'h7f820; 
        10'b0111010001: data <= 19'h7fc52; 
        10'b0111010010: data <= 19'h7fff4; 
        10'b0111010011: data <= 19'h00135; 
        10'b0111010100: data <= 19'h002c5; 
        10'b0111010101: data <= 19'h0041f; 
        10'b0111010110: data <= 19'h005aa; 
        10'b0111010111: data <= 19'h00568; 
        10'b0111011000: data <= 19'h0020f; 
        10'b0111011001: data <= 19'h0001a; 
        10'b0111011010: data <= 19'h7ff54; 
        10'b0111011011: data <= 19'h7ff18; 
        10'b0111011100: data <= 19'h7ff79; 
        10'b0111011101: data <= 19'h0002e; 
        10'b0111011110: data <= 19'h7fec3; 
        10'b0111011111: data <= 19'h7fd98; 
        10'b0111100000: data <= 19'h00034; 
        10'b0111100001: data <= 19'h0042c; 
        10'b0111100010: data <= 19'h0053c; 
        10'b0111100011: data <= 19'h00517; 
        10'b0111100100: data <= 19'h00196; 
        10'b0111100101: data <= 19'h00416; 
        10'b0111100110: data <= 19'h00675; 
        10'b0111100111: data <= 19'h7ff03; 
        10'b0111101000: data <= 19'h7f2e3; 
        10'b0111101001: data <= 19'h7ed39; 
        10'b0111101010: data <= 19'h7ef78; 
        10'b0111101011: data <= 19'h7f625; 
        10'b0111101100: data <= 19'h7feb5; 
        10'b0111101101: data <= 19'h00283; 
        10'b0111101110: data <= 19'h0039f; 
        10'b0111101111: data <= 19'h00356; 
        10'b0111110000: data <= 19'h00441; 
        10'b0111110001: data <= 19'h0033f; 
        10'b0111110010: data <= 19'h00291; 
        10'b0111110011: data <= 19'h002e9; 
        10'b0111110100: data <= 19'h7ffd8; 
        10'b0111110101: data <= 19'h7ff91; 
        10'b0111110110: data <= 19'h0003a; 
        10'b0111110111: data <= 19'h7fefc; 
        10'b0111111000: data <= 19'h7ff4c; 
        10'b0111111001: data <= 19'h0003a; 
        10'b0111111010: data <= 19'h7ff82; 
        10'b0111111011: data <= 19'h7ff14; 
        10'b0111111100: data <= 19'h7ff7f; 
        10'b0111111101: data <= 19'h002aa; 
        10'b0111111110: data <= 19'h0056d; 
        10'b0111111111: data <= 19'h00322; 
        10'b1000000000: data <= 19'h001ed; 
        10'b1000000001: data <= 19'h00565; 
        10'b1000000010: data <= 19'h00a59; 
        10'b1000000011: data <= 19'h00068; 
        10'b1000000100: data <= 19'h7f7a5; 
        10'b1000000101: data <= 19'h7f286; 
        10'b1000000110: data <= 19'h7f69a; 
        10'b1000000111: data <= 19'h7fd23; 
        10'b1000001000: data <= 19'h00308; 
        10'b1000001001: data <= 19'h0033d; 
        10'b1000001010: data <= 19'h00363; 
        10'b1000001011: data <= 19'h001c4; 
        10'b1000001100: data <= 19'h000e1; 
        10'b1000001101: data <= 19'h00178; 
        10'b1000001110: data <= 19'h002d2; 
        10'b1000001111: data <= 19'h001c2; 
        10'b1000010000: data <= 19'h7ffc9; 
        10'b1000010001: data <= 19'h7ff23; 
        10'b1000010010: data <= 19'h0001b; 
        10'b1000010011: data <= 19'h7ff83; 
        10'b1000010100: data <= 19'h7ff91; 
        10'b1000010101: data <= 19'h7ff65; 
        10'b1000010110: data <= 19'h7ff75; 
        10'b1000010111: data <= 19'h7fda7; 
        10'b1000011000: data <= 19'h00101; 
        10'b1000011001: data <= 19'h002eb; 
        10'b1000011010: data <= 19'h006f9; 
        10'b1000011011: data <= 19'h00656; 
        10'b1000011100: data <= 19'h004f4; 
        10'b1000011101: data <= 19'h00693; 
        10'b1000011110: data <= 19'h00a5f; 
        10'b1000011111: data <= 19'h0074b; 
        10'b1000100000: data <= 19'h0018b; 
        10'b1000100001: data <= 19'h7fca5; 
        10'b1000100010: data <= 19'h7fe89; 
        10'b1000100011: data <= 19'h7ff10; 
        10'b1000100100: data <= 19'h00196; 
        10'b1000100101: data <= 19'h7ff45; 
        10'b1000100110: data <= 19'h7fea7; 
        10'b1000100111: data <= 19'h7ff2e; 
        10'b1000101000: data <= 19'h001a2; 
        10'b1000101001: data <= 19'h0017c; 
        10'b1000101010: data <= 19'h002ea; 
        10'b1000101011: data <= 19'h7ff9d; 
        10'b1000101100: data <= 19'h0006b; 
        10'b1000101101: data <= 19'h7ff5d; 
        10'b1000101110: data <= 19'h7fe7f; 
        10'b1000101111: data <= 19'h00085; 
        10'b1000110000: data <= 19'h00083; 
        10'b1000110001: data <= 19'h000ae; 
        10'b1000110010: data <= 19'h7ff84; 
        10'b1000110011: data <= 19'h7fee3; 
        10'b1000110100: data <= 19'h7ff56; 
        10'b1000110101: data <= 19'h002fe; 
        10'b1000110110: data <= 19'h0059b; 
        10'b1000110111: data <= 19'h00421; 
        10'b1000111000: data <= 19'h0051d; 
        10'b1000111001: data <= 19'h00649; 
        10'b1000111010: data <= 19'h009cc; 
        10'b1000111011: data <= 19'h009c8; 
        10'b1000111100: data <= 19'h004e6; 
        10'b1000111101: data <= 19'h0017f; 
        10'b1000111110: data <= 19'h7fefc; 
        10'b1000111111: data <= 19'h000b4; 
        10'b1001000000: data <= 19'h000aa; 
        10'b1001000001: data <= 19'h7fe92; 
        10'b1001000010: data <= 19'h7feea; 
        10'b1001000011: data <= 19'h7fe7a; 
        10'b1001000100: data <= 19'h000cf; 
        10'b1001000101: data <= 19'h00100; 
        10'b1001000110: data <= 19'h0018b; 
        10'b1001000111: data <= 19'h00089; 
        10'b1001001000: data <= 19'h7ff24; 
        10'b1001001001: data <= 19'h7ffce; 
        10'b1001001010: data <= 19'h7feca; 
        10'b1001001011: data <= 19'h7ff5f; 
        10'b1001001100: data <= 19'h7ff1a; 
        10'b1001001101: data <= 19'h7feab; 
        10'b1001001110: data <= 19'h7ff87; 
        10'b1001001111: data <= 19'h7ff1f; 
        10'b1001010000: data <= 19'h7ff71; 
        10'b1001010001: data <= 19'h000c7; 
        10'b1001010010: data <= 19'h00376; 
        10'b1001010011: data <= 19'h005a2; 
        10'b1001010100: data <= 19'h003f3; 
        10'b1001010101: data <= 19'h00449; 
        10'b1001010110: data <= 19'h00863; 
        10'b1001010111: data <= 19'h0097b; 
        10'b1001011000: data <= 19'h0064a; 
        10'b1001011001: data <= 19'h00261; 
        10'b1001011010: data <= 19'h000e3; 
        10'b1001011011: data <= 19'h0002f; 
        10'b1001011100: data <= 19'h7ffd8; 
        10'b1001011101: data <= 19'h7fd68; 
        10'b1001011110: data <= 19'h7fe05; 
        10'b1001011111: data <= 19'h7fedc; 
        10'b1001100000: data <= 19'h000fd; 
        10'b1001100001: data <= 19'h7ffed; 
        10'b1001100010: data <= 19'h7fed3; 
        10'b1001100011: data <= 19'h7fe1e; 
        10'b1001100100: data <= 19'h7ff8a; 
        10'b1001100101: data <= 19'h7ff62; 
        10'b1001100110: data <= 19'h7ff16; 
        10'b1001100111: data <= 19'h7ff38; 
        10'b1001101000: data <= 19'h7fee2; 
        10'b1001101001: data <= 19'h00011; 
        10'b1001101010: data <= 19'h0001b; 
        10'b1001101011: data <= 19'h7ff57; 
        10'b1001101100: data <= 19'h7fed1; 
        10'b1001101101: data <= 19'h0006f; 
        10'b1001101110: data <= 19'h00284; 
        10'b1001101111: data <= 19'h00230; 
        10'b1001110000: data <= 19'h00652; 
        10'b1001110001: data <= 19'h00523; 
        10'b1001110010: data <= 19'h005aa; 
        10'b1001110011: data <= 19'h006bc; 
        10'b1001110100: data <= 19'h005bf; 
        10'b1001110101: data <= 19'h00762; 
        10'b1001110110: data <= 19'h00333; 
        10'b1001110111: data <= 19'h00346; 
        10'b1001111000: data <= 19'h001ca; 
        10'b1001111001: data <= 19'h7fe7b; 
        10'b1001111010: data <= 19'h7feca; 
        10'b1001111011: data <= 19'h7ffea; 
        10'b1001111100: data <= 19'h7fe4a; 
        10'b1001111101: data <= 19'h7fe35; 
        10'b1001111110: data <= 19'h7ff24; 
        10'b1001111111: data <= 19'h7ff11; 
        10'b1010000000: data <= 19'h7ffab; 
        10'b1010000001: data <= 19'h7ff6d; 
        10'b1010000010: data <= 19'h7ff41; 
        10'b1010000011: data <= 19'h7ff9c; 
        10'b1010000100: data <= 19'h7fee0; 
        10'b1010000101: data <= 19'h7ffb2; 
        10'b1010000110: data <= 19'h7fff8; 
        10'b1010000111: data <= 19'h7fea5; 
        10'b1010001000: data <= 19'h7fe9c; 
        10'b1010001001: data <= 19'h7ff99; 
        10'b1010001010: data <= 19'h7ffd6; 
        10'b1010001011: data <= 19'h001c0; 
        10'b1010001100: data <= 19'h00279; 
        10'b1010001101: data <= 19'h005dc; 
        10'b1010001110: data <= 19'h00702; 
        10'b1010001111: data <= 19'h00893; 
        10'b1010010000: data <= 19'h0087c; 
        10'b1010010001: data <= 19'h00516; 
        10'b1010010010: data <= 19'h00425; 
        10'b1010010011: data <= 19'h0024a; 
        10'b1010010100: data <= 19'h000f8; 
        10'b1010010101: data <= 19'h7ffe8; 
        10'b1010010110: data <= 19'h7fcc6; 
        10'b1010010111: data <= 19'h7fbf3; 
        10'b1010011000: data <= 19'h7fcdd; 
        10'b1010011001: data <= 19'h7fe73; 
        10'b1010011010: data <= 19'h7febe; 
        10'b1010011011: data <= 19'h7ffd6; 
        10'b1010011100: data <= 19'h7ff85; 
        10'b1010011101: data <= 19'h00064; 
        10'b1010011110: data <= 19'h7ff54; 
        10'b1010011111: data <= 19'h7fe97; 
        10'b1010100000: data <= 19'h7ff5f; 
        10'b1010100001: data <= 19'h7ffb9; 
        10'b1010100010: data <= 19'h7fe9c; 
        10'b1010100011: data <= 19'h7fff2; 
        10'b1010100100: data <= 19'h7ff9f; 
        10'b1010100101: data <= 19'h7ffa3; 
        10'b1010100110: data <= 19'h7fe55; 
        10'b1010100111: data <= 19'h7fdc6; 
        10'b1010101000: data <= 19'h7fec3; 
        10'b1010101001: data <= 19'h7fee3; 
        10'b1010101010: data <= 19'h0014c; 
        10'b1010101011: data <= 19'h000fa; 
        10'b1010101100: data <= 19'h0025f; 
        10'b1010101101: data <= 19'h00378; 
        10'b1010101110: data <= 19'h001d5; 
        10'b1010101111: data <= 19'h7fe9b; 
        10'b1010110000: data <= 19'h7fdd6; 
        10'b1010110001: data <= 19'h7fd6b; 
        10'b1010110010: data <= 19'h7fdcd; 
        10'b1010110011: data <= 19'h7fcea; 
        10'b1010110100: data <= 19'h7fd0e; 
        10'b1010110101: data <= 19'h7fd38; 
        10'b1010110110: data <= 19'h7ff74; 
        10'b1010110111: data <= 19'h7ff46; 
        10'b1010111000: data <= 19'h7fed5; 
        10'b1010111001: data <= 19'h7ff24; 
        10'b1010111010: data <= 19'h00012; 
        10'b1010111011: data <= 19'h7fefc; 
        10'b1010111100: data <= 19'h7ff26; 
        10'b1010111101: data <= 19'h000cb; 
        10'b1010111110: data <= 19'h7ff94; 
        10'b1010111111: data <= 19'h000a9; 
        10'b1011000000: data <= 19'h000c1; 
        10'b1011000001: data <= 19'h7fff7; 
        10'b1011000010: data <= 19'h7fe7f; 
        10'b1011000011: data <= 19'h7ff58; 
        10'b1011000100: data <= 19'h7fd12; 
        10'b1011000101: data <= 19'h7fd3a; 
        10'b1011000110: data <= 19'h7fc8e; 
        10'b1011000111: data <= 19'h7fb86; 
        10'b1011001000: data <= 19'h7fae3; 
        10'b1011001001: data <= 19'h7fb58; 
        10'b1011001010: data <= 19'h7fa93; 
        10'b1011001011: data <= 19'h7fb1c; 
        10'b1011001100: data <= 19'h7fb60; 
        10'b1011001101: data <= 19'h7fd38; 
        10'b1011001110: data <= 19'h7fdb2; 
        10'b1011001111: data <= 19'h7fe0d; 
        10'b1011010000: data <= 19'h7fdd7; 
        10'b1011010001: data <= 19'h7fe02; 
        10'b1011010010: data <= 19'h7ff55; 
        10'b1011010011: data <= 19'h000c0; 
        10'b1011010100: data <= 19'h0005e; 
        10'b1011010101: data <= 19'h7ff77; 
        10'b1011010110: data <= 19'h7ff49; 
        10'b1011010111: data <= 19'h7ffba; 
        10'b1011011000: data <= 19'h000a1; 
        10'b1011011001: data <= 19'h00091; 
        10'b1011011010: data <= 19'h7ff6d; 
        10'b1011011011: data <= 19'h00009; 
        10'b1011011100: data <= 19'h7ff37; 
        10'b1011011101: data <= 19'h7ff5e; 
        10'b1011011110: data <= 19'h7fea5; 
        10'b1011011111: data <= 19'h00045; 
        10'b1011100000: data <= 19'h7ff48; 
        10'b1011100001: data <= 19'h7fd8c; 
        10'b1011100010: data <= 19'h7fd8a; 
        10'b1011100011: data <= 19'h7fdc6; 
        10'b1011100100: data <= 19'h7ff1a; 
        10'b1011100101: data <= 19'h7fdc7; 
        10'b1011100110: data <= 19'h7fde4; 
        10'b1011100111: data <= 19'h7ff37; 
        10'b1011101000: data <= 19'h7fdc0; 
        10'b1011101001: data <= 19'h7fe2c; 
        10'b1011101010: data <= 19'h7fea3; 
        10'b1011101011: data <= 19'h7fe49; 
        10'b1011101100: data <= 19'h7ff25; 
        10'b1011101101: data <= 19'h7fdf1; 
        10'b1011101110: data <= 19'h7fe43; 
        10'b1011101111: data <= 19'h000ad; 
        10'b1011110000: data <= 19'h7fef0; 
        10'b1011110001: data <= 19'h00033; 
        10'b1011110010: data <= 19'h0008f; 
        10'b1011110011: data <= 19'h7ffdf; 
        10'b1011110100: data <= 19'h7fed7; 
        10'b1011110101: data <= 19'h00077; 
        10'b1011110110: data <= 19'h7ffcd; 
        10'b1011110111: data <= 19'h7ff60; 
        10'b1011111000: data <= 19'h00098; 
        10'b1011111001: data <= 19'h0001e; 
        10'b1011111010: data <= 19'h00035; 
        10'b1011111011: data <= 19'h7fe94; 
        10'b1011111100: data <= 19'h000b2; 
        10'b1011111101: data <= 19'h000ae; 
        10'b1011111110: data <= 19'h0003c; 
        10'b1011111111: data <= 19'h0007d; 
        10'b1100000000: data <= 19'h7ffaa; 
        10'b1100000001: data <= 19'h7ff29; 
        10'b1100000010: data <= 19'h00077; 
        10'b1100000011: data <= 19'h7fec7; 
        10'b1100000100: data <= 19'h7ff8d; 
        10'b1100000101: data <= 19'h7ff24; 
        10'b1100000110: data <= 19'h7ffcb; 
        10'b1100000111: data <= 19'h7ff3e; 
        10'b1100001000: data <= 19'h7fe8d; 
        10'b1100001001: data <= 19'h7feb3; 
        10'b1100001010: data <= 19'h7fe26; 
        10'b1100001011: data <= 19'h7ff92; 
        10'b1100001100: data <= 19'h0004d; 
        10'b1100001101: data <= 19'h7fed3; 
        10'b1100001110: data <= 19'h7fe86; 
        10'b1100001111: data <= 19'h00064; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 14) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 20'hffdee; 
        10'b0000000001: data <= 20'h0012f; 
        10'b0000000010: data <= 20'hfff5b; 
        10'b0000000011: data <= 20'hfffb3; 
        10'b0000000100: data <= 20'h00164; 
        10'b0000000101: data <= 20'hfffdb; 
        10'b0000000110: data <= 20'hffeb0; 
        10'b0000000111: data <= 20'hffe99; 
        10'b0000001000: data <= 20'hfffae; 
        10'b0000001001: data <= 20'hfff4f; 
        10'b0000001010: data <= 20'h0018d; 
        10'b0000001011: data <= 20'hfffe1; 
        10'b0000001100: data <= 20'h000b6; 
        10'b0000001101: data <= 20'hffdfc; 
        10'b0000001110: data <= 20'hfffe3; 
        10'b0000001111: data <= 20'hffd3a; 
        10'b0000010000: data <= 20'hffdb2; 
        10'b0000010001: data <= 20'hfff62; 
        10'b0000010010: data <= 20'hffda0; 
        10'b0000010011: data <= 20'h0018b; 
        10'b0000010100: data <= 20'hffdae; 
        10'b0000010101: data <= 20'hfff42; 
        10'b0000010110: data <= 20'hffd81; 
        10'b0000010111: data <= 20'hfffc0; 
        10'b0000011000: data <= 20'h000c5; 
        10'b0000011001: data <= 20'hfff73; 
        10'b0000011010: data <= 20'hfffe2; 
        10'b0000011011: data <= 20'hfffec; 
        10'b0000011100: data <= 20'h000e1; 
        10'b0000011101: data <= 20'h00115; 
        10'b0000011110: data <= 20'h0005b; 
        10'b0000011111: data <= 20'hffd91; 
        10'b0000100000: data <= 20'hffd72; 
        10'b0000100001: data <= 20'h00022; 
        10'b0000100010: data <= 20'hffdfb; 
        10'b0000100011: data <= 20'hfff70; 
        10'b0000100100: data <= 20'hffe6f; 
        10'b0000100101: data <= 20'hffd25; 
        10'b0000100110: data <= 20'hffe2d; 
        10'b0000100111: data <= 20'h00026; 
        10'b0000101000: data <= 20'h001bd; 
        10'b0000101001: data <= 20'hffd9e; 
        10'b0000101010: data <= 20'hffeb6; 
        10'b0000101011: data <= 20'h000c1; 
        10'b0000101100: data <= 20'hffe06; 
        10'b0000101101: data <= 20'hffd4f; 
        10'b0000101110: data <= 20'h00081; 
        10'b0000101111: data <= 20'h00134; 
        10'b0000110000: data <= 20'hffded; 
        10'b0000110001: data <= 20'h00090; 
        10'b0000110010: data <= 20'hffe3f; 
        10'b0000110011: data <= 20'hffdc6; 
        10'b0000110100: data <= 20'hfff8f; 
        10'b0000110101: data <= 20'h00026; 
        10'b0000110110: data <= 20'hfff4c; 
        10'b0000110111: data <= 20'h00180; 
        10'b0000111000: data <= 20'hffd69; 
        10'b0000111001: data <= 20'hffe68; 
        10'b0000111010: data <= 20'hffe42; 
        10'b0000111011: data <= 20'h000bc; 
        10'b0000111100: data <= 20'h00033; 
        10'b0000111101: data <= 20'hffd53; 
        10'b0000111110: data <= 20'hfff5c; 
        10'b0000111111: data <= 20'h0016e; 
        10'b0001000000: data <= 20'hfff23; 
        10'b0001000001: data <= 20'hffe15; 
        10'b0001000010: data <= 20'hffe27; 
        10'b0001000011: data <= 20'hffcd7; 
        10'b0001000100: data <= 20'hffca3; 
        10'b0001000101: data <= 20'hffed7; 
        10'b0001000110: data <= 20'hffc84; 
        10'b0001000111: data <= 20'hffb87; 
        10'b0001001000: data <= 20'hffcbd; 
        10'b0001001001: data <= 20'hfff25; 
        10'b0001001010: data <= 20'hffd3a; 
        10'b0001001011: data <= 20'hffc6e; 
        10'b0001001100: data <= 20'hfff63; 
        10'b0001001101: data <= 20'h00114; 
        10'b0001001110: data <= 20'h00032; 
        10'b0001001111: data <= 20'hffe07; 
        10'b0001010000: data <= 20'h00159; 
        10'b0001010001: data <= 20'hffd28; 
        10'b0001010010: data <= 20'hfff4f; 
        10'b0001010011: data <= 20'h000a6; 
        10'b0001010100: data <= 20'hffd57; 
        10'b0001010101: data <= 20'hfff60; 
        10'b0001010110: data <= 20'h00181; 
        10'b0001010111: data <= 20'hffd6a; 
        10'b0001011000: data <= 20'hffe25; 
        10'b0001011001: data <= 20'h00138; 
        10'b0001011010: data <= 20'h0007d; 
        10'b0001011011: data <= 20'h0000e; 
        10'b0001011100: data <= 20'h00032; 
        10'b0001011101: data <= 20'hfff51; 
        10'b0001011110: data <= 20'hfff1a; 
        10'b0001011111: data <= 20'hffc7a; 
        10'b0001100000: data <= 20'hffb2c; 
        10'b0001100001: data <= 20'hffd44; 
        10'b0001100010: data <= 20'hffc39; 
        10'b0001100011: data <= 20'hffbba; 
        10'b0001100100: data <= 20'h000b6; 
        10'b0001100101: data <= 20'h00058; 
        10'b0001100110: data <= 20'hffb3d; 
        10'b0001100111: data <= 20'hffbec; 
        10'b0001101000: data <= 20'hffa2a; 
        10'b0001101001: data <= 20'hffbdb; 
        10'b0001101010: data <= 20'hffb00; 
        10'b0001101011: data <= 20'hffc87; 
        10'b0001101100: data <= 20'hffd97; 
        10'b0001101101: data <= 20'h000ea; 
        10'b0001101110: data <= 20'h000e2; 
        10'b0001101111: data <= 20'hffe9f; 
        10'b0001110000: data <= 20'h00059; 
        10'b0001110001: data <= 20'hffd4d; 
        10'b0001110010: data <= 20'hffe1a; 
        10'b0001110011: data <= 20'hffd5c; 
        10'b0001110100: data <= 20'hffd04; 
        10'b0001110101: data <= 20'hfff9c; 
        10'b0001110110: data <= 20'hfff30; 
        10'b0001110111: data <= 20'hffd54; 
        10'b0001111000: data <= 20'hfff19; 
        10'b0001111001: data <= 20'hfff6c; 
        10'b0001111010: data <= 20'hffbac; 
        10'b0001111011: data <= 20'hffbb8; 
        10'b0001111100: data <= 20'hffbca; 
        10'b0001111101: data <= 20'hffbfb; 
        10'b0001111110: data <= 20'hffee7; 
        10'b0001111111: data <= 20'hfff92; 
        10'b0010000000: data <= 20'hffcaf; 
        10'b0010000001: data <= 20'hffce3; 
        10'b0010000010: data <= 20'hffccb; 
        10'b0010000011: data <= 20'hffb85; 
        10'b0010000100: data <= 20'hffe2d; 
        10'b0010000101: data <= 20'hffa3d; 
        10'b0010000110: data <= 20'hffdc2; 
        10'b0010000111: data <= 20'hfffb0; 
        10'b0010001000: data <= 20'hffd7d; 
        10'b0010001001: data <= 20'hffede; 
        10'b0010001010: data <= 20'hffe86; 
        10'b0010001011: data <= 20'hfffc2; 
        10'b0010001100: data <= 20'h000b5; 
        10'b0010001101: data <= 20'hffeba; 
        10'b0010001110: data <= 20'hffff0; 
        10'b0010001111: data <= 20'hffda1; 
        10'b0010010000: data <= 20'hfff5b; 
        10'b0010010001: data <= 20'hffed8; 
        10'b0010010010: data <= 20'hfff28; 
        10'b0010010011: data <= 20'hffe35; 
        10'b0010010100: data <= 20'hfff30; 
        10'b0010010101: data <= 20'hffcc5; 
        10'b0010010110: data <= 20'hffe8b; 
        10'b0010010111: data <= 20'h000f4; 
        10'b0010011000: data <= 20'h003c8; 
        10'b0010011001: data <= 20'h0082a; 
        10'b0010011010: data <= 20'h009de; 
        10'b0010011011: data <= 20'h009c2; 
        10'b0010011100: data <= 20'h00af9; 
        10'b0010011101: data <= 20'h00bcf; 
        10'b0010011110: data <= 20'h00c7f; 
        10'b0010011111: data <= 20'h00467; 
        10'b0010100000: data <= 20'h000c8; 
        10'b0010100001: data <= 20'h00208; 
        10'b0010100010: data <= 20'hffefe; 
        10'b0010100011: data <= 20'hfffdc; 
        10'b0010100100: data <= 20'hffaab; 
        10'b0010100101: data <= 20'hffc20; 
        10'b0010100110: data <= 20'hfffba; 
        10'b0010100111: data <= 20'hffdf0; 
        10'b0010101000: data <= 20'hffeed; 
        10'b0010101001: data <= 20'hfff80; 
        10'b0010101010: data <= 20'h0004a; 
        10'b0010101011: data <= 20'hfff1d; 
        10'b0010101100: data <= 20'h0000b; 
        10'b0010101101: data <= 20'h00022; 
        10'b0010101110: data <= 20'h0004e; 
        10'b0010101111: data <= 20'hfffe1; 
        10'b0010110000: data <= 20'hffd53; 
        10'b0010110001: data <= 20'hffb73; 
        10'b0010110010: data <= 20'h0027d; 
        10'b0010110011: data <= 20'hfff9c; 
        10'b0010110100: data <= 20'h006c4; 
        10'b0010110101: data <= 20'h005fe; 
        10'b0010110110: data <= 20'h005b8; 
        10'b0010110111: data <= 20'h0087d; 
        10'b0010111000: data <= 20'h00a58; 
        10'b0010111001: data <= 20'h00ea9; 
        10'b0010111010: data <= 20'h00da4; 
        10'b0010111011: data <= 20'h00ba1; 
        10'b0010111100: data <= 20'h00b38; 
        10'b0010111101: data <= 20'h00cce; 
        10'b0010111110: data <= 20'h00741; 
        10'b0010111111: data <= 20'h00298; 
        10'b0011000000: data <= 20'hffa71; 
        10'b0011000001: data <= 20'hffa36; 
        10'b0011000010: data <= 20'hffc16; 
        10'b0011000011: data <= 20'h00096; 
        10'b0011000100: data <= 20'h00157; 
        10'b0011000101: data <= 20'h00038; 
        10'b0011000110: data <= 20'hfffb9; 
        10'b0011000111: data <= 20'hffc97; 
        10'b0011001000: data <= 20'hffab7; 
        10'b0011001001: data <= 20'hfff88; 
        10'b0011001010: data <= 20'hffddf; 
        10'b0011001011: data <= 20'h0000a; 
        10'b0011001100: data <= 20'hffd85; 
        10'b0011001101: data <= 20'hfff45; 
        10'b0011001110: data <= 20'h00079; 
        10'b0011001111: data <= 20'h004d5; 
        10'b0011010000: data <= 20'h00a0f; 
        10'b0011010001: data <= 20'h00943; 
        10'b0011010010: data <= 20'h003cc; 
        10'b0011010011: data <= 20'h005e8; 
        10'b0011010100: data <= 20'h0086f; 
        10'b0011010101: data <= 20'h00fbe; 
        10'b0011010110: data <= 20'h00b96; 
        10'b0011010111: data <= 20'h00a23; 
        10'b0011011000: data <= 20'h00425; 
        10'b0011011001: data <= 20'h007f4; 
        10'b0011011010: data <= 20'h008be; 
        10'b0011011011: data <= 20'h00478; 
        10'b0011011100: data <= 20'hffc9c; 
        10'b0011011101: data <= 20'hffa6f; 
        10'b0011011110: data <= 20'hffb00; 
        10'b0011011111: data <= 20'hfffb1; 
        10'b0011100000: data <= 20'h00182; 
        10'b0011100001: data <= 20'h0008d; 
        10'b0011100010: data <= 20'hfff5c; 
        10'b0011100011: data <= 20'hffff9; 
        10'b0011100100: data <= 20'hffc1f; 
        10'b0011100101: data <= 20'hffcfd; 
        10'b0011100110: data <= 20'hffd86; 
        10'b0011100111: data <= 20'hffcf5; 
        10'b0011101000: data <= 20'hffe64; 
        10'b0011101001: data <= 20'hffe50; 
        10'b0011101010: data <= 20'h004c6; 
        10'b0011101011: data <= 20'h00505; 
        10'b0011101100: data <= 20'h00293; 
        10'b0011101101: data <= 20'h00114; 
        10'b0011101110: data <= 20'h001c9; 
        10'b0011101111: data <= 20'h00715; 
        10'b0011110000: data <= 20'h014a6; 
        10'b0011110001: data <= 20'h0106f; 
        10'b0011110010: data <= 20'h00f43; 
        10'b0011110011: data <= 20'h004cc; 
        10'b0011110100: data <= 20'h00409; 
        10'b0011110101: data <= 20'h003b1; 
        10'b0011110110: data <= 20'h0090d; 
        10'b0011110111: data <= 20'h00fc6; 
        10'b0011111000: data <= 20'hffe43; 
        10'b0011111001: data <= 20'hffac0; 
        10'b0011111010: data <= 20'hfff7a; 
        10'b0011111011: data <= 20'hffd3f; 
        10'b0011111100: data <= 20'hfff93; 
        10'b0011111101: data <= 20'hfffbd; 
        10'b0011111110: data <= 20'h00077; 
        10'b0011111111: data <= 20'h00058; 
        10'b0100000000: data <= 20'hffb21; 
        10'b0100000001: data <= 20'hffc87; 
        10'b0100000010: data <= 20'hffb05; 
        10'b0100000011: data <= 20'hffd25; 
        10'b0100000100: data <= 20'hffd2f; 
        10'b0100000101: data <= 20'hffe8e; 
        10'b0100000110: data <= 20'h0036f; 
        10'b0100000111: data <= 20'hffd11; 
        10'b0100001000: data <= 20'h001b4; 
        10'b0100001001: data <= 20'h0052c; 
        10'b0100001010: data <= 20'h00498; 
        10'b0100001011: data <= 20'h003ec; 
        10'b0100001100: data <= 20'h00b50; 
        10'b0100001101: data <= 20'h00f13; 
        10'b0100001110: data <= 20'h01154; 
        10'b0100001111: data <= 20'h00a06; 
        10'b0100010000: data <= 20'h0030d; 
        10'b0100010001: data <= 20'hfff6f; 
        10'b0100010010: data <= 20'h0076f; 
        10'b0100010011: data <= 20'h0100b; 
        10'b0100010100: data <= 20'h004ae; 
        10'b0100010101: data <= 20'hffc0d; 
        10'b0100010110: data <= 20'h0000f; 
        10'b0100010111: data <= 20'hfff84; 
        10'b0100011000: data <= 20'hffd78; 
        10'b0100011001: data <= 20'h0013d; 
        10'b0100011010: data <= 20'hffdde; 
        10'b0100011011: data <= 20'hffc20; 
        10'b0100011100: data <= 20'hffc72; 
        10'b0100011101: data <= 20'hffd2f; 
        10'b0100011110: data <= 20'hffd9e; 
        10'b0100011111: data <= 20'h00050; 
        10'b0100100000: data <= 20'h001a4; 
        10'b0100100001: data <= 20'hfff9f; 
        10'b0100100010: data <= 20'hffd46; 
        10'b0100100011: data <= 20'h000e3; 
        10'b0100100100: data <= 20'h0011d; 
        10'b0100100101: data <= 20'hfff5b; 
        10'b0100100110: data <= 20'hffa8f; 
        10'b0100100111: data <= 20'hff6a4; 
        10'b0100101000: data <= 20'hffa62; 
        10'b0100101001: data <= 20'h0056e; 
        10'b0100101010: data <= 20'h00dc9; 
        10'b0100101011: data <= 20'h00e48; 
        10'b0100101100: data <= 20'h00ca4; 
        10'b0100101101: data <= 20'h00928; 
        10'b0100101110: data <= 20'h00d94; 
        10'b0100101111: data <= 20'h01291; 
        10'b0100110000: data <= 20'h008d7; 
        10'b0100110001: data <= 20'hffc5b; 
        10'b0100110010: data <= 20'hffc57; 
        10'b0100110011: data <= 20'hffd34; 
        10'b0100110100: data <= 20'hffe1b; 
        10'b0100110101: data <= 20'hffd78; 
        10'b0100110110: data <= 20'h00111; 
        10'b0100110111: data <= 20'hfff36; 
        10'b0100111000: data <= 20'hff908; 
        10'b0100111001: data <= 20'hffe84; 
        10'b0100111010: data <= 20'h00117; 
        10'b0100111011: data <= 20'h00542; 
        10'b0100111100: data <= 20'h003f3; 
        10'b0100111101: data <= 20'hffe7d; 
        10'b0100111110: data <= 20'h00162; 
        10'b0100111111: data <= 20'h00024; 
        10'b0101000000: data <= 20'h002b7; 
        10'b0101000001: data <= 20'hffe26; 
        10'b0101000010: data <= 20'hff13c; 
        10'b0101000011: data <= 20'hfe4a5; 
        10'b0101000100: data <= 20'hfe643; 
        10'b0101000101: data <= 20'hff5f2; 
        10'b0101000110: data <= 20'hffea9; 
        10'b0101000111: data <= 20'h00744; 
        10'b0101001000: data <= 20'h00b9f; 
        10'b0101001001: data <= 20'h00ac3; 
        10'b0101001010: data <= 20'h00ead; 
        10'b0101001011: data <= 20'h010a7; 
        10'b0101001100: data <= 20'h00bfa; 
        10'b0101001101: data <= 20'hffdb2; 
        10'b0101001110: data <= 20'hfffd8; 
        10'b0101001111: data <= 20'hffd0a; 
        10'b0101010000: data <= 20'hffe01; 
        10'b0101010001: data <= 20'hfff5d; 
        10'b0101010010: data <= 20'hfff17; 
        10'b0101010011: data <= 20'hfff3e; 
        10'b0101010100: data <= 20'hffc12; 
        10'b0101010101: data <= 20'h000a2; 
        10'b0101010110: data <= 20'h005bb; 
        10'b0101010111: data <= 20'h005fc; 
        10'b0101011000: data <= 20'h002e5; 
        10'b0101011001: data <= 20'hfff32; 
        10'b0101011010: data <= 20'h0041c; 
        10'b0101011011: data <= 20'h002ea; 
        10'b0101011100: data <= 20'h0055f; 
        10'b0101011101: data <= 20'hffb96; 
        10'b0101011110: data <= 20'hfe306; 
        10'b0101011111: data <= 20'hfdc1b; 
        10'b0101100000: data <= 20'hfdc44; 
        10'b0101100001: data <= 20'hfec77; 
        10'b0101100010: data <= 20'hffc8b; 
        10'b0101100011: data <= 20'hffe91; 
        10'b0101100100: data <= 20'h001c2; 
        10'b0101100101: data <= 20'h00501; 
        10'b0101100110: data <= 20'h01309; 
        10'b0101100111: data <= 20'h01168; 
        10'b0101101000: data <= 20'h00c18; 
        10'b0101101001: data <= 20'h0006e; 
        10'b0101101010: data <= 20'hffe19; 
        10'b0101101011: data <= 20'hffe13; 
        10'b0101101100: data <= 20'hffd2a; 
        10'b0101101101: data <= 20'hfffef; 
        10'b0101101110: data <= 20'h000ff; 
        10'b0101101111: data <= 20'hffd49; 
        10'b0101110000: data <= 20'hffef6; 
        10'b0101110001: data <= 20'h0038e; 
        10'b0101110010: data <= 20'h006f1; 
        10'b0101110011: data <= 20'h008f6; 
        10'b0101110100: data <= 20'h006c7; 
        10'b0101110101: data <= 20'h004c0; 
        10'b0101110110: data <= 20'h0067b; 
        10'b0101110111: data <= 20'h00509; 
        10'b0101111000: data <= 20'h003a2; 
        10'b0101111001: data <= 20'hfee5b; 
        10'b0101111010: data <= 20'hfe2f9; 
        10'b0101111011: data <= 20'hfdb1d; 
        10'b0101111100: data <= 20'hfe1b6; 
        10'b0101111101: data <= 20'hff0f7; 
        10'b0101111110: data <= 20'hff8a6; 
        10'b0101111111: data <= 20'hff623; 
        10'b0110000000: data <= 20'hff875; 
        10'b0110000001: data <= 20'h00350; 
        10'b0110000010: data <= 20'h00c7c; 
        10'b0110000011: data <= 20'h0139b; 
        10'b0110000100: data <= 20'h00b21; 
        10'b0110000101: data <= 20'h001cb; 
        10'b0110000110: data <= 20'h00003; 
        10'b0110000111: data <= 20'h00114; 
        10'b0110001000: data <= 20'hfff98; 
        10'b0110001001: data <= 20'h000db; 
        10'b0110001010: data <= 20'hffdd2; 
        10'b0110001011: data <= 20'hffe6c; 
        10'b0110001100: data <= 20'hffc9e; 
        10'b0110001101: data <= 20'h0092b; 
        10'b0110001110: data <= 20'h00be9; 
        10'b0110001111: data <= 20'h00e76; 
        10'b0110010000: data <= 20'h006f0; 
        10'b0110010001: data <= 20'h00857; 
        10'b0110010010: data <= 20'h00c44; 
        10'b0110010011: data <= 20'h0070b; 
        10'b0110010100: data <= 20'h001b9; 
        10'b0110010101: data <= 20'hff0a5; 
        10'b0110010110: data <= 20'hfddc6; 
        10'b0110010111: data <= 20'hfdb03; 
        10'b0110011000: data <= 20'hfe292; 
        10'b0110011001: data <= 20'hfefe6; 
        10'b0110011010: data <= 20'hff8ea; 
        10'b0110011011: data <= 20'hff76f; 
        10'b0110011100: data <= 20'h000c4; 
        10'b0110011101: data <= 20'h006fa; 
        10'b0110011110: data <= 20'h00854; 
        10'b0110011111: data <= 20'h013cf; 
        10'b0110100000: data <= 20'h00a4f; 
        10'b0110100001: data <= 20'hffdea; 
        10'b0110100010: data <= 20'hffef7; 
        10'b0110100011: data <= 20'hffdc6; 
        10'b0110100100: data <= 20'h00127; 
        10'b0110100101: data <= 20'h000a4; 
        10'b0110100110: data <= 20'hffe1e; 
        10'b0110100111: data <= 20'hfff91; 
        10'b0110101000: data <= 20'hfffd8; 
        10'b0110101001: data <= 20'h00cf3; 
        10'b0110101010: data <= 20'h00965; 
        10'b0110101011: data <= 20'h00cee; 
        10'b0110101100: data <= 20'h008ed; 
        10'b0110101101: data <= 20'h00bd6; 
        10'b0110101110: data <= 20'h00ef8; 
        10'b0110101111: data <= 20'h00421; 
        10'b0110110000: data <= 20'hff4bb; 
        10'b0110110001: data <= 20'hfe348; 
        10'b0110110010: data <= 20'hfd9a4; 
        10'b0110110011: data <= 20'hfdb7a; 
        10'b0110110100: data <= 20'hfe754; 
        10'b0110110101: data <= 20'hff3f6; 
        10'b0110110110: data <= 20'hffb82; 
        10'b0110110111: data <= 20'hffba7; 
        10'b0110111000: data <= 20'h003be; 
        10'b0110111001: data <= 20'h0034a; 
        10'b0110111010: data <= 20'h00c94; 
        10'b0110111011: data <= 20'h00eca; 
        10'b0110111100: data <= 20'h007a8; 
        10'b0110111101: data <= 20'hfff3e; 
        10'b0110111110: data <= 20'h00038; 
        10'b0110111111: data <= 20'hffdfa; 
        10'b0111000000: data <= 20'h00055; 
        10'b0111000001: data <= 20'h00173; 
        10'b0111000010: data <= 20'hffd12; 
        10'b0111000011: data <= 20'hffe6a; 
        10'b0111000100: data <= 20'h00230; 
        10'b0111000101: data <= 20'h00bbf; 
        10'b0111000110: data <= 20'h00e99; 
        10'b0111000111: data <= 20'h00b4a; 
        10'b0111001000: data <= 20'h007d7; 
        10'b0111001001: data <= 20'h007e7; 
        10'b0111001010: data <= 20'h00d54; 
        10'b0111001011: data <= 20'hffe40; 
        10'b0111001100: data <= 20'hfea1d; 
        10'b0111001101: data <= 20'hfd9ef; 
        10'b0111001110: data <= 20'hfdaec; 
        10'b0111001111: data <= 20'hfe297; 
        10'b0111010000: data <= 20'hff03f; 
        10'b0111010001: data <= 20'hff8a5; 
        10'b0111010010: data <= 20'hfffe7; 
        10'b0111010011: data <= 20'h0026a; 
        10'b0111010100: data <= 20'h0058b; 
        10'b0111010101: data <= 20'h0083d; 
        10'b0111010110: data <= 20'h00b54; 
        10'b0111010111: data <= 20'h00ad1; 
        10'b0111011000: data <= 20'h0041d; 
        10'b0111011001: data <= 20'h00033; 
        10'b0111011010: data <= 20'hffea8; 
        10'b0111011011: data <= 20'hffe30; 
        10'b0111011100: data <= 20'hffef2; 
        10'b0111011101: data <= 20'h0005b; 
        10'b0111011110: data <= 20'hffd86; 
        10'b0111011111: data <= 20'hffb30; 
        10'b0111100000: data <= 20'h00069; 
        10'b0111100001: data <= 20'h00858; 
        10'b0111100010: data <= 20'h00a78; 
        10'b0111100011: data <= 20'h00a2d; 
        10'b0111100100: data <= 20'h0032d; 
        10'b0111100101: data <= 20'h0082c; 
        10'b0111100110: data <= 20'h00cea; 
        10'b0111100111: data <= 20'hffe06; 
        10'b0111101000: data <= 20'hfe5c7; 
        10'b0111101001: data <= 20'hfda72; 
        10'b0111101010: data <= 20'hfdef0; 
        10'b0111101011: data <= 20'hfec4b; 
        10'b0111101100: data <= 20'hffd69; 
        10'b0111101101: data <= 20'h00506; 
        10'b0111101110: data <= 20'h0073e; 
        10'b0111101111: data <= 20'h006ac; 
        10'b0111110000: data <= 20'h00883; 
        10'b0111110001: data <= 20'h0067d; 
        10'b0111110010: data <= 20'h00521; 
        10'b0111110011: data <= 20'h005d3; 
        10'b0111110100: data <= 20'hfffb0; 
        10'b0111110101: data <= 20'hfff23; 
        10'b0111110110: data <= 20'h00074; 
        10'b0111110111: data <= 20'hffdf8; 
        10'b0111111000: data <= 20'hffe99; 
        10'b0111111001: data <= 20'h00074; 
        10'b0111111010: data <= 20'hfff05; 
        10'b0111111011: data <= 20'hffe28; 
        10'b0111111100: data <= 20'hffefe; 
        10'b0111111101: data <= 20'h00553; 
        10'b0111111110: data <= 20'h00ada; 
        10'b0111111111: data <= 20'h00644; 
        10'b1000000000: data <= 20'h003da; 
        10'b1000000001: data <= 20'h00acb; 
        10'b1000000010: data <= 20'h014b3; 
        10'b1000000011: data <= 20'h000d1; 
        10'b1000000100: data <= 20'hfef4a; 
        10'b1000000101: data <= 20'hfe50c; 
        10'b1000000110: data <= 20'hfed35; 
        10'b1000000111: data <= 20'hffa45; 
        10'b1000001000: data <= 20'h00611; 
        10'b1000001001: data <= 20'h0067a; 
        10'b1000001010: data <= 20'h006c6; 
        10'b1000001011: data <= 20'h00387; 
        10'b1000001100: data <= 20'h001c2; 
        10'b1000001101: data <= 20'h002ef; 
        10'b1000001110: data <= 20'h005a5; 
        10'b1000001111: data <= 20'h00385; 
        10'b1000010000: data <= 20'hfff92; 
        10'b1000010001: data <= 20'hffe45; 
        10'b1000010010: data <= 20'h00035; 
        10'b1000010011: data <= 20'hfff06; 
        10'b1000010100: data <= 20'hfff23; 
        10'b1000010101: data <= 20'hffeca; 
        10'b1000010110: data <= 20'hffeeb; 
        10'b1000010111: data <= 20'hffb4f; 
        10'b1000011000: data <= 20'h00203; 
        10'b1000011001: data <= 20'h005d7; 
        10'b1000011010: data <= 20'h00df1; 
        10'b1000011011: data <= 20'h00cab; 
        10'b1000011100: data <= 20'h009e8; 
        10'b1000011101: data <= 20'h00d26; 
        10'b1000011110: data <= 20'h014be; 
        10'b1000011111: data <= 20'h00e97; 
        10'b1000100000: data <= 20'h00315; 
        10'b1000100001: data <= 20'hff94b; 
        10'b1000100010: data <= 20'hffd11; 
        10'b1000100011: data <= 20'hffe20; 
        10'b1000100100: data <= 20'h0032c; 
        10'b1000100101: data <= 20'hffe8a; 
        10'b1000100110: data <= 20'hffd4e; 
        10'b1000100111: data <= 20'hffe5d; 
        10'b1000101000: data <= 20'h00343; 
        10'b1000101001: data <= 20'h002f8; 
        10'b1000101010: data <= 20'h005d3; 
        10'b1000101011: data <= 20'hfff3a; 
        10'b1000101100: data <= 20'h000d5; 
        10'b1000101101: data <= 20'hffeb9; 
        10'b1000101110: data <= 20'hffcff; 
        10'b1000101111: data <= 20'h0010a; 
        10'b1000110000: data <= 20'h00105; 
        10'b1000110001: data <= 20'h0015c; 
        10'b1000110010: data <= 20'hfff07; 
        10'b1000110011: data <= 20'hffdc5; 
        10'b1000110100: data <= 20'hffeac; 
        10'b1000110101: data <= 20'h005fc; 
        10'b1000110110: data <= 20'h00b35; 
        10'b1000110111: data <= 20'h00841; 
        10'b1000111000: data <= 20'h00a3b; 
        10'b1000111001: data <= 20'h00c91; 
        10'b1000111010: data <= 20'h01397; 
        10'b1000111011: data <= 20'h01391; 
        10'b1000111100: data <= 20'h009cd; 
        10'b1000111101: data <= 20'h002fd; 
        10'b1000111110: data <= 20'hffdf8; 
        10'b1000111111: data <= 20'h00168; 
        10'b1001000000: data <= 20'h00155; 
        10'b1001000001: data <= 20'hffd24; 
        10'b1001000010: data <= 20'hffdd5; 
        10'b1001000011: data <= 20'hffcf5; 
        10'b1001000100: data <= 20'h0019f; 
        10'b1001000101: data <= 20'h00201; 
        10'b1001000110: data <= 20'h00315; 
        10'b1001000111: data <= 20'h00112; 
        10'b1001001000: data <= 20'hffe47; 
        10'b1001001001: data <= 20'hfff9c; 
        10'b1001001010: data <= 20'hffd94; 
        10'b1001001011: data <= 20'hffebe; 
        10'b1001001100: data <= 20'hffe33; 
        10'b1001001101: data <= 20'hffd56; 
        10'b1001001110: data <= 20'hfff0d; 
        10'b1001001111: data <= 20'hffe3e; 
        10'b1001010000: data <= 20'hffee1; 
        10'b1001010001: data <= 20'h0018d; 
        10'b1001010010: data <= 20'h006ed; 
        10'b1001010011: data <= 20'h00b44; 
        10'b1001010100: data <= 20'h007e7; 
        10'b1001010101: data <= 20'h00892; 
        10'b1001010110: data <= 20'h010c5; 
        10'b1001010111: data <= 20'h012f6; 
        10'b1001011000: data <= 20'h00c93; 
        10'b1001011001: data <= 20'h004c2; 
        10'b1001011010: data <= 20'h001c5; 
        10'b1001011011: data <= 20'h0005f; 
        10'b1001011100: data <= 20'hfffb0; 
        10'b1001011101: data <= 20'hffad0; 
        10'b1001011110: data <= 20'hffc0a; 
        10'b1001011111: data <= 20'hffdb9; 
        10'b1001100000: data <= 20'h001fa; 
        10'b1001100001: data <= 20'hfffdb; 
        10'b1001100010: data <= 20'hffda7; 
        10'b1001100011: data <= 20'hffc3c; 
        10'b1001100100: data <= 20'hfff13; 
        10'b1001100101: data <= 20'hffec3; 
        10'b1001100110: data <= 20'hffe2c; 
        10'b1001100111: data <= 20'hffe6f; 
        10'b1001101000: data <= 20'hffdc4; 
        10'b1001101001: data <= 20'h00022; 
        10'b1001101010: data <= 20'h00036; 
        10'b1001101011: data <= 20'hffead; 
        10'b1001101100: data <= 20'hffda3; 
        10'b1001101101: data <= 20'h000df; 
        10'b1001101110: data <= 20'h00509; 
        10'b1001101111: data <= 20'h0045f; 
        10'b1001110000: data <= 20'h00ca3; 
        10'b1001110001: data <= 20'h00a46; 
        10'b1001110010: data <= 20'h00b53; 
        10'b1001110011: data <= 20'h00d78; 
        10'b1001110100: data <= 20'h00b7d; 
        10'b1001110101: data <= 20'h00ec4; 
        10'b1001110110: data <= 20'h00665; 
        10'b1001110111: data <= 20'h0068c; 
        10'b1001111000: data <= 20'h00394; 
        10'b1001111001: data <= 20'hffcf6; 
        10'b1001111010: data <= 20'hffd95; 
        10'b1001111011: data <= 20'hfffd4; 
        10'b1001111100: data <= 20'hffc94; 
        10'b1001111101: data <= 20'hffc6a; 
        10'b1001111110: data <= 20'hffe47; 
        10'b1001111111: data <= 20'hffe22; 
        10'b1010000000: data <= 20'hfff56; 
        10'b1010000001: data <= 20'hffed9; 
        10'b1010000010: data <= 20'hffe83; 
        10'b1010000011: data <= 20'hfff38; 
        10'b1010000100: data <= 20'hffdc0; 
        10'b1010000101: data <= 20'hfff64; 
        10'b1010000110: data <= 20'hffff0; 
        10'b1010000111: data <= 20'hffd49; 
        10'b1010001000: data <= 20'hffd38; 
        10'b1010001001: data <= 20'hfff32; 
        10'b1010001010: data <= 20'hfffab; 
        10'b1010001011: data <= 20'h0037f; 
        10'b1010001100: data <= 20'h004f1; 
        10'b1010001101: data <= 20'h00bb8; 
        10'b1010001110: data <= 20'h00e04; 
        10'b1010001111: data <= 20'h01125; 
        10'b1010010000: data <= 20'h010f9; 
        10'b1010010001: data <= 20'h00a2d; 
        10'b1010010010: data <= 20'h0084a; 
        10'b1010010011: data <= 20'h00494; 
        10'b1010010100: data <= 20'h001f0; 
        10'b1010010101: data <= 20'hfffd0; 
        10'b1010010110: data <= 20'hff98c; 
        10'b1010010111: data <= 20'hff7e7; 
        10'b1010011000: data <= 20'hff9b9; 
        10'b1010011001: data <= 20'hffce6; 
        10'b1010011010: data <= 20'hffd7c; 
        10'b1010011011: data <= 20'hfffad; 
        10'b1010011100: data <= 20'hfff0a; 
        10'b1010011101: data <= 20'h000c9; 
        10'b1010011110: data <= 20'hffea7; 
        10'b1010011111: data <= 20'hffd2e; 
        10'b1010100000: data <= 20'hffebf; 
        10'b1010100001: data <= 20'hfff72; 
        10'b1010100010: data <= 20'hffd38; 
        10'b1010100011: data <= 20'hfffe4; 
        10'b1010100100: data <= 20'hfff3e; 
        10'b1010100101: data <= 20'hfff47; 
        10'b1010100110: data <= 20'hffca9; 
        10'b1010100111: data <= 20'hffb8c; 
        10'b1010101000: data <= 20'hffd86; 
        10'b1010101001: data <= 20'hffdc7; 
        10'b1010101010: data <= 20'h00298; 
        10'b1010101011: data <= 20'h001f5; 
        10'b1010101100: data <= 20'h004bd; 
        10'b1010101101: data <= 20'h006ef; 
        10'b1010101110: data <= 20'h003a9; 
        10'b1010101111: data <= 20'hffd37; 
        10'b1010110000: data <= 20'hffbad; 
        10'b1010110001: data <= 20'hffad6; 
        10'b1010110010: data <= 20'hffb99; 
        10'b1010110011: data <= 20'hff9d3; 
        10'b1010110100: data <= 20'hffa1c; 
        10'b1010110101: data <= 20'hffa70; 
        10'b1010110110: data <= 20'hffee9; 
        10'b1010110111: data <= 20'hffe8b; 
        10'b1010111000: data <= 20'hffdaa; 
        10'b1010111001: data <= 20'hffe48; 
        10'b1010111010: data <= 20'h00023; 
        10'b1010111011: data <= 20'hffdf9; 
        10'b1010111100: data <= 20'hffe4c; 
        10'b1010111101: data <= 20'h00197; 
        10'b1010111110: data <= 20'hfff28; 
        10'b1010111111: data <= 20'h00153; 
        10'b1011000000: data <= 20'h00182; 
        10'b1011000001: data <= 20'hfffed; 
        10'b1011000010: data <= 20'hffcfe; 
        10'b1011000011: data <= 20'hffeaf; 
        10'b1011000100: data <= 20'hffa24; 
        10'b1011000101: data <= 20'hffa74; 
        10'b1011000110: data <= 20'hff91c; 
        10'b1011000111: data <= 20'hff70d; 
        10'b1011001000: data <= 20'hff5c5; 
        10'b1011001001: data <= 20'hff6b0; 
        10'b1011001010: data <= 20'hff527; 
        10'b1011001011: data <= 20'hff637; 
        10'b1011001100: data <= 20'hff6c0; 
        10'b1011001101: data <= 20'hffa70; 
        10'b1011001110: data <= 20'hffb63; 
        10'b1011001111: data <= 20'hffc19; 
        10'b1011010000: data <= 20'hffbad; 
        10'b1011010001: data <= 20'hffc04; 
        10'b1011010010: data <= 20'hffeaa; 
        10'b1011010011: data <= 20'h00180; 
        10'b1011010100: data <= 20'h000bc; 
        10'b1011010101: data <= 20'hffeef; 
        10'b1011010110: data <= 20'hffe93; 
        10'b1011010111: data <= 20'hfff75; 
        10'b1011011000: data <= 20'h00142; 
        10'b1011011001: data <= 20'h00122; 
        10'b1011011010: data <= 20'hffeda; 
        10'b1011011011: data <= 20'h00012; 
        10'b1011011100: data <= 20'hffe6e; 
        10'b1011011101: data <= 20'hffebc; 
        10'b1011011110: data <= 20'hffd4a; 
        10'b1011011111: data <= 20'h00089; 
        10'b1011100000: data <= 20'hffe8f; 
        10'b1011100001: data <= 20'hffb17; 
        10'b1011100010: data <= 20'hffb14; 
        10'b1011100011: data <= 20'hffb8c; 
        10'b1011100100: data <= 20'hffe34; 
        10'b1011100101: data <= 20'hffb8e; 
        10'b1011100110: data <= 20'hffbc8; 
        10'b1011100111: data <= 20'hffe6e; 
        10'b1011101000: data <= 20'hffb81; 
        10'b1011101001: data <= 20'hffc58; 
        10'b1011101010: data <= 20'hffd47; 
        10'b1011101011: data <= 20'hffc92; 
        10'b1011101100: data <= 20'hffe4a; 
        10'b1011101101: data <= 20'hffbe2; 
        10'b1011101110: data <= 20'hffc86; 
        10'b1011101111: data <= 20'h0015a; 
        10'b1011110000: data <= 20'hffddf; 
        10'b1011110001: data <= 20'h00065; 
        10'b1011110010: data <= 20'h0011f; 
        10'b1011110011: data <= 20'hfffbf; 
        10'b1011110100: data <= 20'hffdae; 
        10'b1011110101: data <= 20'h000ee; 
        10'b1011110110: data <= 20'hfff9b; 
        10'b1011110111: data <= 20'hffec0; 
        10'b1011111000: data <= 20'h00130; 
        10'b1011111001: data <= 20'h0003c; 
        10'b1011111010: data <= 20'h0006a; 
        10'b1011111011: data <= 20'hffd28; 
        10'b1011111100: data <= 20'h00164; 
        10'b1011111101: data <= 20'h0015c; 
        10'b1011111110: data <= 20'h00079; 
        10'b1011111111: data <= 20'h000fa; 
        10'b1100000000: data <= 20'hfff53; 
        10'b1100000001: data <= 20'hffe51; 
        10'b1100000010: data <= 20'h000ed; 
        10'b1100000011: data <= 20'hffd8f; 
        10'b1100000100: data <= 20'hfff1a; 
        10'b1100000101: data <= 20'hffe48; 
        10'b1100000110: data <= 20'hfff95; 
        10'b1100000111: data <= 20'hffe7c; 
        10'b1100001000: data <= 20'hffd1a; 
        10'b1100001001: data <= 20'hffd66; 
        10'b1100001010: data <= 20'hffc4c; 
        10'b1100001011: data <= 20'hfff24; 
        10'b1100001100: data <= 20'h00099; 
        10'b1100001101: data <= 20'hffda7; 
        10'b1100001110: data <= 20'hffd0b; 
        10'b1100001111: data <= 20'h000c7; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 15) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 21'h1ffbdc; 
        10'b0000000001: data <= 21'h00025e; 
        10'b0000000010: data <= 21'h1ffeb6; 
        10'b0000000011: data <= 21'h1fff66; 
        10'b0000000100: data <= 21'h0002c8; 
        10'b0000000101: data <= 21'h1fffb6; 
        10'b0000000110: data <= 21'h1ffd5f; 
        10'b0000000111: data <= 21'h1ffd32; 
        10'b0000001000: data <= 21'h1fff5b; 
        10'b0000001001: data <= 21'h1ffe9e; 
        10'b0000001010: data <= 21'h00031a; 
        10'b0000001011: data <= 21'h1fffc1; 
        10'b0000001100: data <= 21'h00016c; 
        10'b0000001101: data <= 21'h1ffbf7; 
        10'b0000001110: data <= 21'h1fffc6; 
        10'b0000001111: data <= 21'h1ffa75; 
        10'b0000010000: data <= 21'h1ffb63; 
        10'b0000010001: data <= 21'h1ffec4; 
        10'b0000010010: data <= 21'h1ffb41; 
        10'b0000010011: data <= 21'h000316; 
        10'b0000010100: data <= 21'h1ffb5c; 
        10'b0000010101: data <= 21'h1ffe85; 
        10'b0000010110: data <= 21'h1ffb01; 
        10'b0000010111: data <= 21'h1fff80; 
        10'b0000011000: data <= 21'h00018b; 
        10'b0000011001: data <= 21'h1ffee5; 
        10'b0000011010: data <= 21'h1fffc5; 
        10'b0000011011: data <= 21'h1fffd8; 
        10'b0000011100: data <= 21'h0001c2; 
        10'b0000011101: data <= 21'h000229; 
        10'b0000011110: data <= 21'h0000b6; 
        10'b0000011111: data <= 21'h1ffb22; 
        10'b0000100000: data <= 21'h1ffae4; 
        10'b0000100001: data <= 21'h000044; 
        10'b0000100010: data <= 21'h1ffbf6; 
        10'b0000100011: data <= 21'h1ffedf; 
        10'b0000100100: data <= 21'h1ffcdf; 
        10'b0000100101: data <= 21'h1ffa4a; 
        10'b0000100110: data <= 21'h1ffc5b; 
        10'b0000100111: data <= 21'h00004c; 
        10'b0000101000: data <= 21'h000379; 
        10'b0000101001: data <= 21'h1ffb3d; 
        10'b0000101010: data <= 21'h1ffd6c; 
        10'b0000101011: data <= 21'h000182; 
        10'b0000101100: data <= 21'h1ffc0d; 
        10'b0000101101: data <= 21'h1ffa9e; 
        10'b0000101110: data <= 21'h000102; 
        10'b0000101111: data <= 21'h000269; 
        10'b0000110000: data <= 21'h1ffbda; 
        10'b0000110001: data <= 21'h000121; 
        10'b0000110010: data <= 21'h1ffc7e; 
        10'b0000110011: data <= 21'h1ffb8c; 
        10'b0000110100: data <= 21'h1fff1e; 
        10'b0000110101: data <= 21'h00004b; 
        10'b0000110110: data <= 21'h1ffe97; 
        10'b0000110111: data <= 21'h0002ff; 
        10'b0000111000: data <= 21'h1ffad1; 
        10'b0000111001: data <= 21'h1ffcd1; 
        10'b0000111010: data <= 21'h1ffc85; 
        10'b0000111011: data <= 21'h000178; 
        10'b0000111100: data <= 21'h000067; 
        10'b0000111101: data <= 21'h1ffaa7; 
        10'b0000111110: data <= 21'h1ffeb9; 
        10'b0000111111: data <= 21'h0002dc; 
        10'b0001000000: data <= 21'h1ffe45; 
        10'b0001000001: data <= 21'h1ffc29; 
        10'b0001000010: data <= 21'h1ffc4f; 
        10'b0001000011: data <= 21'h1ff9ae; 
        10'b0001000100: data <= 21'h1ff945; 
        10'b0001000101: data <= 21'h1ffdad; 
        10'b0001000110: data <= 21'h1ff908; 
        10'b0001000111: data <= 21'h1ff70e; 
        10'b0001001000: data <= 21'h1ff979; 
        10'b0001001001: data <= 21'h1ffe4b; 
        10'b0001001010: data <= 21'h1ffa74; 
        10'b0001001011: data <= 21'h1ff8db; 
        10'b0001001100: data <= 21'h1ffec5; 
        10'b0001001101: data <= 21'h000227; 
        10'b0001001110: data <= 21'h000065; 
        10'b0001001111: data <= 21'h1ffc0e; 
        10'b0001010000: data <= 21'h0002b1; 
        10'b0001010001: data <= 21'h1ffa50; 
        10'b0001010010: data <= 21'h1ffe9e; 
        10'b0001010011: data <= 21'h00014c; 
        10'b0001010100: data <= 21'h1ffaae; 
        10'b0001010101: data <= 21'h1ffec0; 
        10'b0001010110: data <= 21'h000301; 
        10'b0001010111: data <= 21'h1ffad3; 
        10'b0001011000: data <= 21'h1ffc49; 
        10'b0001011001: data <= 21'h00026f; 
        10'b0001011010: data <= 21'h0000fb; 
        10'b0001011011: data <= 21'h00001c; 
        10'b0001011100: data <= 21'h000064; 
        10'b0001011101: data <= 21'h1ffea3; 
        10'b0001011110: data <= 21'h1ffe33; 
        10'b0001011111: data <= 21'h1ff8f4; 
        10'b0001100000: data <= 21'h1ff659; 
        10'b0001100001: data <= 21'h1ffa89; 
        10'b0001100010: data <= 21'h1ff872; 
        10'b0001100011: data <= 21'h1ff773; 
        10'b0001100100: data <= 21'h00016c; 
        10'b0001100101: data <= 21'h0000af; 
        10'b0001100110: data <= 21'h1ff679; 
        10'b0001100111: data <= 21'h1ff7d9; 
        10'b0001101000: data <= 21'h1ff455; 
        10'b0001101001: data <= 21'h1ff7b6; 
        10'b0001101010: data <= 21'h1ff600; 
        10'b0001101011: data <= 21'h1ff90e; 
        10'b0001101100: data <= 21'h1ffb2e; 
        10'b0001101101: data <= 21'h0001d4; 
        10'b0001101110: data <= 21'h0001c5; 
        10'b0001101111: data <= 21'h1ffd3e; 
        10'b0001110000: data <= 21'h0000b1; 
        10'b0001110001: data <= 21'h1ffa99; 
        10'b0001110010: data <= 21'h1ffc33; 
        10'b0001110011: data <= 21'h1ffab9; 
        10'b0001110100: data <= 21'h1ffa09; 
        10'b0001110101: data <= 21'h1fff38; 
        10'b0001110110: data <= 21'h1ffe61; 
        10'b0001110111: data <= 21'h1ffaa8; 
        10'b0001111000: data <= 21'h1ffe32; 
        10'b0001111001: data <= 21'h1ffed8; 
        10'b0001111010: data <= 21'h1ff758; 
        10'b0001111011: data <= 21'h1ff771; 
        10'b0001111100: data <= 21'h1ff793; 
        10'b0001111101: data <= 21'h1ff7f6; 
        10'b0001111110: data <= 21'h1ffdcf; 
        10'b0001111111: data <= 21'h1fff24; 
        10'b0010000000: data <= 21'h1ff95e; 
        10'b0010000001: data <= 21'h1ff9c6; 
        10'b0010000010: data <= 21'h1ff995; 
        10'b0010000011: data <= 21'h1ff70a; 
        10'b0010000100: data <= 21'h1ffc5b; 
        10'b0010000101: data <= 21'h1ff47a; 
        10'b0010000110: data <= 21'h1ffb84; 
        10'b0010000111: data <= 21'h1fff60; 
        10'b0010001000: data <= 21'h1ffafb; 
        10'b0010001001: data <= 21'h1ffdbd; 
        10'b0010001010: data <= 21'h1ffd0d; 
        10'b0010001011: data <= 21'h1fff84; 
        10'b0010001100: data <= 21'h00016a; 
        10'b0010001101: data <= 21'h1ffd75; 
        10'b0010001110: data <= 21'h1fffe0; 
        10'b0010001111: data <= 21'h1ffb43; 
        10'b0010010000: data <= 21'h1ffeb7; 
        10'b0010010001: data <= 21'h1ffdb0; 
        10'b0010010010: data <= 21'h1ffe4f; 
        10'b0010010011: data <= 21'h1ffc6a; 
        10'b0010010100: data <= 21'h1ffe60; 
        10'b0010010101: data <= 21'h1ff98a; 
        10'b0010010110: data <= 21'h1ffd16; 
        10'b0010010111: data <= 21'h0001e7; 
        10'b0010011000: data <= 21'h000790; 
        10'b0010011001: data <= 21'h001055; 
        10'b0010011010: data <= 21'h0013bc; 
        10'b0010011011: data <= 21'h001383; 
        10'b0010011100: data <= 21'h0015f2; 
        10'b0010011101: data <= 21'h00179e; 
        10'b0010011110: data <= 21'h0018fd; 
        10'b0010011111: data <= 21'h0008cf; 
        10'b0010100000: data <= 21'h000190; 
        10'b0010100001: data <= 21'h000410; 
        10'b0010100010: data <= 21'h1ffdfc; 
        10'b0010100011: data <= 21'h1fffb7; 
        10'b0010100100: data <= 21'h1ff555; 
        10'b0010100101: data <= 21'h1ff841; 
        10'b0010100110: data <= 21'h1fff74; 
        10'b0010100111: data <= 21'h1ffbe0; 
        10'b0010101000: data <= 21'h1ffddb; 
        10'b0010101001: data <= 21'h1fff00; 
        10'b0010101010: data <= 21'h000094; 
        10'b0010101011: data <= 21'h1ffe3b; 
        10'b0010101100: data <= 21'h000015; 
        10'b0010101101: data <= 21'h000044; 
        10'b0010101110: data <= 21'h00009c; 
        10'b0010101111: data <= 21'h1fffc2; 
        10'b0010110000: data <= 21'h1ffaa6; 
        10'b0010110001: data <= 21'h1ff6e7; 
        10'b0010110010: data <= 21'h0004fa; 
        10'b0010110011: data <= 21'h1fff38; 
        10'b0010110100: data <= 21'h000d89; 
        10'b0010110101: data <= 21'h000bfb; 
        10'b0010110110: data <= 21'h000b70; 
        10'b0010110111: data <= 21'h0010f9; 
        10'b0010111000: data <= 21'h0014b1; 
        10'b0010111001: data <= 21'h001d52; 
        10'b0010111010: data <= 21'h001b47; 
        10'b0010111011: data <= 21'h001742; 
        10'b0010111100: data <= 21'h001670; 
        10'b0010111101: data <= 21'h00199c; 
        10'b0010111110: data <= 21'h000e83; 
        10'b0010111111: data <= 21'h000530; 
        10'b0011000000: data <= 21'h1ff4e2; 
        10'b0011000001: data <= 21'h1ff46d; 
        10'b0011000010: data <= 21'h1ff82b; 
        10'b0011000011: data <= 21'h00012c; 
        10'b0011000100: data <= 21'h0002ae; 
        10'b0011000101: data <= 21'h00006f; 
        10'b0011000110: data <= 21'h1fff73; 
        10'b0011000111: data <= 21'h1ff92d; 
        10'b0011001000: data <= 21'h1ff56e; 
        10'b0011001001: data <= 21'h1fff11; 
        10'b0011001010: data <= 21'h1ffbbe; 
        10'b0011001011: data <= 21'h000014; 
        10'b0011001100: data <= 21'h1ffb0a; 
        10'b0011001101: data <= 21'h1ffe8a; 
        10'b0011001110: data <= 21'h0000f2; 
        10'b0011001111: data <= 21'h0009aa; 
        10'b0011010000: data <= 21'h00141e; 
        10'b0011010001: data <= 21'h001286; 
        10'b0011010010: data <= 21'h000798; 
        10'b0011010011: data <= 21'h000bd0; 
        10'b0011010100: data <= 21'h0010de; 
        10'b0011010101: data <= 21'h001f7c; 
        10'b0011010110: data <= 21'h00172b; 
        10'b0011010111: data <= 21'h001446; 
        10'b0011011000: data <= 21'h000849; 
        10'b0011011001: data <= 21'h000fe8; 
        10'b0011011010: data <= 21'h00117c; 
        10'b0011011011: data <= 21'h0008f1; 
        10'b0011011100: data <= 21'h1ff937; 
        10'b0011011101: data <= 21'h1ff4de; 
        10'b0011011110: data <= 21'h1ff600; 
        10'b0011011111: data <= 21'h1fff63; 
        10'b0011100000: data <= 21'h000305; 
        10'b0011100001: data <= 21'h00011b; 
        10'b0011100010: data <= 21'h1ffeb8; 
        10'b0011100011: data <= 21'h1ffff3; 
        10'b0011100100: data <= 21'h1ff83e; 
        10'b0011100101: data <= 21'h1ff9fb; 
        10'b0011100110: data <= 21'h1ffb0d; 
        10'b0011100111: data <= 21'h1ff9ea; 
        10'b0011101000: data <= 21'h1ffcc9; 
        10'b0011101001: data <= 21'h1ffca0; 
        10'b0011101010: data <= 21'h00098c; 
        10'b0011101011: data <= 21'h000a0a; 
        10'b0011101100: data <= 21'h000525; 
        10'b0011101101: data <= 21'h000228; 
        10'b0011101110: data <= 21'h000391; 
        10'b0011101111: data <= 21'h000e2a; 
        10'b0011110000: data <= 21'h00294c; 
        10'b0011110001: data <= 21'h0020df; 
        10'b0011110010: data <= 21'h001e85; 
        10'b0011110011: data <= 21'h000998; 
        10'b0011110100: data <= 21'h000812; 
        10'b0011110101: data <= 21'h000763; 
        10'b0011110110: data <= 21'h00121a; 
        10'b0011110111: data <= 21'h001f8b; 
        10'b0011111000: data <= 21'h1ffc87; 
        10'b0011111001: data <= 21'h1ff581; 
        10'b0011111010: data <= 21'h1ffef5; 
        10'b0011111011: data <= 21'h1ffa7e; 
        10'b0011111100: data <= 21'h1fff25; 
        10'b0011111101: data <= 21'h1fff7a; 
        10'b0011111110: data <= 21'h0000ed; 
        10'b0011111111: data <= 21'h0000b0; 
        10'b0100000000: data <= 21'h1ff641; 
        10'b0100000001: data <= 21'h1ff90e; 
        10'b0100000010: data <= 21'h1ff60a; 
        10'b0100000011: data <= 21'h1ffa49; 
        10'b0100000100: data <= 21'h1ffa5e; 
        10'b0100000101: data <= 21'h1ffd1d; 
        10'b0100000110: data <= 21'h0006dd; 
        10'b0100000111: data <= 21'h1ffa23; 
        10'b0100001000: data <= 21'h000368; 
        10'b0100001001: data <= 21'h000a57; 
        10'b0100001010: data <= 21'h000931; 
        10'b0100001011: data <= 21'h0007d8; 
        10'b0100001100: data <= 21'h00169f; 
        10'b0100001101: data <= 21'h001e25; 
        10'b0100001110: data <= 21'h0022a8; 
        10'b0100001111: data <= 21'h00140c; 
        10'b0100010000: data <= 21'h00061a; 
        10'b0100010001: data <= 21'h1ffedf; 
        10'b0100010010: data <= 21'h000ede; 
        10'b0100010011: data <= 21'h002016; 
        10'b0100010100: data <= 21'h00095c; 
        10'b0100010101: data <= 21'h1ff81a; 
        10'b0100010110: data <= 21'h00001d; 
        10'b0100010111: data <= 21'h1fff07; 
        10'b0100011000: data <= 21'h1ffaf0; 
        10'b0100011001: data <= 21'h00027a; 
        10'b0100011010: data <= 21'h1ffbbc; 
        10'b0100011011: data <= 21'h1ff83f; 
        10'b0100011100: data <= 21'h1ff8e4; 
        10'b0100011101: data <= 21'h1ffa5f; 
        10'b0100011110: data <= 21'h1ffb3b; 
        10'b0100011111: data <= 21'h0000a0; 
        10'b0100100000: data <= 21'h000347; 
        10'b0100100001: data <= 21'h1fff3d; 
        10'b0100100010: data <= 21'h1ffa8c; 
        10'b0100100011: data <= 21'h0001c5; 
        10'b0100100100: data <= 21'h000239; 
        10'b0100100101: data <= 21'h1ffeb6; 
        10'b0100100110: data <= 21'h1ff51e; 
        10'b0100100111: data <= 21'h1fed48; 
        10'b0100101000: data <= 21'h1ff4c3; 
        10'b0100101001: data <= 21'h000adc; 
        10'b0100101010: data <= 21'h001b91; 
        10'b0100101011: data <= 21'h001c90; 
        10'b0100101100: data <= 21'h001947; 
        10'b0100101101: data <= 21'h001251; 
        10'b0100101110: data <= 21'h001b28; 
        10'b0100101111: data <= 21'h002523; 
        10'b0100110000: data <= 21'h0011ae; 
        10'b0100110001: data <= 21'h1ff8b6; 
        10'b0100110010: data <= 21'h1ff8af; 
        10'b0100110011: data <= 21'h1ffa68; 
        10'b0100110100: data <= 21'h1ffc36; 
        10'b0100110101: data <= 21'h1ffaef; 
        10'b0100110110: data <= 21'h000221; 
        10'b0100110111: data <= 21'h1ffe6d; 
        10'b0100111000: data <= 21'h1ff211; 
        10'b0100111001: data <= 21'h1ffd07; 
        10'b0100111010: data <= 21'h00022d; 
        10'b0100111011: data <= 21'h000a84; 
        10'b0100111100: data <= 21'h0007e6; 
        10'b0100111101: data <= 21'h1ffcf9; 
        10'b0100111110: data <= 21'h0002c4; 
        10'b0100111111: data <= 21'h000048; 
        10'b0101000000: data <= 21'h00056e; 
        10'b0101000001: data <= 21'h1ffc4d; 
        10'b0101000010: data <= 21'h1fe278; 
        10'b0101000011: data <= 21'h1fc949; 
        10'b0101000100: data <= 21'h1fcc86; 
        10'b0101000101: data <= 21'h1febe4; 
        10'b0101000110: data <= 21'h1ffd52; 
        10'b0101000111: data <= 21'h000e87; 
        10'b0101001000: data <= 21'h00173f; 
        10'b0101001001: data <= 21'h001585; 
        10'b0101001010: data <= 21'h001d59; 
        10'b0101001011: data <= 21'h00214e; 
        10'b0101001100: data <= 21'h0017f3; 
        10'b0101001101: data <= 21'h1ffb65; 
        10'b0101001110: data <= 21'h1fffb1; 
        10'b0101001111: data <= 21'h1ffa13; 
        10'b0101010000: data <= 21'h1ffc01; 
        10'b0101010001: data <= 21'h1ffebb; 
        10'b0101010010: data <= 21'h1ffe2d; 
        10'b0101010011: data <= 21'h1ffe7c; 
        10'b0101010100: data <= 21'h1ff825; 
        10'b0101010101: data <= 21'h000143; 
        10'b0101010110: data <= 21'h000b75; 
        10'b0101010111: data <= 21'h000bf8; 
        10'b0101011000: data <= 21'h0005ca; 
        10'b0101011001: data <= 21'h1ffe65; 
        10'b0101011010: data <= 21'h000837; 
        10'b0101011011: data <= 21'h0005d4; 
        10'b0101011100: data <= 21'h000abf; 
        10'b0101011101: data <= 21'h1ff72b; 
        10'b0101011110: data <= 21'h1fc60c; 
        10'b0101011111: data <= 21'h1fb837; 
        10'b0101100000: data <= 21'h1fb887; 
        10'b0101100001: data <= 21'h1fd8ed; 
        10'b0101100010: data <= 21'h1ff915; 
        10'b0101100011: data <= 21'h1ffd22; 
        10'b0101100100: data <= 21'h000383; 
        10'b0101100101: data <= 21'h000a01; 
        10'b0101100110: data <= 21'h002611; 
        10'b0101100111: data <= 21'h0022d0; 
        10'b0101101000: data <= 21'h001830; 
        10'b0101101001: data <= 21'h0000dd; 
        10'b0101101010: data <= 21'h1ffc32; 
        10'b0101101011: data <= 21'h1ffc25; 
        10'b0101101100: data <= 21'h1ffa53; 
        10'b0101101101: data <= 21'h1fffdf; 
        10'b0101101110: data <= 21'h0001ff; 
        10'b0101101111: data <= 21'h1ffa92; 
        10'b0101110000: data <= 21'h1ffdec; 
        10'b0101110001: data <= 21'h00071c; 
        10'b0101110010: data <= 21'h000de2; 
        10'b0101110011: data <= 21'h0011ec; 
        10'b0101110100: data <= 21'h000d8f; 
        10'b0101110101: data <= 21'h00097f; 
        10'b0101110110: data <= 21'h000cf6; 
        10'b0101110111: data <= 21'h000a13; 
        10'b0101111000: data <= 21'h000744; 
        10'b0101111001: data <= 21'h1fdcb6; 
        10'b0101111010: data <= 21'h1fc5f2; 
        10'b0101111011: data <= 21'h1fb63b; 
        10'b0101111100: data <= 21'h1fc36c; 
        10'b0101111101: data <= 21'h1fe1ed; 
        10'b0101111110: data <= 21'h1ff14c; 
        10'b0101111111: data <= 21'h1fec45; 
        10'b0110000000: data <= 21'h1ff0ea; 
        10'b0110000001: data <= 21'h0006a0; 
        10'b0110000010: data <= 21'h0018f8; 
        10'b0110000011: data <= 21'h002736; 
        10'b0110000100: data <= 21'h001643; 
        10'b0110000101: data <= 21'h000396; 
        10'b0110000110: data <= 21'h000006; 
        10'b0110000111: data <= 21'h000229; 
        10'b0110001000: data <= 21'h1fff30; 
        10'b0110001001: data <= 21'h0001b6; 
        10'b0110001010: data <= 21'h1ffba5; 
        10'b0110001011: data <= 21'h1ffcd9; 
        10'b0110001100: data <= 21'h1ff93c; 
        10'b0110001101: data <= 21'h001257; 
        10'b0110001110: data <= 21'h0017d2; 
        10'b0110001111: data <= 21'h001cec; 
        10'b0110010000: data <= 21'h000de1; 
        10'b0110010001: data <= 21'h0010ad; 
        10'b0110010010: data <= 21'h001888; 
        10'b0110010011: data <= 21'h000e16; 
        10'b0110010100: data <= 21'h000371; 
        10'b0110010101: data <= 21'h1fe149; 
        10'b0110010110: data <= 21'h1fbb8c; 
        10'b0110010111: data <= 21'h1fb606; 
        10'b0110011000: data <= 21'h1fc524; 
        10'b0110011001: data <= 21'h1fdfcd; 
        10'b0110011010: data <= 21'h1ff1d4; 
        10'b0110011011: data <= 21'h1feedd; 
        10'b0110011100: data <= 21'h000188; 
        10'b0110011101: data <= 21'h000df3; 
        10'b0110011110: data <= 21'h0010a8; 
        10'b0110011111: data <= 21'h00279e; 
        10'b0110100000: data <= 21'h00149d; 
        10'b0110100001: data <= 21'h1ffbd5; 
        10'b0110100010: data <= 21'h1ffdee; 
        10'b0110100011: data <= 21'h1ffb8d; 
        10'b0110100100: data <= 21'h00024e; 
        10'b0110100101: data <= 21'h000148; 
        10'b0110100110: data <= 21'h1ffc3b; 
        10'b0110100111: data <= 21'h1fff22; 
        10'b0110101000: data <= 21'h1fffb1; 
        10'b0110101001: data <= 21'h0019e7; 
        10'b0110101010: data <= 21'h0012ca; 
        10'b0110101011: data <= 21'h0019dc; 
        10'b0110101100: data <= 21'h0011db; 
        10'b0110101101: data <= 21'h0017ac; 
        10'b0110101110: data <= 21'h001def; 
        10'b0110101111: data <= 21'h000842; 
        10'b0110110000: data <= 21'h1fe976; 
        10'b0110110001: data <= 21'h1fc68f; 
        10'b0110110010: data <= 21'h1fb348; 
        10'b0110110011: data <= 21'h1fb6f4; 
        10'b0110110100: data <= 21'h1fcea8; 
        10'b0110110101: data <= 21'h1fe7eb; 
        10'b0110110110: data <= 21'h1ff703; 
        10'b0110110111: data <= 21'h1ff74d; 
        10'b0110111000: data <= 21'h00077c; 
        10'b0110111001: data <= 21'h000693; 
        10'b0110111010: data <= 21'h001929; 
        10'b0110111011: data <= 21'h001d94; 
        10'b0110111100: data <= 21'h000f50; 
        10'b0110111101: data <= 21'h1ffe7d; 
        10'b0110111110: data <= 21'h000070; 
        10'b0110111111: data <= 21'h1ffbf4; 
        10'b0111000000: data <= 21'h0000ab; 
        10'b0111000001: data <= 21'h0002e6; 
        10'b0111000010: data <= 21'h1ffa24; 
        10'b0111000011: data <= 21'h1ffcd4; 
        10'b0111000100: data <= 21'h00045f; 
        10'b0111000101: data <= 21'h00177f; 
        10'b0111000110: data <= 21'h001d32; 
        10'b0111000111: data <= 21'h001695; 
        10'b0111001000: data <= 21'h000fae; 
        10'b0111001001: data <= 21'h000fcf; 
        10'b0111001010: data <= 21'h001aa8; 
        10'b0111001011: data <= 21'h1ffc80; 
        10'b0111001100: data <= 21'h1fd439; 
        10'b0111001101: data <= 21'h1fb3dd; 
        10'b0111001110: data <= 21'h1fb5d9; 
        10'b0111001111: data <= 21'h1fc52e; 
        10'b0111010000: data <= 21'h1fe07f; 
        10'b0111010001: data <= 21'h1ff149; 
        10'b0111010010: data <= 21'h1fffce; 
        10'b0111010011: data <= 21'h0004d3; 
        10'b0111010100: data <= 21'h000b16; 
        10'b0111010101: data <= 21'h00107a; 
        10'b0111010110: data <= 21'h0016a9; 
        10'b0111010111: data <= 21'h0015a2; 
        10'b0111011000: data <= 21'h00083a; 
        10'b0111011001: data <= 21'h000067; 
        10'b0111011010: data <= 21'h1ffd50; 
        10'b0111011011: data <= 21'h1ffc61; 
        10'b0111011100: data <= 21'h1ffde5; 
        10'b0111011101: data <= 21'h0000b6; 
        10'b0111011110: data <= 21'h1ffb0c; 
        10'b0111011111: data <= 21'h1ff660; 
        10'b0111100000: data <= 21'h0000d1; 
        10'b0111100001: data <= 21'h0010b1; 
        10'b0111100010: data <= 21'h0014f0; 
        10'b0111100011: data <= 21'h00145b; 
        10'b0111100100: data <= 21'h00065a; 
        10'b0111100101: data <= 21'h001058; 
        10'b0111100110: data <= 21'h0019d4; 
        10'b0111100111: data <= 21'h1ffc0c; 
        10'b0111101000: data <= 21'h1fcb8d; 
        10'b0111101001: data <= 21'h1fb4e5; 
        10'b0111101010: data <= 21'h1fbde0; 
        10'b0111101011: data <= 21'h1fd896; 
        10'b0111101100: data <= 21'h1ffad3; 
        10'b0111101101: data <= 21'h000a0c; 
        10'b0111101110: data <= 21'h000e7b; 
        10'b0111101111: data <= 21'h000d58; 
        10'b0111110000: data <= 21'h001106; 
        10'b0111110001: data <= 21'h000cfa; 
        10'b0111110010: data <= 21'h000a42; 
        10'b0111110011: data <= 21'h000ba6; 
        10'b0111110100: data <= 21'h1fff60; 
        10'b0111110101: data <= 21'h1ffe45; 
        10'b0111110110: data <= 21'h0000e8; 
        10'b0111110111: data <= 21'h1ffbf0; 
        10'b0111111000: data <= 21'h1ffd31; 
        10'b0111111001: data <= 21'h0000e8; 
        10'b0111111010: data <= 21'h1ffe09; 
        10'b0111111011: data <= 21'h1ffc50; 
        10'b0111111100: data <= 21'h1ffdfb; 
        10'b0111111101: data <= 21'h000aa6; 
        10'b0111111110: data <= 21'h0015b5; 
        10'b0111111111: data <= 21'h000c88; 
        10'b1000000000: data <= 21'h0007b3; 
        10'b1000000001: data <= 21'h001596; 
        10'b1000000010: data <= 21'h002965; 
        10'b1000000011: data <= 21'h0001a1; 
        10'b1000000100: data <= 21'h1fde95; 
        10'b1000000101: data <= 21'h1fca17; 
        10'b1000000110: data <= 21'h1fda69; 
        10'b1000000111: data <= 21'h1ff48b; 
        10'b1000001000: data <= 21'h000c22; 
        10'b1000001001: data <= 21'h000cf3; 
        10'b1000001010: data <= 21'h000d8c; 
        10'b1000001011: data <= 21'h00070e; 
        10'b1000001100: data <= 21'h000384; 
        10'b1000001101: data <= 21'h0005de; 
        10'b1000001110: data <= 21'h000b49; 
        10'b1000001111: data <= 21'h00070a; 
        10'b1000010000: data <= 21'h1fff23; 
        10'b1000010001: data <= 21'h1ffc8b; 
        10'b1000010010: data <= 21'h00006b; 
        10'b1000010011: data <= 21'h1ffe0c; 
        10'b1000010100: data <= 21'h1ffe45; 
        10'b1000010101: data <= 21'h1ffd95; 
        10'b1000010110: data <= 21'h1ffdd5; 
        10'b1000010111: data <= 21'h1ff69e; 
        10'b1000011000: data <= 21'h000405; 
        10'b1000011001: data <= 21'h000bae; 
        10'b1000011010: data <= 21'h001be3; 
        10'b1000011011: data <= 21'h001957; 
        10'b1000011100: data <= 21'h0013d1; 
        10'b1000011101: data <= 21'h001a4c; 
        10'b1000011110: data <= 21'h00297d; 
        10'b1000011111: data <= 21'h001d2e; 
        10'b1000100000: data <= 21'h00062b; 
        10'b1000100001: data <= 21'h1ff296; 
        10'b1000100010: data <= 21'h1ffa23; 
        10'b1000100011: data <= 21'h1ffc3f; 
        10'b1000100100: data <= 21'h000658; 
        10'b1000100101: data <= 21'h1ffd14; 
        10'b1000100110: data <= 21'h1ffa9d; 
        10'b1000100111: data <= 21'h1ffcba; 
        10'b1000101000: data <= 21'h000686; 
        10'b1000101001: data <= 21'h0005f0; 
        10'b1000101010: data <= 21'h000ba7; 
        10'b1000101011: data <= 21'h1ffe75; 
        10'b1000101100: data <= 21'h0001ab; 
        10'b1000101101: data <= 21'h1ffd73; 
        10'b1000101110: data <= 21'h1ff9fe; 
        10'b1000101111: data <= 21'h000214; 
        10'b1000110000: data <= 21'h00020b; 
        10'b1000110001: data <= 21'h0002b7; 
        10'b1000110010: data <= 21'h1ffe0f; 
        10'b1000110011: data <= 21'h1ffb8a; 
        10'b1000110100: data <= 21'h1ffd58; 
        10'b1000110101: data <= 21'h000bf8; 
        10'b1000110110: data <= 21'h00166a; 
        10'b1000110111: data <= 21'h001082; 
        10'b1000111000: data <= 21'h001476; 
        10'b1000111001: data <= 21'h001922; 
        10'b1000111010: data <= 21'h00272f; 
        10'b1000111011: data <= 21'h002722; 
        10'b1000111100: data <= 21'h001399; 
        10'b1000111101: data <= 21'h0005fb; 
        10'b1000111110: data <= 21'h1ffbef; 
        10'b1000111111: data <= 21'h0002d0; 
        10'b1001000000: data <= 21'h0002aa; 
        10'b1001000001: data <= 21'h1ffa49; 
        10'b1001000010: data <= 21'h1ffbaa; 
        10'b1001000011: data <= 21'h1ff9ea; 
        10'b1001000100: data <= 21'h00033d; 
        10'b1001000101: data <= 21'h000402; 
        10'b1001000110: data <= 21'h00062a; 
        10'b1001000111: data <= 21'h000224; 
        10'b1001001000: data <= 21'h1ffc8e; 
        10'b1001001001: data <= 21'h1fff37; 
        10'b1001001010: data <= 21'h1ffb28; 
        10'b1001001011: data <= 21'h1ffd7b; 
        10'b1001001100: data <= 21'h1ffc67; 
        10'b1001001101: data <= 21'h1ffaad; 
        10'b1001001110: data <= 21'h1ffe1a; 
        10'b1001001111: data <= 21'h1ffc7c; 
        10'b1001010000: data <= 21'h1ffdc3; 
        10'b1001010001: data <= 21'h00031a; 
        10'b1001010010: data <= 21'h000dd9; 
        10'b1001010011: data <= 21'h001688; 
        10'b1001010100: data <= 21'h000fce; 
        10'b1001010101: data <= 21'h001124; 
        10'b1001010110: data <= 21'h00218b; 
        10'b1001010111: data <= 21'h0025ec; 
        10'b1001011000: data <= 21'h001926; 
        10'b1001011001: data <= 21'h000984; 
        10'b1001011010: data <= 21'h00038b; 
        10'b1001011011: data <= 21'h0000bd; 
        10'b1001011100: data <= 21'h1fff61; 
        10'b1001011101: data <= 21'h1ff5a0; 
        10'b1001011110: data <= 21'h1ff815; 
        10'b1001011111: data <= 21'h1ffb72; 
        10'b1001100000: data <= 21'h0003f4; 
        10'b1001100001: data <= 21'h1fffb6; 
        10'b1001100010: data <= 21'h1ffb4d; 
        10'b1001100011: data <= 21'h1ff879; 
        10'b1001100100: data <= 21'h1ffe27; 
        10'b1001100101: data <= 21'h1ffd87; 
        10'b1001100110: data <= 21'h1ffc58; 
        10'b1001100111: data <= 21'h1ffcdf; 
        10'b1001101000: data <= 21'h1ffb87; 
        10'b1001101001: data <= 21'h000044; 
        10'b1001101010: data <= 21'h00006b; 
        10'b1001101011: data <= 21'h1ffd5b; 
        10'b1001101100: data <= 21'h1ffb46; 
        10'b1001101101: data <= 21'h0001be; 
        10'b1001101110: data <= 21'h000a12; 
        10'b1001101111: data <= 21'h0008bf; 
        10'b1001110000: data <= 21'h001947; 
        10'b1001110001: data <= 21'h00148d; 
        10'b1001110010: data <= 21'h0016a7; 
        10'b1001110011: data <= 21'h001af1; 
        10'b1001110100: data <= 21'h0016fb; 
        10'b1001110101: data <= 21'h001d88; 
        10'b1001110110: data <= 21'h000cca; 
        10'b1001110111: data <= 21'h000d17; 
        10'b1001111000: data <= 21'h000728; 
        10'b1001111001: data <= 21'h1ff9ec; 
        10'b1001111010: data <= 21'h1ffb29; 
        10'b1001111011: data <= 21'h1fffa8; 
        10'b1001111100: data <= 21'h1ff929; 
        10'b1001111101: data <= 21'h1ff8d5; 
        10'b1001111110: data <= 21'h1ffc8f; 
        10'b1001111111: data <= 21'h1ffc45; 
        10'b1010000000: data <= 21'h1ffeac; 
        10'b1010000001: data <= 21'h1ffdb3; 
        10'b1010000010: data <= 21'h1ffd06; 
        10'b1010000011: data <= 21'h1ffe6f; 
        10'b1010000100: data <= 21'h1ffb80; 
        10'b1010000101: data <= 21'h1ffec9; 
        10'b1010000110: data <= 21'h1fffe1; 
        10'b1010000111: data <= 21'h1ffa93; 
        10'b1010001000: data <= 21'h1ffa70; 
        10'b1010001001: data <= 21'h1ffe65; 
        10'b1010001010: data <= 21'h1fff56; 
        10'b1010001011: data <= 21'h0006fe; 
        10'b1010001100: data <= 21'h0009e2; 
        10'b1010001101: data <= 21'h001770; 
        10'b1010001110: data <= 21'h001c09; 
        10'b1010001111: data <= 21'h00224b; 
        10'b1010010000: data <= 21'h0021f2; 
        10'b1010010001: data <= 21'h00145a; 
        10'b1010010010: data <= 21'h001093; 
        10'b1010010011: data <= 21'h000929; 
        10'b1010010100: data <= 21'h0003df; 
        10'b1010010101: data <= 21'h1fff9f; 
        10'b1010010110: data <= 21'h1ff317; 
        10'b1010010111: data <= 21'h1fefcd; 
        10'b1010011000: data <= 21'h1ff373; 
        10'b1010011001: data <= 21'h1ff9cd; 
        10'b1010011010: data <= 21'h1ffaf8; 
        10'b1010011011: data <= 21'h1fff5a; 
        10'b1010011100: data <= 21'h1ffe14; 
        10'b1010011101: data <= 21'h000191; 
        10'b1010011110: data <= 21'h1ffd4e; 
        10'b1010011111: data <= 21'h1ffa5c; 
        10'b1010100000: data <= 21'h1ffd7d; 
        10'b1010100001: data <= 21'h1ffee4; 
        10'b1010100010: data <= 21'h1ffa70; 
        10'b1010100011: data <= 21'h1fffc7; 
        10'b1010100100: data <= 21'h1ffe7c; 
        10'b1010100101: data <= 21'h1ffe8d; 
        10'b1010100110: data <= 21'h1ff952; 
        10'b1010100111: data <= 21'h1ff718; 
        10'b1010101000: data <= 21'h1ffb0c; 
        10'b1010101001: data <= 21'h1ffb8e; 
        10'b1010101010: data <= 21'h00052f; 
        10'b1010101011: data <= 21'h0003e9; 
        10'b1010101100: data <= 21'h00097a; 
        10'b1010101101: data <= 21'h000dde; 
        10'b1010101110: data <= 21'h000752; 
        10'b1010101111: data <= 21'h1ffa6e; 
        10'b1010110000: data <= 21'h1ff75a; 
        10'b1010110001: data <= 21'h1ff5ab; 
        10'b1010110010: data <= 21'h1ff733; 
        10'b1010110011: data <= 21'h1ff3a7; 
        10'b1010110100: data <= 21'h1ff439; 
        10'b1010110101: data <= 21'h1ff4e0; 
        10'b1010110110: data <= 21'h1ffdd2; 
        10'b1010110111: data <= 21'h1ffd16; 
        10'b1010111000: data <= 21'h1ffb53; 
        10'b1010111001: data <= 21'h1ffc8f; 
        10'b1010111010: data <= 21'h000046; 
        10'b1010111011: data <= 21'h1ffbf1; 
        10'b1010111100: data <= 21'h1ffc99; 
        10'b1010111101: data <= 21'h00032d; 
        10'b1010111110: data <= 21'h1ffe50; 
        10'b1010111111: data <= 21'h0002a5; 
        10'b1011000000: data <= 21'h000303; 
        10'b1011000001: data <= 21'h1fffda; 
        10'b1011000010: data <= 21'h1ff9fc; 
        10'b1011000011: data <= 21'h1ffd5e; 
        10'b1011000100: data <= 21'h1ff449; 
        10'b1011000101: data <= 21'h1ff4e8; 
        10'b1011000110: data <= 21'h1ff237; 
        10'b1011000111: data <= 21'h1fee1a; 
        10'b1011001000: data <= 21'h1feb8a; 
        10'b1011001001: data <= 21'h1fed60; 
        10'b1011001010: data <= 21'h1fea4d; 
        10'b1011001011: data <= 21'h1fec6e; 
        10'b1011001100: data <= 21'h1fed80; 
        10'b1011001101: data <= 21'h1ff4df; 
        10'b1011001110: data <= 21'h1ff6c7; 
        10'b1011001111: data <= 21'h1ff832; 
        10'b1011010000: data <= 21'h1ff75a; 
        10'b1011010001: data <= 21'h1ff807; 
        10'b1011010010: data <= 21'h1ffd54; 
        10'b1011010011: data <= 21'h0002ff; 
        10'b1011010100: data <= 21'h000178; 
        10'b1011010101: data <= 21'h1ffddd; 
        10'b1011010110: data <= 21'h1ffd25; 
        10'b1011010111: data <= 21'h1ffeea; 
        10'b1011011000: data <= 21'h000285; 
        10'b1011011001: data <= 21'h000243; 
        10'b1011011010: data <= 21'h1ffdb4; 
        10'b1011011011: data <= 21'h000025; 
        10'b1011011100: data <= 21'h1ffcdc; 
        10'b1011011101: data <= 21'h1ffd78; 
        10'b1011011110: data <= 21'h1ffa94; 
        10'b1011011111: data <= 21'h000113; 
        10'b1011100000: data <= 21'h1ffd1f; 
        10'b1011100001: data <= 21'h1ff62f; 
        10'b1011100010: data <= 21'h1ff628; 
        10'b1011100011: data <= 21'h1ff717; 
        10'b1011100100: data <= 21'h1ffc68; 
        10'b1011100101: data <= 21'h1ff71b; 
        10'b1011100110: data <= 21'h1ff78f; 
        10'b1011100111: data <= 21'h1ffcdb; 
        10'b1011101000: data <= 21'h1ff702; 
        10'b1011101001: data <= 21'h1ff8b0; 
        10'b1011101010: data <= 21'h1ffa8d; 
        10'b1011101011: data <= 21'h1ff923; 
        10'b1011101100: data <= 21'h1ffc94; 
        10'b1011101101: data <= 21'h1ff7c3; 
        10'b1011101110: data <= 21'h1ff90b; 
        10'b1011101111: data <= 21'h0002b4; 
        10'b1011110000: data <= 21'h1ffbbf; 
        10'b1011110001: data <= 21'h0000ca; 
        10'b1011110010: data <= 21'h00023e; 
        10'b1011110011: data <= 21'h1fff7e; 
        10'b1011110100: data <= 21'h1ffb5c; 
        10'b1011110101: data <= 21'h0001dd; 
        10'b1011110110: data <= 21'h1fff36; 
        10'b1011110111: data <= 21'h1ffd7f; 
        10'b1011111000: data <= 21'h000260; 
        10'b1011111001: data <= 21'h000077; 
        10'b1011111010: data <= 21'h0000d5; 
        10'b1011111011: data <= 21'h1ffa50; 
        10'b1011111100: data <= 21'h0002c9; 
        10'b1011111101: data <= 21'h0002b8; 
        10'b1011111110: data <= 21'h0000f1; 
        10'b1011111111: data <= 21'h0001f5; 
        10'b1100000000: data <= 21'h1ffea6; 
        10'b1100000001: data <= 21'h1ffca3; 
        10'b1100000010: data <= 21'h0001da; 
        10'b1100000011: data <= 21'h1ffb1d; 
        10'b1100000100: data <= 21'h1ffe33; 
        10'b1100000101: data <= 21'h1ffc91; 
        10'b1100000110: data <= 21'h1fff2a; 
        10'b1100000111: data <= 21'h1ffcf7; 
        10'b1100001000: data <= 21'h1ffa33; 
        10'b1100001001: data <= 21'h1ffacd; 
        10'b1100001010: data <= 21'h1ff898; 
        10'b1100001011: data <= 21'h1ffe48; 
        10'b1100001100: data <= 21'h000132; 
        10'b1100001101: data <= 21'h1ffb4d; 
        10'b1100001110: data <= 21'h1ffa17; 
        10'b1100001111: data <= 21'h00018e; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 16) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 22'h3ff7b7; 
        10'b0000000001: data <= 22'h0004bd; 
        10'b0000000010: data <= 22'h3ffd6d; 
        10'b0000000011: data <= 22'h3ffecc; 
        10'b0000000100: data <= 22'h000591; 
        10'b0000000101: data <= 22'h3fff6c; 
        10'b0000000110: data <= 22'h3ffabe; 
        10'b0000000111: data <= 22'h3ffa65; 
        10'b0000001000: data <= 22'h3ffeb7; 
        10'b0000001001: data <= 22'h3ffd3c; 
        10'b0000001010: data <= 22'h000634; 
        10'b0000001011: data <= 22'h3fff82; 
        10'b0000001100: data <= 22'h0002d8; 
        10'b0000001101: data <= 22'h3ff7ee; 
        10'b0000001110: data <= 22'h3fff8c; 
        10'b0000001111: data <= 22'h3ff4ea; 
        10'b0000010000: data <= 22'h3ff6c6; 
        10'b0000010001: data <= 22'h3ffd89; 
        10'b0000010010: data <= 22'h3ff682; 
        10'b0000010011: data <= 22'h00062b; 
        10'b0000010100: data <= 22'h3ff6b8; 
        10'b0000010101: data <= 22'h3ffd09; 
        10'b0000010110: data <= 22'h3ff602; 
        10'b0000010111: data <= 22'h3fff00; 
        10'b0000011000: data <= 22'h000316; 
        10'b0000011001: data <= 22'h3ffdcb; 
        10'b0000011010: data <= 22'h3fff89; 
        10'b0000011011: data <= 22'h3fffb0; 
        10'b0000011100: data <= 22'h000384; 
        10'b0000011101: data <= 22'h000452; 
        10'b0000011110: data <= 22'h00016c; 
        10'b0000011111: data <= 22'h3ff644; 
        10'b0000100000: data <= 22'h3ff5c9; 
        10'b0000100001: data <= 22'h000088; 
        10'b0000100010: data <= 22'h3ff7ec; 
        10'b0000100011: data <= 22'h3ffdbf; 
        10'b0000100100: data <= 22'h3ff9be; 
        10'b0000100101: data <= 22'h3ff494; 
        10'b0000100110: data <= 22'h3ff8b6; 
        10'b0000100111: data <= 22'h000098; 
        10'b0000101000: data <= 22'h0006f3; 
        10'b0000101001: data <= 22'h3ff679; 
        10'b0000101010: data <= 22'h3ffad8; 
        10'b0000101011: data <= 22'h000303; 
        10'b0000101100: data <= 22'h3ff819; 
        10'b0000101101: data <= 22'h3ff53c; 
        10'b0000101110: data <= 22'h000205; 
        10'b0000101111: data <= 22'h0004d2; 
        10'b0000110000: data <= 22'h3ff7b5; 
        10'b0000110001: data <= 22'h000242; 
        10'b0000110010: data <= 22'h3ff8fc; 
        10'b0000110011: data <= 22'h3ff717; 
        10'b0000110100: data <= 22'h3ffe3d; 
        10'b0000110101: data <= 22'h000097; 
        10'b0000110110: data <= 22'h3ffd2e; 
        10'b0000110111: data <= 22'h0005ff; 
        10'b0000111000: data <= 22'h3ff5a3; 
        10'b0000111001: data <= 22'h3ff9a2; 
        10'b0000111010: data <= 22'h3ff909; 
        10'b0000111011: data <= 22'h0002f0; 
        10'b0000111100: data <= 22'h0000ce; 
        10'b0000111101: data <= 22'h3ff54d; 
        10'b0000111110: data <= 22'h3ffd71; 
        10'b0000111111: data <= 22'h0005b8; 
        10'b0001000000: data <= 22'h3ffc8b; 
        10'b0001000001: data <= 22'h3ff853; 
        10'b0001000010: data <= 22'h3ff89e; 
        10'b0001000011: data <= 22'h3ff35c; 
        10'b0001000100: data <= 22'h3ff28b; 
        10'b0001000101: data <= 22'h3ffb5b; 
        10'b0001000110: data <= 22'h3ff20f; 
        10'b0001000111: data <= 22'h3fee1c; 
        10'b0001001000: data <= 22'h3ff2f3; 
        10'b0001001001: data <= 22'h3ffc95; 
        10'b0001001010: data <= 22'h3ff4e9; 
        10'b0001001011: data <= 22'h3ff1b7; 
        10'b0001001100: data <= 22'h3ffd8a; 
        10'b0001001101: data <= 22'h00044f; 
        10'b0001001110: data <= 22'h0000c9; 
        10'b0001001111: data <= 22'h3ff81c; 
        10'b0001010000: data <= 22'h000563; 
        10'b0001010001: data <= 22'h3ff4a0; 
        10'b0001010010: data <= 22'h3ffd3c; 
        10'b0001010011: data <= 22'h000299; 
        10'b0001010100: data <= 22'h3ff55b; 
        10'b0001010101: data <= 22'h3ffd7f; 
        10'b0001010110: data <= 22'h000602; 
        10'b0001010111: data <= 22'h3ff5a6; 
        10'b0001011000: data <= 22'h3ff892; 
        10'b0001011001: data <= 22'h0004de; 
        10'b0001011010: data <= 22'h0001f5; 
        10'b0001011011: data <= 22'h000038; 
        10'b0001011100: data <= 22'h0000c8; 
        10'b0001011101: data <= 22'h3ffd46; 
        10'b0001011110: data <= 22'h3ffc66; 
        10'b0001011111: data <= 22'h3ff1e7; 
        10'b0001100000: data <= 22'h3fecb1; 
        10'b0001100001: data <= 22'h3ff511; 
        10'b0001100010: data <= 22'h3ff0e5; 
        10'b0001100011: data <= 22'h3feee7; 
        10'b0001100100: data <= 22'h0002d8; 
        10'b0001100101: data <= 22'h00015f; 
        10'b0001100110: data <= 22'h3fecf3; 
        10'b0001100111: data <= 22'h3fefb2; 
        10'b0001101000: data <= 22'h3fe8aa; 
        10'b0001101001: data <= 22'h3fef6c; 
        10'b0001101010: data <= 22'h3febff; 
        10'b0001101011: data <= 22'h3ff21c; 
        10'b0001101100: data <= 22'h3ff65d; 
        10'b0001101101: data <= 22'h0003a8; 
        10'b0001101110: data <= 22'h00038a; 
        10'b0001101111: data <= 22'h3ffa7d; 
        10'b0001110000: data <= 22'h000163; 
        10'b0001110001: data <= 22'h3ff532; 
        10'b0001110010: data <= 22'h3ff866; 
        10'b0001110011: data <= 22'h3ff572; 
        10'b0001110100: data <= 22'h3ff412; 
        10'b0001110101: data <= 22'h3ffe70; 
        10'b0001110110: data <= 22'h3ffcc2; 
        10'b0001110111: data <= 22'h3ff54f; 
        10'b0001111000: data <= 22'h3ffc64; 
        10'b0001111001: data <= 22'h3ffdb0; 
        10'b0001111010: data <= 22'h3feeaf; 
        10'b0001111011: data <= 22'h3feee1; 
        10'b0001111100: data <= 22'h3fef27; 
        10'b0001111101: data <= 22'h3fefec; 
        10'b0001111110: data <= 22'h3ffb9e; 
        10'b0001111111: data <= 22'h3ffe48; 
        10'b0010000000: data <= 22'h3ff2bc; 
        10'b0010000001: data <= 22'h3ff38c; 
        10'b0010000010: data <= 22'h3ff32a; 
        10'b0010000011: data <= 22'h3fee15; 
        10'b0010000100: data <= 22'h3ff8b5; 
        10'b0010000101: data <= 22'h3fe8f3; 
        10'b0010000110: data <= 22'h3ff707; 
        10'b0010000111: data <= 22'h3ffebf; 
        10'b0010001000: data <= 22'h3ff5f5; 
        10'b0010001001: data <= 22'h3ffb79; 
        10'b0010001010: data <= 22'h3ffa1a; 
        10'b0010001011: data <= 22'h3fff08; 
        10'b0010001100: data <= 22'h0002d5; 
        10'b0010001101: data <= 22'h3ffae9; 
        10'b0010001110: data <= 22'h3fffc1; 
        10'b0010001111: data <= 22'h3ff686; 
        10'b0010010000: data <= 22'h3ffd6e; 
        10'b0010010001: data <= 22'h3ffb60; 
        10'b0010010010: data <= 22'h3ffc9e; 
        10'b0010010011: data <= 22'h3ff8d5; 
        10'b0010010100: data <= 22'h3ffcc0; 
        10'b0010010101: data <= 22'h3ff313; 
        10'b0010010110: data <= 22'h3ffa2d; 
        10'b0010010111: data <= 22'h0003cf; 
        10'b0010011000: data <= 22'h000f1f; 
        10'b0010011001: data <= 22'h0020a9; 
        10'b0010011010: data <= 22'h002778; 
        10'b0010011011: data <= 22'h002706; 
        10'b0010011100: data <= 22'h002be5; 
        10'b0010011101: data <= 22'h002f3c; 
        10'b0010011110: data <= 22'h0031fa; 
        10'b0010011111: data <= 22'h00119e; 
        10'b0010100000: data <= 22'h000320; 
        10'b0010100001: data <= 22'h000821; 
        10'b0010100010: data <= 22'h3ffbf7; 
        10'b0010100011: data <= 22'h3fff6e; 
        10'b0010100100: data <= 22'h3feaab; 
        10'b0010100101: data <= 22'h3ff082; 
        10'b0010100110: data <= 22'h3ffee8; 
        10'b0010100111: data <= 22'h3ff7c0; 
        10'b0010101000: data <= 22'h3ffbb5; 
        10'b0010101001: data <= 22'h3ffdff; 
        10'b0010101010: data <= 22'h000127; 
        10'b0010101011: data <= 22'h3ffc75; 
        10'b0010101100: data <= 22'h00002a; 
        10'b0010101101: data <= 22'h000089; 
        10'b0010101110: data <= 22'h000138; 
        10'b0010101111: data <= 22'h3fff84; 
        10'b0010110000: data <= 22'h3ff54c; 
        10'b0010110001: data <= 22'h3fedcd; 
        10'b0010110010: data <= 22'h0009f4; 
        10'b0010110011: data <= 22'h3ffe70; 
        10'b0010110100: data <= 22'h001b11; 
        10'b0010110101: data <= 22'h0017f6; 
        10'b0010110110: data <= 22'h0016e0; 
        10'b0010110111: data <= 22'h0021f2; 
        10'b0010111000: data <= 22'h002962; 
        10'b0010111001: data <= 22'h003aa3; 
        10'b0010111010: data <= 22'h00368e; 
        10'b0010111011: data <= 22'h002e84; 
        10'b0010111100: data <= 22'h002ce0; 
        10'b0010111101: data <= 22'h003338; 
        10'b0010111110: data <= 22'h001d05; 
        10'b0010111111: data <= 22'h000a60; 
        10'b0011000000: data <= 22'h3fe9c4; 
        10'b0011000001: data <= 22'h3fe8d9; 
        10'b0011000010: data <= 22'h3ff057; 
        10'b0011000011: data <= 22'h000258; 
        10'b0011000100: data <= 22'h00055c; 
        10'b0011000101: data <= 22'h0000de; 
        10'b0011000110: data <= 22'h3ffee5; 
        10'b0011000111: data <= 22'h3ff25a; 
        10'b0011001000: data <= 22'h3feadc; 
        10'b0011001001: data <= 22'h3ffe22; 
        10'b0011001010: data <= 22'h3ff77d; 
        10'b0011001011: data <= 22'h000028; 
        10'b0011001100: data <= 22'h3ff615; 
        10'b0011001101: data <= 22'h3ffd15; 
        10'b0011001110: data <= 22'h0001e4; 
        10'b0011001111: data <= 22'h001355; 
        10'b0011010000: data <= 22'h00283c; 
        10'b0011010001: data <= 22'h00250b; 
        10'b0011010010: data <= 22'h000f2f; 
        10'b0011010011: data <= 22'h0017a0; 
        10'b0011010100: data <= 22'h0021bc; 
        10'b0011010101: data <= 22'h003ef7; 
        10'b0011010110: data <= 22'h002e57; 
        10'b0011010111: data <= 22'h00288d; 
        10'b0011011000: data <= 22'h001092; 
        10'b0011011001: data <= 22'h001fd1; 
        10'b0011011010: data <= 22'h0022f7; 
        10'b0011011011: data <= 22'h0011e1; 
        10'b0011011100: data <= 22'h3ff26e; 
        10'b0011011101: data <= 22'h3fe9bb; 
        10'b0011011110: data <= 22'h3fec01; 
        10'b0011011111: data <= 22'h3ffec6; 
        10'b0011100000: data <= 22'h000609; 
        10'b0011100001: data <= 22'h000235; 
        10'b0011100010: data <= 22'h3ffd70; 
        10'b0011100011: data <= 22'h3fffe5; 
        10'b0011100100: data <= 22'h3ff07c; 
        10'b0011100101: data <= 22'h3ff3f6; 
        10'b0011100110: data <= 22'h3ff61a; 
        10'b0011100111: data <= 22'h3ff3d4; 
        10'b0011101000: data <= 22'h3ff992; 
        10'b0011101001: data <= 22'h3ff940; 
        10'b0011101010: data <= 22'h001317; 
        10'b0011101011: data <= 22'h001415; 
        10'b0011101100: data <= 22'h000a4b; 
        10'b0011101101: data <= 22'h000451; 
        10'b0011101110: data <= 22'h000722; 
        10'b0011101111: data <= 22'h001c53; 
        10'b0011110000: data <= 22'h005298; 
        10'b0011110001: data <= 22'h0041bd; 
        10'b0011110010: data <= 22'h003d0a; 
        10'b0011110011: data <= 22'h001330; 
        10'b0011110100: data <= 22'h001024; 
        10'b0011110101: data <= 22'h000ec6; 
        10'b0011110110: data <= 22'h002435; 
        10'b0011110111: data <= 22'h003f17; 
        10'b0011111000: data <= 22'h3ff90d; 
        10'b0011111001: data <= 22'h3feb02; 
        10'b0011111010: data <= 22'h3ffdea; 
        10'b0011111011: data <= 22'h3ff4fb; 
        10'b0011111100: data <= 22'h3ffe4a; 
        10'b0011111101: data <= 22'h3ffef4; 
        10'b0011111110: data <= 22'h0001da; 
        10'b0011111111: data <= 22'h000161; 
        10'b0100000000: data <= 22'h3fec83; 
        10'b0100000001: data <= 22'h3ff21d; 
        10'b0100000010: data <= 22'h3fec14; 
        10'b0100000011: data <= 22'h3ff492; 
        10'b0100000100: data <= 22'h3ff4bb; 
        10'b0100000101: data <= 22'h3ffa39; 
        10'b0100000110: data <= 22'h000dbb; 
        10'b0100000111: data <= 22'h3ff445; 
        10'b0100001000: data <= 22'h0006d0; 
        10'b0100001001: data <= 22'h0014ae; 
        10'b0100001010: data <= 22'h001261; 
        10'b0100001011: data <= 22'h000fb0; 
        10'b0100001100: data <= 22'h002d3f; 
        10'b0100001101: data <= 22'h003c4a; 
        10'b0100001110: data <= 22'h004550; 
        10'b0100001111: data <= 22'h002818; 
        10'b0100010000: data <= 22'h000c34; 
        10'b0100010001: data <= 22'h3ffdbd; 
        10'b0100010010: data <= 22'h001dbd; 
        10'b0100010011: data <= 22'h00402d; 
        10'b0100010100: data <= 22'h0012b8; 
        10'b0100010101: data <= 22'h3ff034; 
        10'b0100010110: data <= 22'h00003a; 
        10'b0100010111: data <= 22'h3ffe0e; 
        10'b0100011000: data <= 22'h3ff5df; 
        10'b0100011001: data <= 22'h0004f5; 
        10'b0100011010: data <= 22'h3ff777; 
        10'b0100011011: data <= 22'h3ff07e; 
        10'b0100011100: data <= 22'h3ff1c7; 
        10'b0100011101: data <= 22'h3ff4bd; 
        10'b0100011110: data <= 22'h3ff676; 
        10'b0100011111: data <= 22'h000141; 
        10'b0100100000: data <= 22'h00068e; 
        10'b0100100001: data <= 22'h3ffe7a; 
        10'b0100100010: data <= 22'h3ff519; 
        10'b0100100011: data <= 22'h00038b; 
        10'b0100100100: data <= 22'h000473; 
        10'b0100100101: data <= 22'h3ffd6c; 
        10'b0100100110: data <= 22'h3fea3b; 
        10'b0100100111: data <= 22'h3fda90; 
        10'b0100101000: data <= 22'h3fe987; 
        10'b0100101001: data <= 22'h0015b7; 
        10'b0100101010: data <= 22'h003722; 
        10'b0100101011: data <= 22'h003920; 
        10'b0100101100: data <= 22'h00328f; 
        10'b0100101101: data <= 22'h0024a1; 
        10'b0100101110: data <= 22'h00364f; 
        10'b0100101111: data <= 22'h004a45; 
        10'b0100110000: data <= 22'h00235c; 
        10'b0100110001: data <= 22'h3ff16b; 
        10'b0100110010: data <= 22'h3ff15e; 
        10'b0100110011: data <= 22'h3ff4d1; 
        10'b0100110100: data <= 22'h3ff86c; 
        10'b0100110101: data <= 22'h3ff5df; 
        10'b0100110110: data <= 22'h000443; 
        10'b0100110111: data <= 22'h3ffcda; 
        10'b0100111000: data <= 22'h3fe421; 
        10'b0100111001: data <= 22'h3ffa0f; 
        10'b0100111010: data <= 22'h00045b; 
        10'b0100111011: data <= 22'h001507; 
        10'b0100111100: data <= 22'h000fcc; 
        10'b0100111101: data <= 22'h3ff9f3; 
        10'b0100111110: data <= 22'h000588; 
        10'b0100111111: data <= 22'h000090; 
        10'b0101000000: data <= 22'h000add; 
        10'b0101000001: data <= 22'h3ff89a; 
        10'b0101000010: data <= 22'h3fc4f0; 
        10'b0101000011: data <= 22'h3f9293; 
        10'b0101000100: data <= 22'h3f990c; 
        10'b0101000101: data <= 22'h3fd7c7; 
        10'b0101000110: data <= 22'h3ffaa3; 
        10'b0101000111: data <= 22'h001d0f; 
        10'b0101001000: data <= 22'h002e7e; 
        10'b0101001001: data <= 22'h002b0b; 
        10'b0101001010: data <= 22'h003ab3; 
        10'b0101001011: data <= 22'h00429c; 
        10'b0101001100: data <= 22'h002fe7; 
        10'b0101001101: data <= 22'h3ff6ca; 
        10'b0101001110: data <= 22'h3fff61; 
        10'b0101001111: data <= 22'h3ff427; 
        10'b0101010000: data <= 22'h3ff803; 
        10'b0101010001: data <= 22'h3ffd75; 
        10'b0101010010: data <= 22'h3ffc5a; 
        10'b0101010011: data <= 22'h3ffcf8; 
        10'b0101010100: data <= 22'h3ff049; 
        10'b0101010101: data <= 22'h000286; 
        10'b0101010110: data <= 22'h0016ea; 
        10'b0101010111: data <= 22'h0017f0; 
        10'b0101011000: data <= 22'h000b95; 
        10'b0101011001: data <= 22'h3ffcc9; 
        10'b0101011010: data <= 22'h00106f; 
        10'b0101011011: data <= 22'h000ba7; 
        10'b0101011100: data <= 22'h00157e; 
        10'b0101011101: data <= 22'h3fee57; 
        10'b0101011110: data <= 22'h3f8c18; 
        10'b0101011111: data <= 22'h3f706e; 
        10'b0101100000: data <= 22'h3f710f; 
        10'b0101100001: data <= 22'h3fb1da; 
        10'b0101100010: data <= 22'h3ff22a; 
        10'b0101100011: data <= 22'h3ffa44; 
        10'b0101100100: data <= 22'h000706; 
        10'b0101100101: data <= 22'h001403; 
        10'b0101100110: data <= 22'h004c22; 
        10'b0101100111: data <= 22'h0045a1; 
        10'b0101101000: data <= 22'h003060; 
        10'b0101101001: data <= 22'h0001ba; 
        10'b0101101010: data <= 22'h3ff863; 
        10'b0101101011: data <= 22'h3ff84b; 
        10'b0101101100: data <= 22'h3ff4a6; 
        10'b0101101101: data <= 22'h3fffbd; 
        10'b0101101110: data <= 22'h0003fe; 
        10'b0101101111: data <= 22'h3ff524; 
        10'b0101110000: data <= 22'h3ffbd7; 
        10'b0101110001: data <= 22'h000e37; 
        10'b0101110010: data <= 22'h001bc3; 
        10'b0101110011: data <= 22'h0023d9; 
        10'b0101110100: data <= 22'h001b1e; 
        10'b0101110101: data <= 22'h0012fe; 
        10'b0101110110: data <= 22'h0019ec; 
        10'b0101110111: data <= 22'h001425; 
        10'b0101111000: data <= 22'h000e87; 
        10'b0101111001: data <= 22'h3fb96c; 
        10'b0101111010: data <= 22'h3f8be4; 
        10'b0101111011: data <= 22'h3f6c75; 
        10'b0101111100: data <= 22'h3f86d9; 
        10'b0101111101: data <= 22'h3fc3db; 
        10'b0101111110: data <= 22'h3fe298; 
        10'b0101111111: data <= 22'h3fd88a; 
        10'b0110000000: data <= 22'h3fe1d4; 
        10'b0110000001: data <= 22'h000d40; 
        10'b0110000010: data <= 22'h0031f1; 
        10'b0110000011: data <= 22'h004e6c; 
        10'b0110000100: data <= 22'h002c85; 
        10'b0110000101: data <= 22'h00072c; 
        10'b0110000110: data <= 22'h00000d; 
        10'b0110000111: data <= 22'h000452; 
        10'b0110001000: data <= 22'h3ffe61; 
        10'b0110001001: data <= 22'h00036b; 
        10'b0110001010: data <= 22'h3ff74a; 
        10'b0110001011: data <= 22'h3ff9b2; 
        10'b0110001100: data <= 22'h3ff279; 
        10'b0110001101: data <= 22'h0024ad; 
        10'b0110001110: data <= 22'h002fa3; 
        10'b0110001111: data <= 22'h0039d8; 
        10'b0110010000: data <= 22'h001bc2; 
        10'b0110010001: data <= 22'h00215a; 
        10'b0110010010: data <= 22'h00310f; 
        10'b0110010011: data <= 22'h001c2d; 
        10'b0110010100: data <= 22'h0006e2; 
        10'b0110010101: data <= 22'h3fc292; 
        10'b0110010110: data <= 22'h3f7717; 
        10'b0110010111: data <= 22'h3f6c0b; 
        10'b0110011000: data <= 22'h3f8a49; 
        10'b0110011001: data <= 22'h3fbf9a; 
        10'b0110011010: data <= 22'h3fe3a8; 
        10'b0110011011: data <= 22'h3fddba; 
        10'b0110011100: data <= 22'h000311; 
        10'b0110011101: data <= 22'h001be7; 
        10'b0110011110: data <= 22'h00214f; 
        10'b0110011111: data <= 22'h004f3c; 
        10'b0110100000: data <= 22'h00293b; 
        10'b0110100001: data <= 22'h3ff7a9; 
        10'b0110100010: data <= 22'h3ffbdc; 
        10'b0110100011: data <= 22'h3ff719; 
        10'b0110100100: data <= 22'h00049c; 
        10'b0110100101: data <= 22'h000290; 
        10'b0110100110: data <= 22'h3ff877; 
        10'b0110100111: data <= 22'h3ffe43; 
        10'b0110101000: data <= 22'h3fff62; 
        10'b0110101001: data <= 22'h0033ce; 
        10'b0110101010: data <= 22'h002595; 
        10'b0110101011: data <= 22'h0033b9; 
        10'b0110101100: data <= 22'h0023b5; 
        10'b0110101101: data <= 22'h002f59; 
        10'b0110101110: data <= 22'h003bdf; 
        10'b0110101111: data <= 22'h001084; 
        10'b0110110000: data <= 22'h3fd2eb; 
        10'b0110110001: data <= 22'h3f8d1e; 
        10'b0110110010: data <= 22'h3f6691; 
        10'b0110110011: data <= 22'h3f6de9; 
        10'b0110110100: data <= 22'h3f9d51; 
        10'b0110110101: data <= 22'h3fcfd7; 
        10'b0110110110: data <= 22'h3fee07; 
        10'b0110110111: data <= 22'h3fee9b; 
        10'b0110111000: data <= 22'h000ef8; 
        10'b0110111001: data <= 22'h000d26; 
        10'b0110111010: data <= 22'h003252; 
        10'b0110111011: data <= 22'h003b27; 
        10'b0110111100: data <= 22'h001ea0; 
        10'b0110111101: data <= 22'h3ffcf9; 
        10'b0110111110: data <= 22'h0000e0; 
        10'b0110111111: data <= 22'h3ff7e9; 
        10'b0111000000: data <= 22'h000155; 
        10'b0111000001: data <= 22'h0005cc; 
        10'b0111000010: data <= 22'h3ff447; 
        10'b0111000011: data <= 22'h3ff9a9; 
        10'b0111000100: data <= 22'h0008be; 
        10'b0111000101: data <= 22'h002efd; 
        10'b0111000110: data <= 22'h003a65; 
        10'b0111000111: data <= 22'h002d29; 
        10'b0111001000: data <= 22'h001f5c; 
        10'b0111001001: data <= 22'h001f9e; 
        10'b0111001010: data <= 22'h003550; 
        10'b0111001011: data <= 22'h3ff900; 
        10'b0111001100: data <= 22'h3fa872; 
        10'b0111001101: data <= 22'h3f67ba; 
        10'b0111001110: data <= 22'h3f6bb2; 
        10'b0111001111: data <= 22'h3f8a5c; 
        10'b0111010000: data <= 22'h3fc0fd; 
        10'b0111010001: data <= 22'h3fe293; 
        10'b0111010010: data <= 22'h3fff9d; 
        10'b0111010011: data <= 22'h0009a6; 
        10'b0111010100: data <= 22'h00162c; 
        10'b0111010101: data <= 22'h0020f4; 
        10'b0111010110: data <= 22'h002d52; 
        10'b0111010111: data <= 22'h002b43; 
        10'b0111011000: data <= 22'h001075; 
        10'b0111011001: data <= 22'h0000cd; 
        10'b0111011010: data <= 22'h3ffaa1; 
        10'b0111011011: data <= 22'h3ff8c2; 
        10'b0111011100: data <= 22'h3ffbc9; 
        10'b0111011101: data <= 22'h00016d; 
        10'b0111011110: data <= 22'h3ff618; 
        10'b0111011111: data <= 22'h3fecc0; 
        10'b0111100000: data <= 22'h0001a3; 
        10'b0111100001: data <= 22'h002161; 
        10'b0111100010: data <= 22'h0029e1; 
        10'b0111100011: data <= 22'h0028b6; 
        10'b0111100100: data <= 22'h000cb3; 
        10'b0111100101: data <= 22'h0020b0; 
        10'b0111100110: data <= 22'h0033a8; 
        10'b0111100111: data <= 22'h3ff818; 
        10'b0111101000: data <= 22'h3f971b; 
        10'b0111101001: data <= 22'h3f69ca; 
        10'b0111101010: data <= 22'h3f7bc0; 
        10'b0111101011: data <= 22'h3fb12b; 
        10'b0111101100: data <= 22'h3ff5a6; 
        10'b0111101101: data <= 22'h001418; 
        10'b0111101110: data <= 22'h001cf6; 
        10'b0111101111: data <= 22'h001ab1; 
        10'b0111110000: data <= 22'h00220c; 
        10'b0111110001: data <= 22'h0019f5; 
        10'b0111110010: data <= 22'h001485; 
        10'b0111110011: data <= 22'h00174c; 
        10'b0111110100: data <= 22'h3ffec0; 
        10'b0111110101: data <= 22'h3ffc8b; 
        10'b0111110110: data <= 22'h0001d0; 
        10'b0111110111: data <= 22'h3ff7df; 
        10'b0111111000: data <= 22'h3ffa62; 
        10'b0111111001: data <= 22'h0001d0; 
        10'b0111111010: data <= 22'h3ffc12; 
        10'b0111111011: data <= 22'h3ff8a1; 
        10'b0111111100: data <= 22'h3ffbf6; 
        10'b0111111101: data <= 22'h00154d; 
        10'b0111111110: data <= 22'h002b69; 
        10'b0111111111: data <= 22'h001911; 
        10'b1000000000: data <= 22'h000f66; 
        10'b1000000001: data <= 22'h002b2c; 
        10'b1000000010: data <= 22'h0052cb; 
        10'b1000000011: data <= 22'h000342; 
        10'b1000000100: data <= 22'h3fbd2a; 
        10'b1000000101: data <= 22'h3f942e; 
        10'b1000000110: data <= 22'h3fb4d2; 
        10'b1000000111: data <= 22'h3fe915; 
        10'b1000001000: data <= 22'h001843; 
        10'b1000001001: data <= 22'h0019e7; 
        10'b1000001010: data <= 22'h001b18; 
        10'b1000001011: data <= 22'h000e1d; 
        10'b1000001100: data <= 22'h000708; 
        10'b1000001101: data <= 22'h000bbd; 
        10'b1000001110: data <= 22'h001693; 
        10'b1000001111: data <= 22'h000e13; 
        10'b1000010000: data <= 22'h3ffe46; 
        10'b1000010001: data <= 22'h3ff916; 
        10'b1000010010: data <= 22'h0000d5; 
        10'b1000010011: data <= 22'h3ffc19; 
        10'b1000010100: data <= 22'h3ffc8a; 
        10'b1000010101: data <= 22'h3ffb29; 
        10'b1000010110: data <= 22'h3ffbab; 
        10'b1000010111: data <= 22'h3fed3c; 
        10'b1000011000: data <= 22'h00080a; 
        10'b1000011001: data <= 22'h00175c; 
        10'b1000011010: data <= 22'h0037c5; 
        10'b1000011011: data <= 22'h0032ad; 
        10'b1000011100: data <= 22'h0027a2; 
        10'b1000011101: data <= 22'h003499; 
        10'b1000011110: data <= 22'h0052fa; 
        10'b1000011111: data <= 22'h003a5b; 
        10'b1000100000: data <= 22'h000c55; 
        10'b1000100001: data <= 22'h3fe52c; 
        10'b1000100010: data <= 22'h3ff446; 
        10'b1000100011: data <= 22'h3ff87e; 
        10'b1000100100: data <= 22'h000cb0; 
        10'b1000100101: data <= 22'h3ffa28; 
        10'b1000100110: data <= 22'h3ff539; 
        10'b1000100111: data <= 22'h3ff974; 
        10'b1000101000: data <= 22'h000d0d; 
        10'b1000101001: data <= 22'h000be1; 
        10'b1000101010: data <= 22'h00174e; 
        10'b1000101011: data <= 22'h3ffcea; 
        10'b1000101100: data <= 22'h000355; 
        10'b1000101101: data <= 22'h3ffae5; 
        10'b1000101110: data <= 22'h3ff3fb; 
        10'b1000101111: data <= 22'h000428; 
        10'b1000110000: data <= 22'h000415; 
        10'b1000110001: data <= 22'h00056e; 
        10'b1000110010: data <= 22'h3ffc1d; 
        10'b1000110011: data <= 22'h3ff714; 
        10'b1000110100: data <= 22'h3ffab0; 
        10'b1000110101: data <= 22'h0017ef; 
        10'b1000110110: data <= 22'h002cd5; 
        10'b1000110111: data <= 22'h002104; 
        10'b1000111000: data <= 22'h0028eb; 
        10'b1000111001: data <= 22'h003244; 
        10'b1000111010: data <= 22'h004e5d; 
        10'b1000111011: data <= 22'h004e44; 
        10'b1000111100: data <= 22'h002733; 
        10'b1000111101: data <= 22'h000bf5; 
        10'b1000111110: data <= 22'h3ff7df; 
        10'b1000111111: data <= 22'h0005a1; 
        10'b1001000000: data <= 22'h000554; 
        10'b1001000001: data <= 22'h3ff492; 
        10'b1001000010: data <= 22'h3ff754; 
        10'b1001000011: data <= 22'h3ff3d4; 
        10'b1001000100: data <= 22'h00067a; 
        10'b1001000101: data <= 22'h000804; 
        10'b1001000110: data <= 22'h000c54; 
        10'b1001000111: data <= 22'h000448; 
        10'b1001001000: data <= 22'h3ff91c; 
        10'b1001001001: data <= 22'h3ffe6f; 
        10'b1001001010: data <= 22'h3ff64f; 
        10'b1001001011: data <= 22'h3ffaf6; 
        10'b1001001100: data <= 22'h3ff8ce; 
        10'b1001001101: data <= 22'h3ff55a; 
        10'b1001001110: data <= 22'h3ffc35; 
        10'b1001001111: data <= 22'h3ff8f8; 
        10'b1001010000: data <= 22'h3ffb86; 
        10'b1001010001: data <= 22'h000634; 
        10'b1001010010: data <= 22'h001bb2; 
        10'b1001010011: data <= 22'h002d10; 
        10'b1001010100: data <= 22'h001f9c; 
        10'b1001010101: data <= 22'h002249; 
        10'b1001010110: data <= 22'h004316; 
        10'b1001010111: data <= 22'h004bd8; 
        10'b1001011000: data <= 22'h00324c; 
        10'b1001011001: data <= 22'h001308; 
        10'b1001011010: data <= 22'h000716; 
        10'b1001011011: data <= 22'h00017a; 
        10'b1001011100: data <= 22'h3ffec2; 
        10'b1001011101: data <= 22'h3feb3f; 
        10'b1001011110: data <= 22'h3ff02a; 
        10'b1001011111: data <= 22'h3ff6e3; 
        10'b1001100000: data <= 22'h0007e8; 
        10'b1001100001: data <= 22'h3fff6b; 
        10'b1001100010: data <= 22'h3ff69a; 
        10'b1001100011: data <= 22'h3ff0f2; 
        10'b1001100100: data <= 22'h3ffc4e; 
        10'b1001100101: data <= 22'h3ffb0e; 
        10'b1001100110: data <= 22'h3ff8b0; 
        10'b1001100111: data <= 22'h3ff9be; 
        10'b1001101000: data <= 22'h3ff70e; 
        10'b1001101001: data <= 22'h000089; 
        10'b1001101010: data <= 22'h0000d7; 
        10'b1001101011: data <= 22'h3ffab6; 
        10'b1001101100: data <= 22'h3ff68b; 
        10'b1001101101: data <= 22'h00037b; 
        10'b1001101110: data <= 22'h001423; 
        10'b1001101111: data <= 22'h00117d; 
        10'b1001110000: data <= 22'h00328d; 
        10'b1001110001: data <= 22'h00291a; 
        10'b1001110010: data <= 22'h002d4e; 
        10'b1001110011: data <= 22'h0035e2; 
        10'b1001110100: data <= 22'h002df6; 
        10'b1001110101: data <= 22'h003b11; 
        10'b1001110110: data <= 22'h001994; 
        10'b1001110111: data <= 22'h001a2e; 
        10'b1001111000: data <= 22'h000e50; 
        10'b1001111001: data <= 22'h3ff3d8; 
        10'b1001111010: data <= 22'h3ff652; 
        10'b1001111011: data <= 22'h3fff50; 
        10'b1001111100: data <= 22'h3ff252; 
        10'b1001111101: data <= 22'h3ff1aa; 
        10'b1001111110: data <= 22'h3ff91d; 
        10'b1001111111: data <= 22'h3ff889; 
        10'b1010000000: data <= 22'h3ffd58; 
        10'b1010000001: data <= 22'h3ffb65; 
        10'b1010000010: data <= 22'h3ffa0b; 
        10'b1010000011: data <= 22'h3ffcde; 
        10'b1010000100: data <= 22'h3ff701; 
        10'b1010000101: data <= 22'h3ffd92; 
        10'b1010000110: data <= 22'h3fffc2; 
        10'b1010000111: data <= 22'h3ff526; 
        10'b1010001000: data <= 22'h3ff4e1; 
        10'b1010001001: data <= 22'h3ffcc9; 
        10'b1010001010: data <= 22'h3ffeac; 
        10'b1010001011: data <= 22'h000dfd; 
        10'b1010001100: data <= 22'h0013c4; 
        10'b1010001101: data <= 22'h002ee0; 
        10'b1010001110: data <= 22'h003811; 
        10'b1010001111: data <= 22'h004496; 
        10'b1010010000: data <= 22'h0043e4; 
        10'b1010010001: data <= 22'h0028b4; 
        10'b1010010010: data <= 22'h002126; 
        10'b1010010011: data <= 22'h001251; 
        10'b1010010100: data <= 22'h0007bf; 
        10'b1010010101: data <= 22'h3fff3f; 
        10'b1010010110: data <= 22'h3fe62f; 
        10'b1010010111: data <= 22'h3fdf9a; 
        10'b1010011000: data <= 22'h3fe6e5; 
        10'b1010011001: data <= 22'h3ff399; 
        10'b1010011010: data <= 22'h3ff5ef; 
        10'b1010011011: data <= 22'h3ffeb4; 
        10'b1010011100: data <= 22'h3ffc29; 
        10'b1010011101: data <= 22'h000322; 
        10'b1010011110: data <= 22'h3ffa9d; 
        10'b1010011111: data <= 22'h3ff4b7; 
        10'b1010100000: data <= 22'h3ffafa; 
        10'b1010100001: data <= 22'h3ffdc8; 
        10'b1010100010: data <= 22'h3ff4e1; 
        10'b1010100011: data <= 22'h3fff8f; 
        10'b1010100100: data <= 22'h3ffcf7; 
        10'b1010100101: data <= 22'h3ffd1b; 
        10'b1010100110: data <= 22'h3ff2a4; 
        10'b1010100111: data <= 22'h3fee2f; 
        10'b1010101000: data <= 22'h3ff617; 
        10'b1010101001: data <= 22'h3ff71c; 
        10'b1010101010: data <= 22'h000a5e; 
        10'b1010101011: data <= 22'h0007d2; 
        10'b1010101100: data <= 22'h0012f4; 
        10'b1010101101: data <= 22'h001bbc; 
        10'b1010101110: data <= 22'h000ea5; 
        10'b1010101111: data <= 22'h3ff4dc; 
        10'b1010110000: data <= 22'h3feeb4; 
        10'b1010110001: data <= 22'h3feb56; 
        10'b1010110010: data <= 22'h3fee66; 
        10'b1010110011: data <= 22'h3fe74d; 
        10'b1010110100: data <= 22'h3fe871; 
        10'b1010110101: data <= 22'h3fe9c0; 
        10'b1010110110: data <= 22'h3ffba3; 
        10'b1010110111: data <= 22'h3ffa2d; 
        10'b1010111000: data <= 22'h3ff6a7; 
        10'b1010111001: data <= 22'h3ff91f; 
        10'b1010111010: data <= 22'h00008c; 
        10'b1010111011: data <= 22'h3ff7e2; 
        10'b1010111100: data <= 22'h3ff931; 
        10'b1010111101: data <= 22'h00065a; 
        10'b1010111110: data <= 22'h3ffc9f; 
        10'b1010111111: data <= 22'h00054b; 
        10'b1011000000: data <= 22'h000606; 
        10'b1011000001: data <= 22'h3fffb4; 
        10'b1011000010: data <= 22'h3ff3f8; 
        10'b1011000011: data <= 22'h3ffabd; 
        10'b1011000100: data <= 22'h3fe891; 
        10'b1011000101: data <= 22'h3fe9d1; 
        10'b1011000110: data <= 22'h3fe46e; 
        10'b1011000111: data <= 22'h3fdc34; 
        10'b1011001000: data <= 22'h3fd715; 
        10'b1011001001: data <= 22'h3fdabf; 
        10'b1011001010: data <= 22'h3fd49b; 
        10'b1011001011: data <= 22'h3fd8dc; 
        10'b1011001100: data <= 22'h3fdb00; 
        10'b1011001101: data <= 22'h3fe9bf; 
        10'b1011001110: data <= 22'h3fed8e; 
        10'b1011001111: data <= 22'h3ff065; 
        10'b1011010000: data <= 22'h3feeb5; 
        10'b1011010001: data <= 22'h3ff00f; 
        10'b1011010010: data <= 22'h3ffaa8; 
        10'b1011010011: data <= 22'h0005ff; 
        10'b1011010100: data <= 22'h0002ef; 
        10'b1011010101: data <= 22'h3ffbbb; 
        10'b1011010110: data <= 22'h3ffa4b; 
        10'b1011010111: data <= 22'h3ffdd3; 
        10'b1011011000: data <= 22'h00050a; 
        10'b1011011001: data <= 22'h000486; 
        10'b1011011010: data <= 22'h3ffb68; 
        10'b1011011011: data <= 22'h00004a; 
        10'b1011011100: data <= 22'h3ff9b9; 
        10'b1011011101: data <= 22'h3ffaf1; 
        10'b1011011110: data <= 22'h3ff529; 
        10'b1011011111: data <= 22'h000226; 
        10'b1011100000: data <= 22'h3ffa3e; 
        10'b1011100001: data <= 22'h3fec5d; 
        10'b1011100010: data <= 22'h3fec4f; 
        10'b1011100011: data <= 22'h3fee2f; 
        10'b1011100100: data <= 22'h3ff8d1; 
        10'b1011100101: data <= 22'h3fee36; 
        10'b1011100110: data <= 22'h3fef1e; 
        10'b1011100111: data <= 22'h3ff9b7; 
        10'b1011101000: data <= 22'h3fee03; 
        10'b1011101001: data <= 22'h3ff160; 
        10'b1011101010: data <= 22'h3ff51b; 
        10'b1011101011: data <= 22'h3ff246; 
        10'b1011101100: data <= 22'h3ff928; 
        10'b1011101101: data <= 22'h3fef87; 
        10'b1011101110: data <= 22'h3ff216; 
        10'b1011101111: data <= 22'h000568; 
        10'b1011110000: data <= 22'h3ff77d; 
        10'b1011110001: data <= 22'h000195; 
        10'b1011110010: data <= 22'h00047c; 
        10'b1011110011: data <= 22'h3ffefb; 
        10'b1011110100: data <= 22'h3ff6b9; 
        10'b1011110101: data <= 22'h0003b9; 
        10'b1011110110: data <= 22'h3ffe6c; 
        10'b1011110111: data <= 22'h3ffaff; 
        10'b1011111000: data <= 22'h0004c1; 
        10'b1011111001: data <= 22'h0000ee; 
        10'b1011111010: data <= 22'h0001a9; 
        10'b1011111011: data <= 22'h3ff4a0; 
        10'b1011111100: data <= 22'h000592; 
        10'b1011111101: data <= 22'h000570; 
        10'b1011111110: data <= 22'h0001e2; 
        10'b1011111111: data <= 22'h0003ea; 
        10'b1100000000: data <= 22'h3ffd4d; 
        10'b1100000001: data <= 22'h3ff946; 
        10'b1100000010: data <= 22'h0003b5; 
        10'b1100000011: data <= 22'h3ff63a; 
        10'b1100000100: data <= 22'h3ffc67; 
        10'b1100000101: data <= 22'h3ff922; 
        10'b1100000110: data <= 22'h3ffe54; 
        10'b1100000111: data <= 22'h3ff9ef; 
        10'b1100001000: data <= 22'h3ff467; 
        10'b1100001001: data <= 22'h3ff59a; 
        10'b1100001010: data <= 22'h3ff131; 
        10'b1100001011: data <= 22'h3ffc91; 
        10'b1100001100: data <= 22'h000265; 
        10'b1100001101: data <= 22'h3ff69b; 
        10'b1100001110: data <= 22'h3ff42e; 
        10'b1100001111: data <= 22'h00031c; 
      endcase 
    end 
  end 
endgenerate 
assign dout = data; 
endmodule
