logic [BITS - 1 : 0] arr_0_digit_7 [0 : WIDTH-1]= '{-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-688,912,496,368,-1072,-1456,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1504,2016,2016,2016,2016,1808,1120,1120,1120,1120,1120,1120,1120,1120,672,-1200,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-960,-208,-880,-208,560,1584,2016,1552,2016,2016,2016,1952,1616,2016,2016,192,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1760,-976,-1808,-960,-960,-960,-1088,-1696,1728,2016,-336,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-704,2000,1296,-1744,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1680,1680,2048,-704,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,16,2016,1760,-1328,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1088,1936,2016,-1040,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,80,2016,944,-1952,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1888,1232,1920,-1104,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-16,2016,864,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-832,1968,1792,-1120,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1728,1488,2016,608,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1984,1200,2016,1456,-1472,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1424,2016,2016,-800,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1536,1536,2016,-192,-2016,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,80,2016,2016,-1200,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1056,1824,2016,2016,-1200,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-96,2016,2016,1456,-1392,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-96,2016,1264,-1744,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,}; 
logic [BITS - 1 : 0] arr_1_digit_2 [0 : WIDTH-1]= '{-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-176,-32,688,2048,2048,352,-544,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,656,2000,2000,2000,2000,2000,2000,1440,-1552,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,656,2000,2000,2000,1360,224,768,2000,2000,-80,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1200,1952,2000,1312,-1520,-1840,-2048,-1936,1248,2000,192,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-800,1968,1312,-1632,-2048,-2048,-2048,-80,1920,2000,-992,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1536,-1744,-2048,-2048,-2048,-2048,1296,2000,2000,-992,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-160,1904,2000,1120,-1872,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-816,1904,2000,1648,-1024,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,0,2000,2000,256,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,768,1888,2000,496,-1840,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1632,1696,2000,1680,-1472,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1120,2000,2000,208,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-784,1920,2000,976,-1840,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1728,1152,2000,2000,208,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,96,2000,2000,720,-1840,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1920,2000,2000,-1632,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1920,2000,2000,-1344,-1712,-1712,-1712,-1712,-1952,-2048,-1952,-1712,-1712,-1440,352,352,352,304,-1872,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1920,2000,2000,2000,2000,2000,2000,2000,640,240,608,2000,2000,2000,2000,2000,2000,2000,-64,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,736,2000,2000,2000,2000,2000,2000,2000,2000,2000,2000,2000,1936,1904,1904,656,-160,-160,-1120,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-144,-64,-64,-64,608,2000,2000,2000,432,-64,-64,-1376,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,}; 
logic [BITS - 1 : 0] arr_2_digit_1 [0 : WIDTH-1]= '{-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1424,2016,-288,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-640,1984,-720,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,112,1808,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1312,1856,352,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-688,2016,-1024,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1184,1520,-1856,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1520,2016,1408,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-512,2016,1072,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,192,2016,-800,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1120,1744,1232,-1904,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-48,2048,592,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,688,2016,-736,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1648,1664,1392,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-112,2016,496,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,368,2016,224,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1600,2016,-976,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1056,1968,2016,-976,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,208,2016,1232,-1984,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1872,1392,2016,-96,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1952,1120,768,-1872,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,}; 
logic [BITS - 1 : 0] arr_3_digit_0 [0 : WIDTH-1]= '{-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1856,352,2000,1184,-1536,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1440,1968,1968,2000,-320,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1696,1104,1968,1968,2000,-320,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-272,992,1968,1968,1968,2000,656,-288,-1040,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,2000,1968,1968,1968,1968,2000,1968,1968,1472,-1216,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,864,2048,2000,2000,2000,2000,1696,1504,2000,2000,2000,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1024,1488,2000,1968,1968,1968,304,-800,-1040,0,1968,1968,-352,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1520,1648,1968,2000,1968,1472,144,-1872,-2048,-2048,-1536,1632,1968,1840,-224,-1952,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1440,1968,1968,2000,960,-1712,-2048,-2048,-2048,-2048,-2048,-288,1968,2000,1968,-1472,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1440,1968,1968,1168,-1552,-2048,-2048,-2048,-2048,-2048,-2048,-1536,1152,2000,1968,-1472,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1440,2000,2000,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1520,1184,2048,2000,576,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,192,1968,1968,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-288,1968,2000,1968,-1472,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1424,1968,1968,-2048,-2048,-2048,-2048,-2048,-2048,-1696,-1024,1648,1968,2000,1632,-1552,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1424,1968,1968,-2048,-2048,-2048,-2048,-2048,-2048,256,1968,1968,1968,1488,-1056,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1424,1968,1968,-2048,-2048,-2048,-2048,-2048,864,1488,1968,1968,1968,832,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1440,2000,2000,-864,-864,1600,2000,2000,2048,2000,2000,2000,2000,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-224,1968,1968,2000,1968,1968,1968,1968,2000,1968,1968,1968,304,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1536,1632,1968,2000,1968,1968,1968,1968,2000,1632,976,-1472,-1872,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1040,224,2000,1968,1968,1968,1968,2000,-320,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-880,736,1968,720,-896,-880,-1552,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,}; 
logic [BITS - 1 : 0] arr_4_digit_4 [0 : WIDTH-1]= '{-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1232,1536,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-912,-1568,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-96,1648,-2048,-2048,-2048,-2048,-2048,-2048,-2048,320,640,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1968,1072,1648,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-496,1312,-1856,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-928,1984,96,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-208,1984,-1696,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1312,1728,1424,-1840,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1024,1984,-1696,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,640,1904,-1184,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1744,2048,2000,-1696,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-688,1824,1328,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,208,2000,976,-1952,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,656,1984,-336,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1520,1664,1952,-976,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1792,1552,1984,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,96,1984,1328,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1680,1984,576,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,656,1984,624,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1888,1216,1296,-1744,-2048,-2048,-2048,-2048,-2048,-2048,-1680,2000,2000,-320,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,656,1984,1136,-672,-672,-672,-672,16,576,1072,1984,1984,-336,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1376,672,1872,1984,1984,1984,1984,1664,1648,1968,1984,1984,-1888,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1248,-688,-688,-688,-688,-2048,-2048,528,1984,1984,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,0,1984,1984,-1312,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,0,2000,2000,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,0,1984,1984,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,112,1984,1856,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1664,1728,-256,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,816,-976,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,}; 
logic [BITS - 1 : 0] arr_5_digit_1 [0 : WIDTH-1]= '{-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-800,2016,-320,-1984,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1728,1584,2016,2016,-1888,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-736,2016,2016,592,-2016,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1920,1200,2016,2016,-864,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1184,2016,2016,1952,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,96,2016,2016,832,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1088,2016,1920,-1264,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1104,2016,2016,1744,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-256,2016,2016,64,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,560,2016,1760,-1584,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1072,1984,2016,1520,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-768,2016,2016,416,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,560,2016,1760,-1184,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1584,1984,2016,1312,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-656,2016,2016,48,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-352,2016,1696,-1712,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,752,2016,1216,-1952,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1952,1328,2016,1088,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1984,480,2016,512,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1616,464,-320,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,}; 
logic [BITS - 1 : 0] arr_6_digit_4 [0 : WIDTH-1]= '{-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1680,1024,96,-1520,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1792,-800,-1952,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1760,1712,1952,656,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1792,1472,1808,-1440,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1712,976,2000,304,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,176,2000,-432,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-912,2000,2000,-1696,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1344,2016,720,-1824,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1680,400,2000,-496,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1344,1648,2016,-560,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,560,2048,1216,-1856,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-368,2016,480,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,544,2000,800,-1952,-2048,-2048,-2048,-2048,-2048,-2048,-1888,48,1744,2000,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,544,2000,2000,1008,752,-912,-912,-912,-912,80,1104,2000,2000,656,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1216,1600,2000,2000,2016,2000,2000,2000,2000,2016,2000,2000,1456,-1472,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1760,-992,144,2016,1664,144,144,144,-1328,2000,2000,528,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1488,2016,1248,-1696,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,512,2000,-928,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-672,2016,1808,-1232,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,480,2016,592,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1648,1856,-1232,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-368,2016,1664,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1280,2000,464,-2048,-1824,-1552,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1280,2000,416,-576,1216,528,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1280,2000,2016,2000,416,-1568,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1056,992,0,-1664,-1936,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,}; 
logic [BITS - 1 : 0] arr_7_digit_9 [0 : WIDTH-1]= '{-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1808,336,1040,-1952,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-576,1536,2000,2000,-1728,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1584,1712,2016,2000,2000,608,-1744,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,256,2000,2016,2000,2000,2000,1760,-192,-1936,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1536,1808,2000,1280,912,2000,2000,2000,1648,-1648,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-768,2016,1040,-2048,-1904,-464,1456,2016,2048,1168,-1744,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-656,2000,-752,-2048,-2048,-2048,864,2000,2016,1008,-1840,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,752,2000,432,-2048,-2048,-2048,1696,2000,2016,112,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-656,2000,1280,-1392,-672,608,1968,1744,2016,1728,-1360,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1744,1760,2000,2016,2000,2000,912,-1456,1408,2000,384,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-944,1792,2048,2016,272,-1904,-2048,96,2016,1520,-1472,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-944,480,224,-1840,-2048,-2048,-1888,752,2000,528,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-624,2000,1568,-1744,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2000,608,2000,-16,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1264,1872,2000,-1424,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-192,2016,704,-1888,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1696,1440,2016,-1296,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1552,2016,592,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,928,1856,-1360,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1808,1520,-784,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,}; 
logic [BITS - 1 : 0] arr_8_digit_5 [0 : WIDTH-1]= '{-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1760,-1280,-1280,-1280,-1776,16,-672,-1280,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-832,400,1424,2000,2000,2000,1392,1888,2000,2000,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1472,224,1856,1984,2000,2000,2000,2000,2000,2000,2000,2000,2000,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1024,2000,2000,2000,2000,2000,2000,2000,1360,672,672,672,672,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1712,64,-880,-2048,-1120,1760,1584,1760,640,-48,-928,-1712,-1856,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1856,1248,2000,-784,-2048,-2048,-1520,-2048,-1552,-2000,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1936,784,2000,64,-1872,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1840,80,2000,1680,-1792,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-560,2000,1520,-1584,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,352,2000,736,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1696,2000,1888,0,-1248,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,2048,2000,2000,2000,1968,304,-576,-96,-672,-1360,-1360,-672,-1584,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,176,2000,2000,2000,2000,2000,2000,2000,2000,2000,2000,2000,1664,640,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1984,-1184,1440,1504,1968,2000,2000,2000,2000,2000,2000,2000,2000,1984,-48,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-960,-880,1152,2000,2000,2000,2000,2000,2000,2000,752,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-112,2000,1936,384,-1216,576,2000,2000,752,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1232,2000,2000,2000,960,1984,2000,2000,320,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1888,624,2000,2000,2000,2000,1952,752,-1856,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1664,832,1648,2000,1488,0,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-544,336,-1680,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,}; 
logic [BITS - 1 : 0] arr_9_digit_9 [0 : WIDTH-1]= '{-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1456,-1136,144,1168,1136,-512,-1440,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1312,384,1696,2016,2016,2016,2016,2016,1952,1328,368,-1936,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1296,400,1792,2016,2016,1584,608,80,1968,1152,2016,1616,1552,-368,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,400,1696,2016,2016,944,224,-1904,-2048,-2048,1008,-1392,1120,1888,1520,2000,-1696,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1904,-16,2000,2016,1680,0,-1856,-2048,-2048,-2048,-2048,1312,-1344,-912,2016,2016,2016,-1696,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-880,1840,2016,1600,-1168,-2048,-2048,-2048,-2048,-1984,-1520,-176,1552,1824,2016,2048,544,-1952,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-832,1792,2016,1520,-288,160,800,800,656,1312,1968,1648,2016,2016,2016,1664,-1424,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1888,752,1856,2000,2048,2016,2016,1968,2016,2016,2016,2016,2016,1984,688,-1632,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1776,128,1072,768,288,400,1152,2016,2016,2016,2016,352,-1776,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,544,2016,2016,1808,-448,-1984,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-144,1952,2016,2016,-592,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-432,1824,2016,2016,1328,-1920,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1168,1808,2016,2016,1824,-1088,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,48,2016,2016,1856,-1008,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1824,1936,2016,2016,384,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-1840,1600,2016,2016,1280,-1904,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-784,2048,2016,2016,-976,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1296,2016,2016,144,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,1584,2048,1680,-1632,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-224,2048,-304,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,}; 
