`timescale 1ns / 1ps 
 
////////////////////////////////////////////////////////////////////////////////// 
// WEIGHT MEMORY (ROM) 
////////////////////////////////////////////////////////////////////////////////// 
module ROM_weights_3 #( 
    parameter int WGHT_INT = 6, // integer part 
    parameter int WGHT_FRC = 16 // fractional part 
)( 
    input logic clk, // clock 
    input logic [9:0] address,
    output [WGHT_INT + WGHT_FRC-1:0] dout 
); 

(* rom_style = "block" *) reg [WGHT_INT + WGHT_FRC-1:0] data;
generate 
  if (WGHT_FRC == 1) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 7'h00; 
        10'b0000000001: data <= 7'h00; 
        10'b0000000010: data <= 7'h00; 
        10'b0000000011: data <= 7'h00; 
        10'b0000000100: data <= 7'h00; 
        10'b0000000101: data <= 7'h00; 
        10'b0000000110: data <= 7'h00; 
        10'b0000000111: data <= 7'h00; 
        10'b0000001000: data <= 7'h00; 
        10'b0000001001: data <= 7'h00; 
        10'b0000001010: data <= 7'h00; 
        10'b0000001011: data <= 7'h00; 
        10'b0000001100: data <= 7'h00; 
        10'b0000001101: data <= 7'h00; 
        10'b0000001110: data <= 7'h00; 
        10'b0000001111: data <= 7'h00; 
        10'b0000010000: data <= 7'h00; 
        10'b0000010001: data <= 7'h00; 
        10'b0000010010: data <= 7'h00; 
        10'b0000010011: data <= 7'h00; 
        10'b0000010100: data <= 7'h00; 
        10'b0000010101: data <= 7'h00; 
        10'b0000010110: data <= 7'h00; 
        10'b0000010111: data <= 7'h00; 
        10'b0000011000: data <= 7'h00; 
        10'b0000011001: data <= 7'h00; 
        10'b0000011010: data <= 7'h00; 
        10'b0000011011: data <= 7'h00; 
        10'b0000011100: data <= 7'h00; 
        10'b0000011101: data <= 7'h00; 
        10'b0000011110: data <= 7'h00; 
        10'b0000011111: data <= 7'h00; 
        10'b0000100000: data <= 7'h00; 
        10'b0000100001: data <= 7'h00; 
        10'b0000100010: data <= 7'h00; 
        10'b0000100011: data <= 7'h00; 
        10'b0000100100: data <= 7'h00; 
        10'b0000100101: data <= 7'h00; 
        10'b0000100110: data <= 7'h00; 
        10'b0000100111: data <= 7'h00; 
        10'b0000101000: data <= 7'h00; 
        10'b0000101001: data <= 7'h00; 
        10'b0000101010: data <= 7'h00; 
        10'b0000101011: data <= 7'h00; 
        10'b0000101100: data <= 7'h00; 
        10'b0000101101: data <= 7'h00; 
        10'b0000101110: data <= 7'h00; 
        10'b0000101111: data <= 7'h00; 
        10'b0000110000: data <= 7'h00; 
        10'b0000110001: data <= 7'h00; 
        10'b0000110010: data <= 7'h00; 
        10'b0000110011: data <= 7'h00; 
        10'b0000110100: data <= 7'h00; 
        10'b0000110101: data <= 7'h00; 
        10'b0000110110: data <= 7'h00; 
        10'b0000110111: data <= 7'h00; 
        10'b0000111000: data <= 7'h00; 
        10'b0000111001: data <= 7'h00; 
        10'b0000111010: data <= 7'h00; 
        10'b0000111011: data <= 7'h00; 
        10'b0000111100: data <= 7'h00; 
        10'b0000111101: data <= 7'h00; 
        10'b0000111110: data <= 7'h00; 
        10'b0000111111: data <= 7'h00; 
        10'b0001000000: data <= 7'h00; 
        10'b0001000001: data <= 7'h00; 
        10'b0001000010: data <= 7'h00; 
        10'b0001000011: data <= 7'h00; 
        10'b0001000100: data <= 7'h00; 
        10'b0001000101: data <= 7'h00; 
        10'b0001000110: data <= 7'h00; 
        10'b0001000111: data <= 7'h00; 
        10'b0001001000: data <= 7'h00; 
        10'b0001001001: data <= 7'h00; 
        10'b0001001010: data <= 7'h00; 
        10'b0001001011: data <= 7'h00; 
        10'b0001001100: data <= 7'h00; 
        10'b0001001101: data <= 7'h00; 
        10'b0001001110: data <= 7'h00; 
        10'b0001001111: data <= 7'h00; 
        10'b0001010000: data <= 7'h00; 
        10'b0001010001: data <= 7'h00; 
        10'b0001010010: data <= 7'h00; 
        10'b0001010011: data <= 7'h00; 
        10'b0001010100: data <= 7'h00; 
        10'b0001010101: data <= 7'h00; 
        10'b0001010110: data <= 7'h00; 
        10'b0001010111: data <= 7'h00; 
        10'b0001011000: data <= 7'h00; 
        10'b0001011001: data <= 7'h00; 
        10'b0001011010: data <= 7'h00; 
        10'b0001011011: data <= 7'h00; 
        10'b0001011100: data <= 7'h00; 
        10'b0001011101: data <= 7'h00; 
        10'b0001011110: data <= 7'h00; 
        10'b0001011111: data <= 7'h00; 
        10'b0001100000: data <= 7'h00; 
        10'b0001100001: data <= 7'h00; 
        10'b0001100010: data <= 7'h00; 
        10'b0001100011: data <= 7'h00; 
        10'b0001100100: data <= 7'h00; 
        10'b0001100101: data <= 7'h00; 
        10'b0001100110: data <= 7'h00; 
        10'b0001100111: data <= 7'h00; 
        10'b0001101000: data <= 7'h00; 
        10'b0001101001: data <= 7'h00; 
        10'b0001101010: data <= 7'h00; 
        10'b0001101011: data <= 7'h00; 
        10'b0001101100: data <= 7'h00; 
        10'b0001101101: data <= 7'h00; 
        10'b0001101110: data <= 7'h00; 
        10'b0001101111: data <= 7'h00; 
        10'b0001110000: data <= 7'h00; 
        10'b0001110001: data <= 7'h00; 
        10'b0001110010: data <= 7'h00; 
        10'b0001110011: data <= 7'h00; 
        10'b0001110100: data <= 7'h00; 
        10'b0001110101: data <= 7'h00; 
        10'b0001110110: data <= 7'h00; 
        10'b0001110111: data <= 7'h00; 
        10'b0001111000: data <= 7'h00; 
        10'b0001111001: data <= 7'h00; 
        10'b0001111010: data <= 7'h00; 
        10'b0001111011: data <= 7'h01; 
        10'b0001111100: data <= 7'h01; 
        10'b0001111101: data <= 7'h01; 
        10'b0001111110: data <= 7'h01; 
        10'b0001111111: data <= 7'h00; 
        10'b0010000000: data <= 7'h00; 
        10'b0010000001: data <= 7'h00; 
        10'b0010000010: data <= 7'h00; 
        10'b0010000011: data <= 7'h00; 
        10'b0010000100: data <= 7'h00; 
        10'b0010000101: data <= 7'h00; 
        10'b0010000110: data <= 7'h00; 
        10'b0010000111: data <= 7'h00; 
        10'b0010001000: data <= 7'h00; 
        10'b0010001001: data <= 7'h00; 
        10'b0010001010: data <= 7'h00; 
        10'b0010001011: data <= 7'h00; 
        10'b0010001100: data <= 7'h00; 
        10'b0010001101: data <= 7'h00; 
        10'b0010001110: data <= 7'h00; 
        10'b0010001111: data <= 7'h00; 
        10'b0010010000: data <= 7'h00; 
        10'b0010010001: data <= 7'h00; 
        10'b0010010010: data <= 7'h00; 
        10'b0010010011: data <= 7'h00; 
        10'b0010010100: data <= 7'h00; 
        10'b0010010101: data <= 7'h00; 
        10'b0010010110: data <= 7'h00; 
        10'b0010010111: data <= 7'h00; 
        10'b0010011000: data <= 7'h00; 
        10'b0010011001: data <= 7'h00; 
        10'b0010011010: data <= 7'h00; 
        10'b0010011011: data <= 7'h00; 
        10'b0010011100: data <= 7'h00; 
        10'b0010011101: data <= 7'h00; 
        10'b0010011110: data <= 7'h00; 
        10'b0010011111: data <= 7'h00; 
        10'b0010100000: data <= 7'h00; 
        10'b0010100001: data <= 7'h00; 
        10'b0010100010: data <= 7'h7f; 
        10'b0010100011: data <= 7'h00; 
        10'b0010100100: data <= 7'h00; 
        10'b0010100101: data <= 7'h00; 
        10'b0010100110: data <= 7'h00; 
        10'b0010100111: data <= 7'h00; 
        10'b0010101000: data <= 7'h00; 
        10'b0010101001: data <= 7'h00; 
        10'b0010101010: data <= 7'h00; 
        10'b0010101011: data <= 7'h00; 
        10'b0010101100: data <= 7'h00; 
        10'b0010101101: data <= 7'h00; 
        10'b0010101110: data <= 7'h00; 
        10'b0010101111: data <= 7'h00; 
        10'b0010110000: data <= 7'h00; 
        10'b0010110001: data <= 7'h00; 
        10'b0010110010: data <= 7'h00; 
        10'b0010110011: data <= 7'h00; 
        10'b0010110100: data <= 7'h00; 
        10'b0010110101: data <= 7'h01; 
        10'b0010110110: data <= 7'h00; 
        10'b0010110111: data <= 7'h00; 
        10'b0010111000: data <= 7'h00; 
        10'b0010111001: data <= 7'h00; 
        10'b0010111010: data <= 7'h00; 
        10'b0010111011: data <= 7'h00; 
        10'b0010111100: data <= 7'h00; 
        10'b0010111101: data <= 7'h00; 
        10'b0010111110: data <= 7'h00; 
        10'b0010111111: data <= 7'h00; 
        10'b0011000000: data <= 7'h00; 
        10'b0011000001: data <= 7'h00; 
        10'b0011000010: data <= 7'h00; 
        10'b0011000011: data <= 7'h00; 
        10'b0011000100: data <= 7'h00; 
        10'b0011000101: data <= 7'h00; 
        10'b0011000110: data <= 7'h00; 
        10'b0011000111: data <= 7'h00; 
        10'b0011001000: data <= 7'h01; 
        10'b0011001001: data <= 7'h01; 
        10'b0011001010: data <= 7'h00; 
        10'b0011001011: data <= 7'h00; 
        10'b0011001100: data <= 7'h00; 
        10'b0011001101: data <= 7'h00; 
        10'b0011001110: data <= 7'h00; 
        10'b0011001111: data <= 7'h00; 
        10'b0011010000: data <= 7'h00; 
        10'b0011010001: data <= 7'h00; 
        10'b0011010010: data <= 7'h00; 
        10'b0011010011: data <= 7'h00; 
        10'b0011010100: data <= 7'h00; 
        10'b0011010101: data <= 7'h00; 
        10'b0011010110: data <= 7'h00; 
        10'b0011010111: data <= 7'h00; 
        10'b0011011000: data <= 7'h00; 
        10'b0011011001: data <= 7'h00; 
        10'b0011011010: data <= 7'h00; 
        10'b0011011011: data <= 7'h7f; 
        10'b0011011100: data <= 7'h00; 
        10'b0011011101: data <= 7'h00; 
        10'b0011011110: data <= 7'h00; 
        10'b0011011111: data <= 7'h00; 
        10'b0011100000: data <= 7'h00; 
        10'b0011100001: data <= 7'h00; 
        10'b0011100010: data <= 7'h00; 
        10'b0011100011: data <= 7'h00; 
        10'b0011100100: data <= 7'h00; 
        10'b0011100101: data <= 7'h00; 
        10'b0011100110: data <= 7'h00; 
        10'b0011100111: data <= 7'h00; 
        10'b0011101000: data <= 7'h00; 
        10'b0011101001: data <= 7'h00; 
        10'b0011101010: data <= 7'h00; 
        10'b0011101011: data <= 7'h00; 
        10'b0011101100: data <= 7'h00; 
        10'b0011101101: data <= 7'h00; 
        10'b0011101110: data <= 7'h01; 
        10'b0011101111: data <= 7'h00; 
        10'b0011110000: data <= 7'h00; 
        10'b0011110001: data <= 7'h00; 
        10'b0011110010: data <= 7'h00; 
        10'b0011110011: data <= 7'h00; 
        10'b0011110100: data <= 7'h00; 
        10'b0011110101: data <= 7'h00; 
        10'b0011110110: data <= 7'h00; 
        10'b0011110111: data <= 7'h00; 
        10'b0011111000: data <= 7'h00; 
        10'b0011111001: data <= 7'h00; 
        10'b0011111010: data <= 7'h00; 
        10'b0011111011: data <= 7'h00; 
        10'b0011111100: data <= 7'h00; 
        10'b0011111101: data <= 7'h00; 
        10'b0011111110: data <= 7'h00; 
        10'b0011111111: data <= 7'h00; 
        10'b0100000000: data <= 7'h00; 
        10'b0100000001: data <= 7'h00; 
        10'b0100000010: data <= 7'h00; 
        10'b0100000011: data <= 7'h00; 
        10'b0100000100: data <= 7'h00; 
        10'b0100000101: data <= 7'h00; 
        10'b0100000110: data <= 7'h00; 
        10'b0100000111: data <= 7'h7f; 
        10'b0100001000: data <= 7'h7f; 
        10'b0100001001: data <= 7'h00; 
        10'b0100001010: data <= 7'h01; 
        10'b0100001011: data <= 7'h01; 
        10'b0100001100: data <= 7'h01; 
        10'b0100001101: data <= 7'h00; 
        10'b0100001110: data <= 7'h00; 
        10'b0100001111: data <= 7'h00; 
        10'b0100010000: data <= 7'h00; 
        10'b0100010001: data <= 7'h00; 
        10'b0100010010: data <= 7'h00; 
        10'b0100010011: data <= 7'h00; 
        10'b0100010100: data <= 7'h00; 
        10'b0100010101: data <= 7'h00; 
        10'b0100010110: data <= 7'h00; 
        10'b0100010111: data <= 7'h00; 
        10'b0100011000: data <= 7'h00; 
        10'b0100011001: data <= 7'h00; 
        10'b0100011010: data <= 7'h00; 
        10'b0100011011: data <= 7'h00; 
        10'b0100011100: data <= 7'h00; 
        10'b0100011101: data <= 7'h00; 
        10'b0100011110: data <= 7'h00; 
        10'b0100011111: data <= 7'h00; 
        10'b0100100000: data <= 7'h7f; 
        10'b0100100001: data <= 7'h7f; 
        10'b0100100010: data <= 7'h7f; 
        10'b0100100011: data <= 7'h7f; 
        10'b0100100100: data <= 7'h7f; 
        10'b0100100101: data <= 7'h00; 
        10'b0100100110: data <= 7'h00; 
        10'b0100100111: data <= 7'h01; 
        10'b0100101000: data <= 7'h00; 
        10'b0100101001: data <= 7'h00; 
        10'b0100101010: data <= 7'h00; 
        10'b0100101011: data <= 7'h00; 
        10'b0100101100: data <= 7'h00; 
        10'b0100101101: data <= 7'h00; 
        10'b0100101110: data <= 7'h00; 
        10'b0100101111: data <= 7'h00; 
        10'b0100110000: data <= 7'h00; 
        10'b0100110001: data <= 7'h00; 
        10'b0100110010: data <= 7'h00; 
        10'b0100110011: data <= 7'h00; 
        10'b0100110100: data <= 7'h00; 
        10'b0100110101: data <= 7'h00; 
        10'b0100110110: data <= 7'h00; 
        10'b0100110111: data <= 7'h00; 
        10'b0100111000: data <= 7'h00; 
        10'b0100111001: data <= 7'h00; 
        10'b0100111010: data <= 7'h7f; 
        10'b0100111011: data <= 7'h7f; 
        10'b0100111100: data <= 7'h7f; 
        10'b0100111101: data <= 7'h7f; 
        10'b0100111110: data <= 7'h7f; 
        10'b0100111111: data <= 7'h00; 
        10'b0101000000: data <= 7'h00; 
        10'b0101000001: data <= 7'h00; 
        10'b0101000010: data <= 7'h00; 
        10'b0101000011: data <= 7'h00; 
        10'b0101000100: data <= 7'h00; 
        10'b0101000101: data <= 7'h00; 
        10'b0101000110: data <= 7'h00; 
        10'b0101000111: data <= 7'h00; 
        10'b0101001000: data <= 7'h00; 
        10'b0101001001: data <= 7'h00; 
        10'b0101001010: data <= 7'h00; 
        10'b0101001011: data <= 7'h00; 
        10'b0101001100: data <= 7'h00; 
        10'b0101001101: data <= 7'h00; 
        10'b0101001110: data <= 7'h00; 
        10'b0101001111: data <= 7'h00; 
        10'b0101010000: data <= 7'h00; 
        10'b0101010001: data <= 7'h00; 
        10'b0101010010: data <= 7'h00; 
        10'b0101010011: data <= 7'h00; 
        10'b0101010100: data <= 7'h00; 
        10'b0101010101: data <= 7'h00; 
        10'b0101010110: data <= 7'h7f; 
        10'b0101010111: data <= 7'h7f; 
        10'b0101011000: data <= 7'h7f; 
        10'b0101011001: data <= 7'h00; 
        10'b0101011010: data <= 7'h00; 
        10'b0101011011: data <= 7'h00; 
        10'b0101011100: data <= 7'h00; 
        10'b0101011101: data <= 7'h00; 
        10'b0101011110: data <= 7'h01; 
        10'b0101011111: data <= 7'h00; 
        10'b0101100000: data <= 7'h00; 
        10'b0101100001: data <= 7'h00; 
        10'b0101100010: data <= 7'h00; 
        10'b0101100011: data <= 7'h00; 
        10'b0101100100: data <= 7'h00; 
        10'b0101100101: data <= 7'h00; 
        10'b0101100110: data <= 7'h00; 
        10'b0101100111: data <= 7'h00; 
        10'b0101101000: data <= 7'h00; 
        10'b0101101001: data <= 7'h00; 
        10'b0101101010: data <= 7'h00; 
        10'b0101101011: data <= 7'h00; 
        10'b0101101100: data <= 7'h00; 
        10'b0101101101: data <= 7'h00; 
        10'b0101101110: data <= 7'h00; 
        10'b0101101111: data <= 7'h00; 
        10'b0101110000: data <= 7'h00; 
        10'b0101110001: data <= 7'h00; 
        10'b0101110010: data <= 7'h7f; 
        10'b0101110011: data <= 7'h7f; 
        10'b0101110100: data <= 7'h00; 
        10'b0101110101: data <= 7'h00; 
        10'b0101110110: data <= 7'h00; 
        10'b0101110111: data <= 7'h00; 
        10'b0101111000: data <= 7'h00; 
        10'b0101111001: data <= 7'h00; 
        10'b0101111010: data <= 7'h00; 
        10'b0101111011: data <= 7'h00; 
        10'b0101111100: data <= 7'h00; 
        10'b0101111101: data <= 7'h00; 
        10'b0101111110: data <= 7'h00; 
        10'b0101111111: data <= 7'h00; 
        10'b0110000000: data <= 7'h00; 
        10'b0110000001: data <= 7'h00; 
        10'b0110000010: data <= 7'h00; 
        10'b0110000011: data <= 7'h00; 
        10'b0110000100: data <= 7'h00; 
        10'b0110000101: data <= 7'h00; 
        10'b0110000110: data <= 7'h00; 
        10'b0110000111: data <= 7'h00; 
        10'b0110001000: data <= 7'h00; 
        10'b0110001001: data <= 7'h00; 
        10'b0110001010: data <= 7'h00; 
        10'b0110001011: data <= 7'h00; 
        10'b0110001100: data <= 7'h00; 
        10'b0110001101: data <= 7'h00; 
        10'b0110001110: data <= 7'h00; 
        10'b0110001111: data <= 7'h00; 
        10'b0110010000: data <= 7'h00; 
        10'b0110010001: data <= 7'h00; 
        10'b0110010010: data <= 7'h00; 
        10'b0110010011: data <= 7'h00; 
        10'b0110010100: data <= 7'h00; 
        10'b0110010101: data <= 7'h00; 
        10'b0110010110: data <= 7'h00; 
        10'b0110010111: data <= 7'h00; 
        10'b0110011000: data <= 7'h00; 
        10'b0110011001: data <= 7'h00; 
        10'b0110011010: data <= 7'h00; 
        10'b0110011011: data <= 7'h00; 
        10'b0110011100: data <= 7'h00; 
        10'b0110011101: data <= 7'h00; 
        10'b0110011110: data <= 7'h00; 
        10'b0110011111: data <= 7'h00; 
        10'b0110100000: data <= 7'h00; 
        10'b0110100001: data <= 7'h00; 
        10'b0110100010: data <= 7'h00; 
        10'b0110100011: data <= 7'h00; 
        10'b0110100100: data <= 7'h00; 
        10'b0110100101: data <= 7'h00; 
        10'b0110100110: data <= 7'h00; 
        10'b0110100111: data <= 7'h00; 
        10'b0110101000: data <= 7'h00; 
        10'b0110101001: data <= 7'h00; 
        10'b0110101010: data <= 7'h00; 
        10'b0110101011: data <= 7'h00; 
        10'b0110101100: data <= 7'h00; 
        10'b0110101101: data <= 7'h00; 
        10'b0110101110: data <= 7'h00; 
        10'b0110101111: data <= 7'h00; 
        10'b0110110000: data <= 7'h00; 
        10'b0110110001: data <= 7'h00; 
        10'b0110110010: data <= 7'h00; 
        10'b0110110011: data <= 7'h00; 
        10'b0110110100: data <= 7'h00; 
        10'b0110110101: data <= 7'h00; 
        10'b0110110110: data <= 7'h00; 
        10'b0110110111: data <= 7'h00; 
        10'b0110111000: data <= 7'h00; 
        10'b0110111001: data <= 7'h00; 
        10'b0110111010: data <= 7'h00; 
        10'b0110111011: data <= 7'h00; 
        10'b0110111100: data <= 7'h00; 
        10'b0110111101: data <= 7'h00; 
        10'b0110111110: data <= 7'h00; 
        10'b0110111111: data <= 7'h00; 
        10'b0111000000: data <= 7'h00; 
        10'b0111000001: data <= 7'h00; 
        10'b0111000010: data <= 7'h00; 
        10'b0111000011: data <= 7'h00; 
        10'b0111000100: data <= 7'h00; 
        10'b0111000101: data <= 7'h00; 
        10'b0111000110: data <= 7'h00; 
        10'b0111000111: data <= 7'h00; 
        10'b0111001000: data <= 7'h7f; 
        10'b0111001001: data <= 7'h7f; 
        10'b0111001010: data <= 7'h7f; 
        10'b0111001011: data <= 7'h00; 
        10'b0111001100: data <= 7'h00; 
        10'b0111001101: data <= 7'h00; 
        10'b0111001110: data <= 7'h00; 
        10'b0111001111: data <= 7'h00; 
        10'b0111010000: data <= 7'h00; 
        10'b0111010001: data <= 7'h00; 
        10'b0111010010: data <= 7'h00; 
        10'b0111010011: data <= 7'h00; 
        10'b0111010100: data <= 7'h00; 
        10'b0111010101: data <= 7'h00; 
        10'b0111010110: data <= 7'h00; 
        10'b0111010111: data <= 7'h00; 
        10'b0111011000: data <= 7'h00; 
        10'b0111011001: data <= 7'h00; 
        10'b0111011010: data <= 7'h00; 
        10'b0111011011: data <= 7'h00; 
        10'b0111011100: data <= 7'h00; 
        10'b0111011101: data <= 7'h00; 
        10'b0111011110: data <= 7'h00; 
        10'b0111011111: data <= 7'h00; 
        10'b0111100000: data <= 7'h00; 
        10'b0111100001: data <= 7'h00; 
        10'b0111100010: data <= 7'h00; 
        10'b0111100011: data <= 7'h00; 
        10'b0111100100: data <= 7'h7f; 
        10'b0111100101: data <= 7'h7f; 
        10'b0111100110: data <= 7'h7f; 
        10'b0111100111: data <= 7'h7f; 
        10'b0111101000: data <= 7'h7f; 
        10'b0111101001: data <= 7'h7f; 
        10'b0111101010: data <= 7'h7f; 
        10'b0111101011: data <= 7'h00; 
        10'b0111101100: data <= 7'h00; 
        10'b0111101101: data <= 7'h00; 
        10'b0111101110: data <= 7'h00; 
        10'b0111101111: data <= 7'h00; 
        10'b0111110000: data <= 7'h00; 
        10'b0111110001: data <= 7'h00; 
        10'b0111110010: data <= 7'h00; 
        10'b0111110011: data <= 7'h00; 
        10'b0111110100: data <= 7'h00; 
        10'b0111110101: data <= 7'h00; 
        10'b0111110110: data <= 7'h00; 
        10'b0111110111: data <= 7'h00; 
        10'b0111111000: data <= 7'h00; 
        10'b0111111001: data <= 7'h00; 
        10'b0111111010: data <= 7'h00; 
        10'b0111111011: data <= 7'h00; 
        10'b0111111100: data <= 7'h00; 
        10'b0111111101: data <= 7'h00; 
        10'b0111111110: data <= 7'h00; 
        10'b0111111111: data <= 7'h00; 
        10'b1000000000: data <= 7'h00; 
        10'b1000000001: data <= 7'h7f; 
        10'b1000000010: data <= 7'h7f; 
        10'b1000000011: data <= 7'h7f; 
        10'b1000000100: data <= 7'h7f; 
        10'b1000000101: data <= 7'h7f; 
        10'b1000000110: data <= 7'h7f; 
        10'b1000000111: data <= 7'h00; 
        10'b1000001000: data <= 7'h00; 
        10'b1000001001: data <= 7'h00; 
        10'b1000001010: data <= 7'h00; 
        10'b1000001011: data <= 7'h00; 
        10'b1000001100: data <= 7'h00; 
        10'b1000001101: data <= 7'h01; 
        10'b1000001110: data <= 7'h01; 
        10'b1000001111: data <= 7'h00; 
        10'b1000010000: data <= 7'h00; 
        10'b1000010001: data <= 7'h00; 
        10'b1000010010: data <= 7'h00; 
        10'b1000010011: data <= 7'h00; 
        10'b1000010100: data <= 7'h00; 
        10'b1000010101: data <= 7'h00; 
        10'b1000010110: data <= 7'h00; 
        10'b1000010111: data <= 7'h00; 
        10'b1000011000: data <= 7'h00; 
        10'b1000011001: data <= 7'h00; 
        10'b1000011010: data <= 7'h00; 
        10'b1000011011: data <= 7'h00; 
        10'b1000011100: data <= 7'h00; 
        10'b1000011101: data <= 7'h00; 
        10'b1000011110: data <= 7'h00; 
        10'b1000011111: data <= 7'h00; 
        10'b1000100000: data <= 7'h7f; 
        10'b1000100001: data <= 7'h7f; 
        10'b1000100010: data <= 7'h00; 
        10'b1000100011: data <= 7'h00; 
        10'b1000100100: data <= 7'h00; 
        10'b1000100101: data <= 7'h00; 
        10'b1000100110: data <= 7'h01; 
        10'b1000100111: data <= 7'h00; 
        10'b1000101000: data <= 7'h00; 
        10'b1000101001: data <= 7'h00; 
        10'b1000101010: data <= 7'h00; 
        10'b1000101011: data <= 7'h00; 
        10'b1000101100: data <= 7'h00; 
        10'b1000101101: data <= 7'h00; 
        10'b1000101110: data <= 7'h00; 
        10'b1000101111: data <= 7'h00; 
        10'b1000110000: data <= 7'h00; 
        10'b1000110001: data <= 7'h00; 
        10'b1000110010: data <= 7'h00; 
        10'b1000110011: data <= 7'h00; 
        10'b1000110100: data <= 7'h01; 
        10'b1000110101: data <= 7'h01; 
        10'b1000110110: data <= 7'h01; 
        10'b1000110111: data <= 7'h00; 
        10'b1000111000: data <= 7'h00; 
        10'b1000111001: data <= 7'h00; 
        10'b1000111010: data <= 7'h00; 
        10'b1000111011: data <= 7'h00; 
        10'b1000111100: data <= 7'h00; 
        10'b1000111101: data <= 7'h00; 
        10'b1000111110: data <= 7'h00; 
        10'b1000111111: data <= 7'h00; 
        10'b1001000000: data <= 7'h00; 
        10'b1001000001: data <= 7'h00; 
        10'b1001000010: data <= 7'h00; 
        10'b1001000011: data <= 7'h00; 
        10'b1001000100: data <= 7'h00; 
        10'b1001000101: data <= 7'h00; 
        10'b1001000110: data <= 7'h00; 
        10'b1001000111: data <= 7'h00; 
        10'b1001001000: data <= 7'h00; 
        10'b1001001001: data <= 7'h00; 
        10'b1001001010: data <= 7'h00; 
        10'b1001001011: data <= 7'h00; 
        10'b1001001100: data <= 7'h00; 
        10'b1001001101: data <= 7'h00; 
        10'b1001001110: data <= 7'h00; 
        10'b1001001111: data <= 7'h00; 
        10'b1001010000: data <= 7'h01; 
        10'b1001010001: data <= 7'h01; 
        10'b1001010010: data <= 7'h00; 
        10'b1001010011: data <= 7'h00; 
        10'b1001010100: data <= 7'h00; 
        10'b1001010101: data <= 7'h00; 
        10'b1001010110: data <= 7'h00; 
        10'b1001010111: data <= 7'h00; 
        10'b1001011000: data <= 7'h00; 
        10'b1001011001: data <= 7'h00; 
        10'b1001011010: data <= 7'h00; 
        10'b1001011011: data <= 7'h00; 
        10'b1001011100: data <= 7'h00; 
        10'b1001011101: data <= 7'h00; 
        10'b1001011110: data <= 7'h00; 
        10'b1001011111: data <= 7'h00; 
        10'b1001100000: data <= 7'h00; 
        10'b1001100001: data <= 7'h00; 
        10'b1001100010: data <= 7'h00; 
        10'b1001100011: data <= 7'h00; 
        10'b1001100100: data <= 7'h00; 
        10'b1001100101: data <= 7'h00; 
        10'b1001100110: data <= 7'h00; 
        10'b1001100111: data <= 7'h00; 
        10'b1001101000: data <= 7'h00; 
        10'b1001101001: data <= 7'h00; 
        10'b1001101010: data <= 7'h00; 
        10'b1001101011: data <= 7'h00; 
        10'b1001101100: data <= 7'h00; 
        10'b1001101101: data <= 7'h00; 
        10'b1001101110: data <= 7'h00; 
        10'b1001101111: data <= 7'h00; 
        10'b1001110000: data <= 7'h00; 
        10'b1001110001: data <= 7'h00; 
        10'b1001110010: data <= 7'h00; 
        10'b1001110011: data <= 7'h00; 
        10'b1001110100: data <= 7'h00; 
        10'b1001110101: data <= 7'h00; 
        10'b1001110110: data <= 7'h00; 
        10'b1001110111: data <= 7'h00; 
        10'b1001111000: data <= 7'h00; 
        10'b1001111001: data <= 7'h00; 
        10'b1001111010: data <= 7'h00; 
        10'b1001111011: data <= 7'h00; 
        10'b1001111100: data <= 7'h00; 
        10'b1001111101: data <= 7'h00; 
        10'b1001111110: data <= 7'h00; 
        10'b1001111111: data <= 7'h00; 
        10'b1010000000: data <= 7'h00; 
        10'b1010000001: data <= 7'h00; 
        10'b1010000010: data <= 7'h00; 
        10'b1010000011: data <= 7'h00; 
        10'b1010000100: data <= 7'h00; 
        10'b1010000101: data <= 7'h00; 
        10'b1010000110: data <= 7'h00; 
        10'b1010000111: data <= 7'h00; 
        10'b1010001000: data <= 7'h00; 
        10'b1010001001: data <= 7'h00; 
        10'b1010001010: data <= 7'h00; 
        10'b1010001011: data <= 7'h00; 
        10'b1010001100: data <= 7'h00; 
        10'b1010001101: data <= 7'h00; 
        10'b1010001110: data <= 7'h00; 
        10'b1010001111: data <= 7'h00; 
        10'b1010010000: data <= 7'h00; 
        10'b1010010001: data <= 7'h00; 
        10'b1010010010: data <= 7'h00; 
        10'b1010010011: data <= 7'h00; 
        10'b1010010100: data <= 7'h00; 
        10'b1010010101: data <= 7'h00; 
        10'b1010010110: data <= 7'h00; 
        10'b1010010111: data <= 7'h00; 
        10'b1010011000: data <= 7'h00; 
        10'b1010011001: data <= 7'h00; 
        10'b1010011010: data <= 7'h00; 
        10'b1010011011: data <= 7'h00; 
        10'b1010011100: data <= 7'h00; 
        10'b1010011101: data <= 7'h00; 
        10'b1010011110: data <= 7'h00; 
        10'b1010011111: data <= 7'h00; 
        10'b1010100000: data <= 7'h00; 
        10'b1010100001: data <= 7'h00; 
        10'b1010100010: data <= 7'h00; 
        10'b1010100011: data <= 7'h00; 
        10'b1010100100: data <= 7'h00; 
        10'b1010100101: data <= 7'h00; 
        10'b1010100110: data <= 7'h00; 
        10'b1010100111: data <= 7'h00; 
        10'b1010101000: data <= 7'h00; 
        10'b1010101001: data <= 7'h00; 
        10'b1010101010: data <= 7'h00; 
        10'b1010101011: data <= 7'h01; 
        10'b1010101100: data <= 7'h01; 
        10'b1010101101: data <= 7'h00; 
        10'b1010101110: data <= 7'h00; 
        10'b1010101111: data <= 7'h00; 
        10'b1010110000: data <= 7'h00; 
        10'b1010110001: data <= 7'h00; 
        10'b1010110010: data <= 7'h00; 
        10'b1010110011: data <= 7'h00; 
        10'b1010110100: data <= 7'h00; 
        10'b1010110101: data <= 7'h00; 
        10'b1010110110: data <= 7'h00; 
        10'b1010110111: data <= 7'h00; 
        10'b1010111000: data <= 7'h00; 
        10'b1010111001: data <= 7'h00; 
        10'b1010111010: data <= 7'h00; 
        10'b1010111011: data <= 7'h00; 
        10'b1010111100: data <= 7'h00; 
        10'b1010111101: data <= 7'h00; 
        10'b1010111110: data <= 7'h00; 
        10'b1010111111: data <= 7'h00; 
        10'b1011000000: data <= 7'h00; 
        10'b1011000001: data <= 7'h00; 
        10'b1011000010: data <= 7'h00; 
        10'b1011000011: data <= 7'h00; 
        10'b1011000100: data <= 7'h00; 
        10'b1011000101: data <= 7'h00; 
        10'b1011000110: data <= 7'h00; 
        10'b1011000111: data <= 7'h00; 
        10'b1011001000: data <= 7'h01; 
        10'b1011001001: data <= 7'h00; 
        10'b1011001010: data <= 7'h00; 
        10'b1011001011: data <= 7'h00; 
        10'b1011001100: data <= 7'h00; 
        10'b1011001101: data <= 7'h00; 
        10'b1011001110: data <= 7'h00; 
        10'b1011001111: data <= 7'h00; 
        10'b1011010000: data <= 7'h00; 
        10'b1011010001: data <= 7'h00; 
        10'b1011010010: data <= 7'h00; 
        10'b1011010011: data <= 7'h00; 
        10'b1011010100: data <= 7'h00; 
        10'b1011010101: data <= 7'h00; 
        10'b1011010110: data <= 7'h00; 
        10'b1011010111: data <= 7'h00; 
        10'b1011011000: data <= 7'h00; 
        10'b1011011001: data <= 7'h00; 
        10'b1011011010: data <= 7'h00; 
        10'b1011011011: data <= 7'h00; 
        10'b1011011100: data <= 7'h00; 
        10'b1011011101: data <= 7'h00; 
        10'b1011011110: data <= 7'h00; 
        10'b1011011111: data <= 7'h00; 
        10'b1011100000: data <= 7'h00; 
        10'b1011100001: data <= 7'h00; 
        10'b1011100010: data <= 7'h00; 
        10'b1011100011: data <= 7'h00; 
        10'b1011100100: data <= 7'h00; 
        10'b1011100101: data <= 7'h00; 
        10'b1011100110: data <= 7'h00; 
        10'b1011100111: data <= 7'h00; 
        10'b1011101000: data <= 7'h00; 
        10'b1011101001: data <= 7'h00; 
        10'b1011101010: data <= 7'h00; 
        10'b1011101011: data <= 7'h00; 
        10'b1011101100: data <= 7'h00; 
        10'b1011101101: data <= 7'h00; 
        10'b1011101110: data <= 7'h00; 
        10'b1011101111: data <= 7'h00; 
        10'b1011110000: data <= 7'h00; 
        10'b1011110001: data <= 7'h00; 
        10'b1011110010: data <= 7'h00; 
        10'b1011110011: data <= 7'h00; 
        10'b1011110100: data <= 7'h00; 
        10'b1011110101: data <= 7'h00; 
        10'b1011110110: data <= 7'h00; 
        10'b1011110111: data <= 7'h00; 
        10'b1011111000: data <= 7'h00; 
        10'b1011111001: data <= 7'h00; 
        10'b1011111010: data <= 7'h00; 
        10'b1011111011: data <= 7'h00; 
        10'b1011111100: data <= 7'h00; 
        10'b1011111101: data <= 7'h00; 
        10'b1011111110: data <= 7'h00; 
        10'b1011111111: data <= 7'h00; 
        10'b1100000000: data <= 7'h00; 
        10'b1100000001: data <= 7'h00; 
        10'b1100000010: data <= 7'h00; 
        10'b1100000011: data <= 7'h00; 
        10'b1100000100: data <= 7'h00; 
        10'b1100000101: data <= 7'h00; 
        10'b1100000110: data <= 7'h00; 
        10'b1100000111: data <= 7'h00; 
        10'b1100001000: data <= 7'h00; 
        10'b1100001001: data <= 7'h00; 
        10'b1100001010: data <= 7'h00; 
        10'b1100001011: data <= 7'h00; 
        10'b1100001100: data <= 7'h00; 
        10'b1100001101: data <= 7'h00; 
        10'b1100001110: data <= 7'h00; 
        10'b1100001111: data <= 7'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 2) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 8'h00; 
        10'b0000000001: data <= 8'h00; 
        10'b0000000010: data <= 8'h00; 
        10'b0000000011: data <= 8'h00; 
        10'b0000000100: data <= 8'h00; 
        10'b0000000101: data <= 8'h00; 
        10'b0000000110: data <= 8'h00; 
        10'b0000000111: data <= 8'h00; 
        10'b0000001000: data <= 8'h00; 
        10'b0000001001: data <= 8'h00; 
        10'b0000001010: data <= 8'h00; 
        10'b0000001011: data <= 8'h00; 
        10'b0000001100: data <= 8'h00; 
        10'b0000001101: data <= 8'h00; 
        10'b0000001110: data <= 8'h00; 
        10'b0000001111: data <= 8'h00; 
        10'b0000010000: data <= 8'h00; 
        10'b0000010001: data <= 8'h00; 
        10'b0000010010: data <= 8'h00; 
        10'b0000010011: data <= 8'h00; 
        10'b0000010100: data <= 8'h00; 
        10'b0000010101: data <= 8'h00; 
        10'b0000010110: data <= 8'h00; 
        10'b0000010111: data <= 8'h00; 
        10'b0000011000: data <= 8'h00; 
        10'b0000011001: data <= 8'h00; 
        10'b0000011010: data <= 8'h00; 
        10'b0000011011: data <= 8'h00; 
        10'b0000011100: data <= 8'h00; 
        10'b0000011101: data <= 8'h00; 
        10'b0000011110: data <= 8'h00; 
        10'b0000011111: data <= 8'h00; 
        10'b0000100000: data <= 8'h00; 
        10'b0000100001: data <= 8'h00; 
        10'b0000100010: data <= 8'h00; 
        10'b0000100011: data <= 8'h00; 
        10'b0000100100: data <= 8'h00; 
        10'b0000100101: data <= 8'h00; 
        10'b0000100110: data <= 8'h00; 
        10'b0000100111: data <= 8'h00; 
        10'b0000101000: data <= 8'h00; 
        10'b0000101001: data <= 8'h00; 
        10'b0000101010: data <= 8'h00; 
        10'b0000101011: data <= 8'h00; 
        10'b0000101100: data <= 8'h00; 
        10'b0000101101: data <= 8'h00; 
        10'b0000101110: data <= 8'h00; 
        10'b0000101111: data <= 8'h00; 
        10'b0000110000: data <= 8'h00; 
        10'b0000110001: data <= 8'h00; 
        10'b0000110010: data <= 8'h00; 
        10'b0000110011: data <= 8'h00; 
        10'b0000110100: data <= 8'h00; 
        10'b0000110101: data <= 8'h00; 
        10'b0000110110: data <= 8'h00; 
        10'b0000110111: data <= 8'h00; 
        10'b0000111000: data <= 8'h00; 
        10'b0000111001: data <= 8'h00; 
        10'b0000111010: data <= 8'h00; 
        10'b0000111011: data <= 8'h00; 
        10'b0000111100: data <= 8'h00; 
        10'b0000111101: data <= 8'h00; 
        10'b0000111110: data <= 8'h00; 
        10'b0000111111: data <= 8'h00; 
        10'b0001000000: data <= 8'h00; 
        10'b0001000001: data <= 8'h00; 
        10'b0001000010: data <= 8'h00; 
        10'b0001000011: data <= 8'h00; 
        10'b0001000100: data <= 8'h00; 
        10'b0001000101: data <= 8'h00; 
        10'b0001000110: data <= 8'h00; 
        10'b0001000111: data <= 8'h00; 
        10'b0001001000: data <= 8'h00; 
        10'b0001001001: data <= 8'h00; 
        10'b0001001010: data <= 8'h00; 
        10'b0001001011: data <= 8'h00; 
        10'b0001001100: data <= 8'h00; 
        10'b0001001101: data <= 8'h00; 
        10'b0001001110: data <= 8'h00; 
        10'b0001001111: data <= 8'h00; 
        10'b0001010000: data <= 8'h00; 
        10'b0001010001: data <= 8'h00; 
        10'b0001010010: data <= 8'h00; 
        10'b0001010011: data <= 8'h00; 
        10'b0001010100: data <= 8'h00; 
        10'b0001010101: data <= 8'h00; 
        10'b0001010110: data <= 8'h00; 
        10'b0001010111: data <= 8'h00; 
        10'b0001011000: data <= 8'h00; 
        10'b0001011001: data <= 8'h00; 
        10'b0001011010: data <= 8'h00; 
        10'b0001011011: data <= 8'h00; 
        10'b0001011100: data <= 8'h00; 
        10'b0001011101: data <= 8'h00; 
        10'b0001011110: data <= 8'h00; 
        10'b0001011111: data <= 8'h00; 
        10'b0001100000: data <= 8'h01; 
        10'b0001100001: data <= 8'h01; 
        10'b0001100010: data <= 8'h01; 
        10'b0001100011: data <= 8'h01; 
        10'b0001100100: data <= 8'h00; 
        10'b0001100101: data <= 8'h00; 
        10'b0001100110: data <= 8'h00; 
        10'b0001100111: data <= 8'h00; 
        10'b0001101000: data <= 8'h00; 
        10'b0001101001: data <= 8'h00; 
        10'b0001101010: data <= 8'h00; 
        10'b0001101011: data <= 8'h00; 
        10'b0001101100: data <= 8'h00; 
        10'b0001101101: data <= 8'h00; 
        10'b0001101110: data <= 8'h00; 
        10'b0001101111: data <= 8'h00; 
        10'b0001110000: data <= 8'h00; 
        10'b0001110001: data <= 8'h00; 
        10'b0001110010: data <= 8'h00; 
        10'b0001110011: data <= 8'h00; 
        10'b0001110100: data <= 8'h00; 
        10'b0001110101: data <= 8'h00; 
        10'b0001110110: data <= 8'h00; 
        10'b0001110111: data <= 8'h00; 
        10'b0001111000: data <= 8'h01; 
        10'b0001111001: data <= 8'h01; 
        10'b0001111010: data <= 8'h01; 
        10'b0001111011: data <= 8'h01; 
        10'b0001111100: data <= 8'h01; 
        10'b0001111101: data <= 8'h01; 
        10'b0001111110: data <= 8'h01; 
        10'b0001111111: data <= 8'h01; 
        10'b0010000000: data <= 8'h00; 
        10'b0010000001: data <= 8'h00; 
        10'b0010000010: data <= 8'h01; 
        10'b0010000011: data <= 8'h00; 
        10'b0010000100: data <= 8'h00; 
        10'b0010000101: data <= 8'hff; 
        10'b0010000110: data <= 8'hff; 
        10'b0010000111: data <= 8'hff; 
        10'b0010001000: data <= 8'h00; 
        10'b0010001001: data <= 8'h00; 
        10'b0010001010: data <= 8'h00; 
        10'b0010001011: data <= 8'h00; 
        10'b0010001100: data <= 8'h00; 
        10'b0010001101: data <= 8'h00; 
        10'b0010001110: data <= 8'h00; 
        10'b0010001111: data <= 8'h00; 
        10'b0010010000: data <= 8'h00; 
        10'b0010010001: data <= 8'h00; 
        10'b0010010010: data <= 8'h01; 
        10'b0010010011: data <= 8'h01; 
        10'b0010010100: data <= 8'h01; 
        10'b0010010101: data <= 8'h01; 
        10'b0010010110: data <= 8'h00; 
        10'b0010010111: data <= 8'h01; 
        10'b0010011000: data <= 8'h01; 
        10'b0010011001: data <= 8'h01; 
        10'b0010011010: data <= 8'h00; 
        10'b0010011011: data <= 8'h01; 
        10'b0010011100: data <= 8'h01; 
        10'b0010011101: data <= 8'h00; 
        10'b0010011110: data <= 8'h00; 
        10'b0010011111: data <= 8'h00; 
        10'b0010100000: data <= 8'h00; 
        10'b0010100001: data <= 8'hff; 
        10'b0010100010: data <= 8'hff; 
        10'b0010100011: data <= 8'hff; 
        10'b0010100100: data <= 8'h00; 
        10'b0010100101: data <= 8'h00; 
        10'b0010100110: data <= 8'h00; 
        10'b0010100111: data <= 8'h00; 
        10'b0010101000: data <= 8'h00; 
        10'b0010101001: data <= 8'h00; 
        10'b0010101010: data <= 8'h00; 
        10'b0010101011: data <= 8'h00; 
        10'b0010101100: data <= 8'h00; 
        10'b0010101101: data <= 8'h01; 
        10'b0010101110: data <= 8'h01; 
        10'b0010101111: data <= 8'h01; 
        10'b0010110000: data <= 8'h01; 
        10'b0010110001: data <= 8'h01; 
        10'b0010110010: data <= 8'h01; 
        10'b0010110011: data <= 8'h01; 
        10'b0010110100: data <= 8'h01; 
        10'b0010110101: data <= 8'h01; 
        10'b0010110110: data <= 8'h01; 
        10'b0010110111: data <= 8'h00; 
        10'b0010111000: data <= 8'h01; 
        10'b0010111001: data <= 8'h01; 
        10'b0010111010: data <= 8'h01; 
        10'b0010111011: data <= 8'h00; 
        10'b0010111100: data <= 8'h00; 
        10'b0010111101: data <= 8'h00; 
        10'b0010111110: data <= 8'hff; 
        10'b0010111111: data <= 8'hff; 
        10'b0011000000: data <= 8'hff; 
        10'b0011000001: data <= 8'h00; 
        10'b0011000010: data <= 8'h00; 
        10'b0011000011: data <= 8'h00; 
        10'b0011000100: data <= 8'h00; 
        10'b0011000101: data <= 8'h00; 
        10'b0011000110: data <= 8'h00; 
        10'b0011000111: data <= 8'h00; 
        10'b0011001000: data <= 8'h01; 
        10'b0011001001: data <= 8'h01; 
        10'b0011001010: data <= 8'h01; 
        10'b0011001011: data <= 8'h00; 
        10'b0011001100: data <= 8'h00; 
        10'b0011001101: data <= 8'h00; 
        10'b0011001110: data <= 8'h00; 
        10'b0011001111: data <= 8'h00; 
        10'b0011010000: data <= 8'h01; 
        10'b0011010001: data <= 8'h01; 
        10'b0011010010: data <= 8'h01; 
        10'b0011010011: data <= 8'h01; 
        10'b0011010100: data <= 8'h00; 
        10'b0011010101: data <= 8'h00; 
        10'b0011010110: data <= 8'h00; 
        10'b0011010111: data <= 8'h00; 
        10'b0011011000: data <= 8'h00; 
        10'b0011011001: data <= 8'h00; 
        10'b0011011010: data <= 8'h00; 
        10'b0011011011: data <= 8'hff; 
        10'b0011011100: data <= 8'hff; 
        10'b0011011101: data <= 8'h00; 
        10'b0011011110: data <= 8'h00; 
        10'b0011011111: data <= 8'h00; 
        10'b0011100000: data <= 8'h00; 
        10'b0011100001: data <= 8'h00; 
        10'b0011100010: data <= 8'h00; 
        10'b0011100011: data <= 8'h00; 
        10'b0011100100: data <= 8'h01; 
        10'b0011100101: data <= 8'h01; 
        10'b0011100110: data <= 8'h01; 
        10'b0011100111: data <= 8'h00; 
        10'b0011101000: data <= 8'h00; 
        10'b0011101001: data <= 8'h00; 
        10'b0011101010: data <= 8'h01; 
        10'b0011101011: data <= 8'h00; 
        10'b0011101100: data <= 8'h00; 
        10'b0011101101: data <= 8'h00; 
        10'b0011101110: data <= 8'h01; 
        10'b0011101111: data <= 8'h01; 
        10'b0011110000: data <= 8'h00; 
        10'b0011110001: data <= 8'h00; 
        10'b0011110010: data <= 8'h01; 
        10'b0011110011: data <= 8'h00; 
        10'b0011110100: data <= 8'h01; 
        10'b0011110101: data <= 8'h00; 
        10'b0011110110: data <= 8'h00; 
        10'b0011110111: data <= 8'hff; 
        10'b0011111000: data <= 8'hff; 
        10'b0011111001: data <= 8'h00; 
        10'b0011111010: data <= 8'h00; 
        10'b0011111011: data <= 8'h00; 
        10'b0011111100: data <= 8'h00; 
        10'b0011111101: data <= 8'h00; 
        10'b0011111110: data <= 8'h00; 
        10'b0011111111: data <= 8'h00; 
        10'b0100000000: data <= 8'h00; 
        10'b0100000001: data <= 8'h01; 
        10'b0100000010: data <= 8'h00; 
        10'b0100000011: data <= 8'h00; 
        10'b0100000100: data <= 8'h00; 
        10'b0100000101: data <= 8'h00; 
        10'b0100000110: data <= 8'hff; 
        10'b0100000111: data <= 8'hfe; 
        10'b0100001000: data <= 8'hff; 
        10'b0100001001: data <= 8'h00; 
        10'b0100001010: data <= 8'h01; 
        10'b0100001011: data <= 8'h02; 
        10'b0100001100: data <= 8'h01; 
        10'b0100001101: data <= 8'h01; 
        10'b0100001110: data <= 8'h01; 
        10'b0100001111: data <= 8'h01; 
        10'b0100010000: data <= 8'h01; 
        10'b0100010001: data <= 8'h01; 
        10'b0100010010: data <= 8'h00; 
        10'b0100010011: data <= 8'hff; 
        10'b0100010100: data <= 8'h00; 
        10'b0100010101: data <= 8'h00; 
        10'b0100010110: data <= 8'h00; 
        10'b0100010111: data <= 8'h00; 
        10'b0100011000: data <= 8'h00; 
        10'b0100011001: data <= 8'h00; 
        10'b0100011010: data <= 8'h00; 
        10'b0100011011: data <= 8'h00; 
        10'b0100011100: data <= 8'h00; 
        10'b0100011101: data <= 8'h00; 
        10'b0100011110: data <= 8'h00; 
        10'b0100011111: data <= 8'hff; 
        10'b0100100000: data <= 8'hff; 
        10'b0100100001: data <= 8'hfe; 
        10'b0100100010: data <= 8'hfe; 
        10'b0100100011: data <= 8'hfe; 
        10'b0100100100: data <= 8'hfe; 
        10'b0100100101: data <= 8'h00; 
        10'b0100100110: data <= 8'h01; 
        10'b0100100111: data <= 8'h01; 
        10'b0100101000: data <= 8'h01; 
        10'b0100101001: data <= 8'h01; 
        10'b0100101010: data <= 8'h01; 
        10'b0100101011: data <= 8'h01; 
        10'b0100101100: data <= 8'h01; 
        10'b0100101101: data <= 8'h00; 
        10'b0100101110: data <= 8'h00; 
        10'b0100101111: data <= 8'hff; 
        10'b0100110000: data <= 8'h00; 
        10'b0100110001: data <= 8'h00; 
        10'b0100110010: data <= 8'h00; 
        10'b0100110011: data <= 8'h00; 
        10'b0100110100: data <= 8'h00; 
        10'b0100110101: data <= 8'h00; 
        10'b0100110110: data <= 8'h00; 
        10'b0100110111: data <= 8'h00; 
        10'b0100111000: data <= 8'h00; 
        10'b0100111001: data <= 8'hff; 
        10'b0100111010: data <= 8'hff; 
        10'b0100111011: data <= 8'hfe; 
        10'b0100111100: data <= 8'hfe; 
        10'b0100111101: data <= 8'hfe; 
        10'b0100111110: data <= 8'hff; 
        10'b0100111111: data <= 8'hff; 
        10'b0101000000: data <= 8'h00; 
        10'b0101000001: data <= 8'h00; 
        10'b0101000010: data <= 8'h01; 
        10'b0101000011: data <= 8'h01; 
        10'b0101000100: data <= 8'h00; 
        10'b0101000101: data <= 8'h01; 
        10'b0101000110: data <= 8'h01; 
        10'b0101000111: data <= 8'h01; 
        10'b0101001000: data <= 8'h01; 
        10'b0101001001: data <= 8'h00; 
        10'b0101001010: data <= 8'h00; 
        10'b0101001011: data <= 8'h00; 
        10'b0101001100: data <= 8'h00; 
        10'b0101001101: data <= 8'h00; 
        10'b0101001110: data <= 8'h00; 
        10'b0101001111: data <= 8'h00; 
        10'b0101010000: data <= 8'h00; 
        10'b0101010001: data <= 8'h00; 
        10'b0101010010: data <= 8'h00; 
        10'b0101010011: data <= 8'h00; 
        10'b0101010100: data <= 8'h00; 
        10'b0101010101: data <= 8'hff; 
        10'b0101010110: data <= 8'hff; 
        10'b0101010111: data <= 8'hfe; 
        10'b0101011000: data <= 8'hff; 
        10'b0101011001: data <= 8'hff; 
        10'b0101011010: data <= 8'h00; 
        10'b0101011011: data <= 8'h00; 
        10'b0101011100: data <= 8'h00; 
        10'b0101011101: data <= 8'h00; 
        10'b0101011110: data <= 8'h01; 
        10'b0101011111: data <= 8'h01; 
        10'b0101100000: data <= 8'h00; 
        10'b0101100001: data <= 8'h01; 
        10'b0101100010: data <= 8'h00; 
        10'b0101100011: data <= 8'h00; 
        10'b0101100100: data <= 8'hff; 
        10'b0101100101: data <= 8'hff; 
        10'b0101100110: data <= 8'hff; 
        10'b0101100111: data <= 8'hff; 
        10'b0101101000: data <= 8'h00; 
        10'b0101101001: data <= 8'h00; 
        10'b0101101010: data <= 8'h00; 
        10'b0101101011: data <= 8'h00; 
        10'b0101101100: data <= 8'h00; 
        10'b0101101101: data <= 8'h00; 
        10'b0101101110: data <= 8'h00; 
        10'b0101101111: data <= 8'h00; 
        10'b0101110000: data <= 8'h00; 
        10'b0101110001: data <= 8'h00; 
        10'b0101110010: data <= 8'hff; 
        10'b0101110011: data <= 8'hff; 
        10'b0101110100: data <= 8'hff; 
        10'b0101110101: data <= 8'h00; 
        10'b0101110110: data <= 8'h00; 
        10'b0101110111: data <= 8'hff; 
        10'b0101111000: data <= 8'h00; 
        10'b0101111001: data <= 8'h01; 
        10'b0101111010: data <= 8'h01; 
        10'b0101111011: data <= 8'h00; 
        10'b0101111100: data <= 8'h00; 
        10'b0101111101: data <= 8'h00; 
        10'b0101111110: data <= 8'h00; 
        10'b0101111111: data <= 8'h00; 
        10'b0110000000: data <= 8'hff; 
        10'b0110000001: data <= 8'hff; 
        10'b0110000010: data <= 8'hff; 
        10'b0110000011: data <= 8'h00; 
        10'b0110000100: data <= 8'h00; 
        10'b0110000101: data <= 8'h00; 
        10'b0110000110: data <= 8'h00; 
        10'b0110000111: data <= 8'h00; 
        10'b0110001000: data <= 8'h00; 
        10'b0110001001: data <= 8'h00; 
        10'b0110001010: data <= 8'h00; 
        10'b0110001011: data <= 8'h00; 
        10'b0110001100: data <= 8'h00; 
        10'b0110001101: data <= 8'h00; 
        10'b0110001110: data <= 8'hff; 
        10'b0110001111: data <= 8'hff; 
        10'b0110010000: data <= 8'hff; 
        10'b0110010001: data <= 8'h00; 
        10'b0110010010: data <= 8'hff; 
        10'b0110010011: data <= 8'hff; 
        10'b0110010100: data <= 8'h00; 
        10'b0110010101: data <= 8'h00; 
        10'b0110010110: data <= 8'h00; 
        10'b0110010111: data <= 8'h00; 
        10'b0110011000: data <= 8'h00; 
        10'b0110011001: data <= 8'h00; 
        10'b0110011010: data <= 8'h00; 
        10'b0110011011: data <= 8'h00; 
        10'b0110011100: data <= 8'hff; 
        10'b0110011101: data <= 8'h00; 
        10'b0110011110: data <= 8'h00; 
        10'b0110011111: data <= 8'h00; 
        10'b0110100000: data <= 8'h00; 
        10'b0110100001: data <= 8'h00; 
        10'b0110100010: data <= 8'h00; 
        10'b0110100011: data <= 8'h00; 
        10'b0110100100: data <= 8'h00; 
        10'b0110100101: data <= 8'h00; 
        10'b0110100110: data <= 8'h00; 
        10'b0110100111: data <= 8'h00; 
        10'b0110101000: data <= 8'h00; 
        10'b0110101001: data <= 8'h00; 
        10'b0110101010: data <= 8'hff; 
        10'b0110101011: data <= 8'hff; 
        10'b0110101100: data <= 8'hff; 
        10'b0110101101: data <= 8'h00; 
        10'b0110101110: data <= 8'h00; 
        10'b0110101111: data <= 8'h00; 
        10'b0110110000: data <= 8'h00; 
        10'b0110110001: data <= 8'h01; 
        10'b0110110010: data <= 8'h00; 
        10'b0110110011: data <= 8'h00; 
        10'b0110110100: data <= 8'hff; 
        10'b0110110101: data <= 8'h00; 
        10'b0110110110: data <= 8'h00; 
        10'b0110110111: data <= 8'h00; 
        10'b0110111000: data <= 8'h00; 
        10'b0110111001: data <= 8'h00; 
        10'b0110111010: data <= 8'h00; 
        10'b0110111011: data <= 8'h00; 
        10'b0110111100: data <= 8'h00; 
        10'b0110111101: data <= 8'h00; 
        10'b0110111110: data <= 8'h00; 
        10'b0110111111: data <= 8'h00; 
        10'b0111000000: data <= 8'h00; 
        10'b0111000001: data <= 8'h00; 
        10'b0111000010: data <= 8'h00; 
        10'b0111000011: data <= 8'h00; 
        10'b0111000100: data <= 8'h00; 
        10'b0111000101: data <= 8'h00; 
        10'b0111000110: data <= 8'h00; 
        10'b0111000111: data <= 8'hff; 
        10'b0111001000: data <= 8'hff; 
        10'b0111001001: data <= 8'hff; 
        10'b0111001010: data <= 8'hff; 
        10'b0111001011: data <= 8'h00; 
        10'b0111001100: data <= 8'h00; 
        10'b0111001101: data <= 8'h01; 
        10'b0111001110: data <= 8'h00; 
        10'b0111001111: data <= 8'hff; 
        10'b0111010000: data <= 8'hff; 
        10'b0111010001: data <= 8'h00; 
        10'b0111010010: data <= 8'h00; 
        10'b0111010011: data <= 8'h01; 
        10'b0111010100: data <= 8'h01; 
        10'b0111010101: data <= 8'h01; 
        10'b0111010110: data <= 8'h01; 
        10'b0111010111: data <= 8'h00; 
        10'b0111011000: data <= 8'h00; 
        10'b0111011001: data <= 8'h00; 
        10'b0111011010: data <= 8'h00; 
        10'b0111011011: data <= 8'h00; 
        10'b0111011100: data <= 8'h00; 
        10'b0111011101: data <= 8'h00; 
        10'b0111011110: data <= 8'h00; 
        10'b0111011111: data <= 8'h00; 
        10'b0111100000: data <= 8'h00; 
        10'b0111100001: data <= 8'h00; 
        10'b0111100010: data <= 8'h00; 
        10'b0111100011: data <= 8'hff; 
        10'b0111100100: data <= 8'hff; 
        10'b0111100101: data <= 8'hfe; 
        10'b0111100110: data <= 8'hfd; 
        10'b0111100111: data <= 8'hfd; 
        10'b0111101000: data <= 8'hfe; 
        10'b0111101001: data <= 8'hff; 
        10'b0111101010: data <= 8'hff; 
        10'b0111101011: data <= 8'hff; 
        10'b0111101100: data <= 8'h00; 
        10'b0111101101: data <= 8'h00; 
        10'b0111101110: data <= 8'h01; 
        10'b0111101111: data <= 8'h01; 
        10'b0111110000: data <= 8'h00; 
        10'b0111110001: data <= 8'h01; 
        10'b0111110010: data <= 8'h01; 
        10'b0111110011: data <= 8'h00; 
        10'b0111110100: data <= 8'h00; 
        10'b0111110101: data <= 8'h00; 
        10'b0111110110: data <= 8'h00; 
        10'b0111110111: data <= 8'h00; 
        10'b0111111000: data <= 8'h00; 
        10'b0111111001: data <= 8'h00; 
        10'b0111111010: data <= 8'h00; 
        10'b0111111011: data <= 8'h01; 
        10'b0111111100: data <= 8'h00; 
        10'b0111111101: data <= 8'h00; 
        10'b0111111110: data <= 8'h00; 
        10'b0111111111: data <= 8'h00; 
        10'b1000000000: data <= 8'h00; 
        10'b1000000001: data <= 8'hfe; 
        10'b1000000010: data <= 8'hfe; 
        10'b1000000011: data <= 8'hfe; 
        10'b1000000100: data <= 8'hfd; 
        10'b1000000101: data <= 8'hfe; 
        10'b1000000110: data <= 8'hff; 
        10'b1000000111: data <= 8'h00; 
        10'b1000001000: data <= 8'h01; 
        10'b1000001001: data <= 8'h01; 
        10'b1000001010: data <= 8'h01; 
        10'b1000001011: data <= 8'h01; 
        10'b1000001100: data <= 8'h01; 
        10'b1000001101: data <= 8'h01; 
        10'b1000001110: data <= 8'h01; 
        10'b1000001111: data <= 8'h00; 
        10'b1000010000: data <= 8'h00; 
        10'b1000010001: data <= 8'h00; 
        10'b1000010010: data <= 8'h00; 
        10'b1000010011: data <= 8'h00; 
        10'b1000010100: data <= 8'h00; 
        10'b1000010101: data <= 8'h00; 
        10'b1000010110: data <= 8'h00; 
        10'b1000010111: data <= 8'h01; 
        10'b1000011000: data <= 8'h01; 
        10'b1000011001: data <= 8'h01; 
        10'b1000011010: data <= 8'h01; 
        10'b1000011011: data <= 8'h00; 
        10'b1000011100: data <= 8'h00; 
        10'b1000011101: data <= 8'h00; 
        10'b1000011110: data <= 8'h00; 
        10'b1000011111: data <= 8'hff; 
        10'b1000100000: data <= 8'hff; 
        10'b1000100001: data <= 8'hff; 
        10'b1000100010: data <= 8'hff; 
        10'b1000100011: data <= 8'h00; 
        10'b1000100100: data <= 8'h01; 
        10'b1000100101: data <= 8'h01; 
        10'b1000100110: data <= 8'h01; 
        10'b1000100111: data <= 8'h01; 
        10'b1000101000: data <= 8'h01; 
        10'b1000101001: data <= 8'h01; 
        10'b1000101010: data <= 8'h00; 
        10'b1000101011: data <= 8'h00; 
        10'b1000101100: data <= 8'h00; 
        10'b1000101101: data <= 8'h00; 
        10'b1000101110: data <= 8'h00; 
        10'b1000101111: data <= 8'h00; 
        10'b1000110000: data <= 8'h00; 
        10'b1000110001: data <= 8'h00; 
        10'b1000110010: data <= 8'h00; 
        10'b1000110011: data <= 8'h01; 
        10'b1000110100: data <= 8'h01; 
        10'b1000110101: data <= 8'h01; 
        10'b1000110110: data <= 8'h01; 
        10'b1000110111: data <= 8'h01; 
        10'b1000111000: data <= 8'h01; 
        10'b1000111001: data <= 8'h01; 
        10'b1000111010: data <= 8'h00; 
        10'b1000111011: data <= 8'h00; 
        10'b1000111100: data <= 8'h00; 
        10'b1000111101: data <= 8'h00; 
        10'b1000111110: data <= 8'h00; 
        10'b1000111111: data <= 8'h00; 
        10'b1001000000: data <= 8'h00; 
        10'b1001000001: data <= 8'h01; 
        10'b1001000010: data <= 8'h01; 
        10'b1001000011: data <= 8'h01; 
        10'b1001000100: data <= 8'h01; 
        10'b1001000101: data <= 8'h01; 
        10'b1001000110: data <= 8'h00; 
        10'b1001000111: data <= 8'h00; 
        10'b1001001000: data <= 8'h00; 
        10'b1001001001: data <= 8'h00; 
        10'b1001001010: data <= 8'h00; 
        10'b1001001011: data <= 8'h00; 
        10'b1001001100: data <= 8'h00; 
        10'b1001001101: data <= 8'h00; 
        10'b1001001110: data <= 8'h00; 
        10'b1001001111: data <= 8'h00; 
        10'b1001010000: data <= 8'h01; 
        10'b1001010001: data <= 8'h01; 
        10'b1001010010: data <= 8'h01; 
        10'b1001010011: data <= 8'h01; 
        10'b1001010100: data <= 8'h01; 
        10'b1001010101: data <= 8'h00; 
        10'b1001010110: data <= 8'h00; 
        10'b1001010111: data <= 8'h00; 
        10'b1001011000: data <= 8'h00; 
        10'b1001011001: data <= 8'h00; 
        10'b1001011010: data <= 8'h00; 
        10'b1001011011: data <= 8'h00; 
        10'b1001011100: data <= 8'h00; 
        10'b1001011101: data <= 8'h00; 
        10'b1001011110: data <= 8'h00; 
        10'b1001011111: data <= 8'h01; 
        10'b1001100000: data <= 8'h00; 
        10'b1001100001: data <= 8'h00; 
        10'b1001100010: data <= 8'h00; 
        10'b1001100011: data <= 8'h00; 
        10'b1001100100: data <= 8'h00; 
        10'b1001100101: data <= 8'h00; 
        10'b1001100110: data <= 8'h00; 
        10'b1001100111: data <= 8'h00; 
        10'b1001101000: data <= 8'h00; 
        10'b1001101001: data <= 8'h00; 
        10'b1001101010: data <= 8'h00; 
        10'b1001101011: data <= 8'h00; 
        10'b1001101100: data <= 8'h01; 
        10'b1001101101: data <= 8'h01; 
        10'b1001101110: data <= 8'h01; 
        10'b1001101111: data <= 8'h00; 
        10'b1001110000: data <= 8'h00; 
        10'b1001110001: data <= 8'h00; 
        10'b1001110010: data <= 8'h00; 
        10'b1001110011: data <= 8'h00; 
        10'b1001110100: data <= 8'h00; 
        10'b1001110101: data <= 8'h00; 
        10'b1001110110: data <= 8'h00; 
        10'b1001110111: data <= 8'h00; 
        10'b1001111000: data <= 8'h00; 
        10'b1001111001: data <= 8'h00; 
        10'b1001111010: data <= 8'h00; 
        10'b1001111011: data <= 8'h01; 
        10'b1001111100: data <= 8'h00; 
        10'b1001111101: data <= 8'h00; 
        10'b1001111110: data <= 8'h00; 
        10'b1001111111: data <= 8'h00; 
        10'b1010000000: data <= 8'h00; 
        10'b1010000001: data <= 8'h00; 
        10'b1010000010: data <= 8'h00; 
        10'b1010000011: data <= 8'h00; 
        10'b1010000100: data <= 8'h00; 
        10'b1010000101: data <= 8'h00; 
        10'b1010000110: data <= 8'h00; 
        10'b1010000111: data <= 8'h00; 
        10'b1010001000: data <= 8'h01; 
        10'b1010001001: data <= 8'h01; 
        10'b1010001010: data <= 8'h01; 
        10'b1010001011: data <= 8'h01; 
        10'b1010001100: data <= 8'h00; 
        10'b1010001101: data <= 8'h00; 
        10'b1010001110: data <= 8'h00; 
        10'b1010001111: data <= 8'h00; 
        10'b1010010000: data <= 8'h00; 
        10'b1010010001: data <= 8'h00; 
        10'b1010010010: data <= 8'h00; 
        10'b1010010011: data <= 8'h00; 
        10'b1010010100: data <= 8'h00; 
        10'b1010010101: data <= 8'h00; 
        10'b1010010110: data <= 8'h01; 
        10'b1010010111: data <= 8'h00; 
        10'b1010011000: data <= 8'h00; 
        10'b1010011001: data <= 8'h00; 
        10'b1010011010: data <= 8'h00; 
        10'b1010011011: data <= 8'h00; 
        10'b1010011100: data <= 8'h00; 
        10'b1010011101: data <= 8'h00; 
        10'b1010011110: data <= 8'h00; 
        10'b1010011111: data <= 8'h00; 
        10'b1010100000: data <= 8'h00; 
        10'b1010100001: data <= 8'h00; 
        10'b1010100010: data <= 8'h00; 
        10'b1010100011: data <= 8'h00; 
        10'b1010100100: data <= 8'h00; 
        10'b1010100101: data <= 8'h01; 
        10'b1010100110: data <= 8'h01; 
        10'b1010100111: data <= 8'h01; 
        10'b1010101000: data <= 8'h01; 
        10'b1010101001: data <= 8'h01; 
        10'b1010101010: data <= 8'h01; 
        10'b1010101011: data <= 8'h01; 
        10'b1010101100: data <= 8'h01; 
        10'b1010101101: data <= 8'h01; 
        10'b1010101110: data <= 8'h01; 
        10'b1010101111: data <= 8'h01; 
        10'b1010110000: data <= 8'h01; 
        10'b1010110001: data <= 8'h00; 
        10'b1010110010: data <= 8'h00; 
        10'b1010110011: data <= 8'hff; 
        10'b1010110100: data <= 8'hff; 
        10'b1010110101: data <= 8'h00; 
        10'b1010110110: data <= 8'h00; 
        10'b1010110111: data <= 8'h00; 
        10'b1010111000: data <= 8'h00; 
        10'b1010111001: data <= 8'h00; 
        10'b1010111010: data <= 8'h00; 
        10'b1010111011: data <= 8'h00; 
        10'b1010111100: data <= 8'h00; 
        10'b1010111101: data <= 8'h00; 
        10'b1010111110: data <= 8'h00; 
        10'b1010111111: data <= 8'h00; 
        10'b1011000000: data <= 8'h00; 
        10'b1011000001: data <= 8'h00; 
        10'b1011000010: data <= 8'h00; 
        10'b1011000011: data <= 8'h00; 
        10'b1011000100: data <= 8'h00; 
        10'b1011000101: data <= 8'h00; 
        10'b1011000110: data <= 8'h01; 
        10'b1011000111: data <= 8'h01; 
        10'b1011001000: data <= 8'h01; 
        10'b1011001001: data <= 8'h01; 
        10'b1011001010: data <= 8'h01; 
        10'b1011001011: data <= 8'h00; 
        10'b1011001100: data <= 8'h00; 
        10'b1011001101: data <= 8'h00; 
        10'b1011001110: data <= 8'h00; 
        10'b1011001111: data <= 8'h00; 
        10'b1011010000: data <= 8'h00; 
        10'b1011010001: data <= 8'h00; 
        10'b1011010010: data <= 8'h00; 
        10'b1011010011: data <= 8'h00; 
        10'b1011010100: data <= 8'h00; 
        10'b1011010101: data <= 8'h00; 
        10'b1011010110: data <= 8'h00; 
        10'b1011010111: data <= 8'h00; 
        10'b1011011000: data <= 8'h00; 
        10'b1011011001: data <= 8'h00; 
        10'b1011011010: data <= 8'h00; 
        10'b1011011011: data <= 8'h00; 
        10'b1011011100: data <= 8'h00; 
        10'b1011011101: data <= 8'h00; 
        10'b1011011110: data <= 8'h00; 
        10'b1011011111: data <= 8'h00; 
        10'b1011100000: data <= 8'h00; 
        10'b1011100001: data <= 8'h00; 
        10'b1011100010: data <= 8'h00; 
        10'b1011100011: data <= 8'h00; 
        10'b1011100100: data <= 8'h00; 
        10'b1011100101: data <= 8'h00; 
        10'b1011100110: data <= 8'h00; 
        10'b1011100111: data <= 8'h00; 
        10'b1011101000: data <= 8'h00; 
        10'b1011101001: data <= 8'h00; 
        10'b1011101010: data <= 8'h00; 
        10'b1011101011: data <= 8'h00; 
        10'b1011101100: data <= 8'h00; 
        10'b1011101101: data <= 8'h00; 
        10'b1011101110: data <= 8'h00; 
        10'b1011101111: data <= 8'h00; 
        10'b1011110000: data <= 8'h00; 
        10'b1011110001: data <= 8'h00; 
        10'b1011110010: data <= 8'h00; 
        10'b1011110011: data <= 8'h00; 
        10'b1011110100: data <= 8'h00; 
        10'b1011110101: data <= 8'h00; 
        10'b1011110110: data <= 8'h00; 
        10'b1011110111: data <= 8'h00; 
        10'b1011111000: data <= 8'h00; 
        10'b1011111001: data <= 8'h00; 
        10'b1011111010: data <= 8'h00; 
        10'b1011111011: data <= 8'h00; 
        10'b1011111100: data <= 8'h00; 
        10'b1011111101: data <= 8'h00; 
        10'b1011111110: data <= 8'h00; 
        10'b1011111111: data <= 8'h00; 
        10'b1100000000: data <= 8'h00; 
        10'b1100000001: data <= 8'h00; 
        10'b1100000010: data <= 8'h00; 
        10'b1100000011: data <= 8'h00; 
        10'b1100000100: data <= 8'h00; 
        10'b1100000101: data <= 8'h00; 
        10'b1100000110: data <= 8'h00; 
        10'b1100000111: data <= 8'h00; 
        10'b1100001000: data <= 8'h00; 
        10'b1100001001: data <= 8'h00; 
        10'b1100001010: data <= 8'h00; 
        10'b1100001011: data <= 8'h00; 
        10'b1100001100: data <= 8'h00; 
        10'b1100001101: data <= 8'h00; 
        10'b1100001110: data <= 8'h00; 
        10'b1100001111: data <= 8'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 3) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 9'h000; 
        10'b0000000001: data <= 9'h000; 
        10'b0000000010: data <= 9'h000; 
        10'b0000000011: data <= 9'h000; 
        10'b0000000100: data <= 9'h000; 
        10'b0000000101: data <= 9'h000; 
        10'b0000000110: data <= 9'h000; 
        10'b0000000111: data <= 9'h000; 
        10'b0000001000: data <= 9'h000; 
        10'b0000001001: data <= 9'h000; 
        10'b0000001010: data <= 9'h000; 
        10'b0000001011: data <= 9'h000; 
        10'b0000001100: data <= 9'h000; 
        10'b0000001101: data <= 9'h000; 
        10'b0000001110: data <= 9'h000; 
        10'b0000001111: data <= 9'h000; 
        10'b0000010000: data <= 9'h000; 
        10'b0000010001: data <= 9'h000; 
        10'b0000010010: data <= 9'h000; 
        10'b0000010011: data <= 9'h000; 
        10'b0000010100: data <= 9'h000; 
        10'b0000010101: data <= 9'h000; 
        10'b0000010110: data <= 9'h1ff; 
        10'b0000010111: data <= 9'h000; 
        10'b0000011000: data <= 9'h000; 
        10'b0000011001: data <= 9'h000; 
        10'b0000011010: data <= 9'h000; 
        10'b0000011011: data <= 9'h000; 
        10'b0000011100: data <= 9'h000; 
        10'b0000011101: data <= 9'h000; 
        10'b0000011110: data <= 9'h000; 
        10'b0000011111: data <= 9'h000; 
        10'b0000100000: data <= 9'h000; 
        10'b0000100001: data <= 9'h000; 
        10'b0000100010: data <= 9'h000; 
        10'b0000100011: data <= 9'h000; 
        10'b0000100100: data <= 9'h000; 
        10'b0000100101: data <= 9'h1ff; 
        10'b0000100110: data <= 9'h000; 
        10'b0000100111: data <= 9'h000; 
        10'b0000101000: data <= 9'h000; 
        10'b0000101001: data <= 9'h000; 
        10'b0000101010: data <= 9'h000; 
        10'b0000101011: data <= 9'h000; 
        10'b0000101100: data <= 9'h000; 
        10'b0000101101: data <= 9'h000; 
        10'b0000101110: data <= 9'h000; 
        10'b0000101111: data <= 9'h000; 
        10'b0000110000: data <= 9'h000; 
        10'b0000110001: data <= 9'h000; 
        10'b0000110010: data <= 9'h000; 
        10'b0000110011: data <= 9'h000; 
        10'b0000110100: data <= 9'h000; 
        10'b0000110101: data <= 9'h000; 
        10'b0000110110: data <= 9'h000; 
        10'b0000110111: data <= 9'h000; 
        10'b0000111000: data <= 9'h000; 
        10'b0000111001: data <= 9'h000; 
        10'b0000111010: data <= 9'h000; 
        10'b0000111011: data <= 9'h000; 
        10'b0000111100: data <= 9'h000; 
        10'b0000111101: data <= 9'h000; 
        10'b0000111110: data <= 9'h000; 
        10'b0000111111: data <= 9'h000; 
        10'b0001000000: data <= 9'h000; 
        10'b0001000001: data <= 9'h000; 
        10'b0001000010: data <= 9'h000; 
        10'b0001000011: data <= 9'h000; 
        10'b0001000100: data <= 9'h000; 
        10'b0001000101: data <= 9'h000; 
        10'b0001000110: data <= 9'h000; 
        10'b0001000111: data <= 9'h000; 
        10'b0001001000: data <= 9'h000; 
        10'b0001001001: data <= 9'h000; 
        10'b0001001010: data <= 9'h000; 
        10'b0001001011: data <= 9'h000; 
        10'b0001001100: data <= 9'h000; 
        10'b0001001101: data <= 9'h000; 
        10'b0001001110: data <= 9'h000; 
        10'b0001001111: data <= 9'h000; 
        10'b0001010000: data <= 9'h000; 
        10'b0001010001: data <= 9'h000; 
        10'b0001010010: data <= 9'h000; 
        10'b0001010011: data <= 9'h000; 
        10'b0001010100: data <= 9'h000; 
        10'b0001010101: data <= 9'h000; 
        10'b0001010110: data <= 9'h000; 
        10'b0001010111: data <= 9'h000; 
        10'b0001011000: data <= 9'h000; 
        10'b0001011001: data <= 9'h000; 
        10'b0001011010: data <= 9'h000; 
        10'b0001011011: data <= 9'h000; 
        10'b0001011100: data <= 9'h000; 
        10'b0001011101: data <= 9'h000; 
        10'b0001011110: data <= 9'h000; 
        10'b0001011111: data <= 9'h001; 
        10'b0001100000: data <= 9'h001; 
        10'b0001100001: data <= 9'h001; 
        10'b0001100010: data <= 9'h001; 
        10'b0001100011: data <= 9'h001; 
        10'b0001100100: data <= 9'h001; 
        10'b0001100101: data <= 9'h001; 
        10'b0001100110: data <= 9'h001; 
        10'b0001100111: data <= 9'h000; 
        10'b0001101000: data <= 9'h000; 
        10'b0001101001: data <= 9'h1ff; 
        10'b0001101010: data <= 9'h000; 
        10'b0001101011: data <= 9'h000; 
        10'b0001101100: data <= 9'h000; 
        10'b0001101101: data <= 9'h000; 
        10'b0001101110: data <= 9'h000; 
        10'b0001101111: data <= 9'h000; 
        10'b0001110000: data <= 9'h000; 
        10'b0001110001: data <= 9'h000; 
        10'b0001110010: data <= 9'h000; 
        10'b0001110011: data <= 9'h000; 
        10'b0001110100: data <= 9'h000; 
        10'b0001110101: data <= 9'h000; 
        10'b0001110110: data <= 9'h001; 
        10'b0001110111: data <= 9'h001; 
        10'b0001111000: data <= 9'h002; 
        10'b0001111001: data <= 9'h001; 
        10'b0001111010: data <= 9'h002; 
        10'b0001111011: data <= 9'h002; 
        10'b0001111100: data <= 9'h002; 
        10'b0001111101: data <= 9'h003; 
        10'b0001111110: data <= 9'h002; 
        10'b0001111111: data <= 9'h002; 
        10'b0010000000: data <= 9'h001; 
        10'b0010000001: data <= 9'h001; 
        10'b0010000010: data <= 9'h001; 
        10'b0010000011: data <= 9'h000; 
        10'b0010000100: data <= 9'h1ff; 
        10'b0010000101: data <= 9'h1ff; 
        10'b0010000110: data <= 9'h1ff; 
        10'b0010000111: data <= 9'h1ff; 
        10'b0010001000: data <= 9'h000; 
        10'b0010001001: data <= 9'h000; 
        10'b0010001010: data <= 9'h000; 
        10'b0010001011: data <= 9'h000; 
        10'b0010001100: data <= 9'h000; 
        10'b0010001101: data <= 9'h000; 
        10'b0010001110: data <= 9'h000; 
        10'b0010001111: data <= 9'h000; 
        10'b0010010000: data <= 9'h000; 
        10'b0010010001: data <= 9'h001; 
        10'b0010010010: data <= 9'h001; 
        10'b0010010011: data <= 9'h001; 
        10'b0010010100: data <= 9'h001; 
        10'b0010010101: data <= 9'h001; 
        10'b0010010110: data <= 9'h001; 
        10'b0010010111: data <= 9'h001; 
        10'b0010011000: data <= 9'h001; 
        10'b0010011001: data <= 9'h002; 
        10'b0010011010: data <= 9'h000; 
        10'b0010011011: data <= 9'h001; 
        10'b0010011100: data <= 9'h001; 
        10'b0010011101: data <= 9'h000; 
        10'b0010011110: data <= 9'h000; 
        10'b0010011111: data <= 9'h1ff; 
        10'b0010100000: data <= 9'h1ff; 
        10'b0010100001: data <= 9'h1fe; 
        10'b0010100010: data <= 9'h1fe; 
        10'b0010100011: data <= 9'h1fe; 
        10'b0010100100: data <= 9'h1ff; 
        10'b0010100101: data <= 9'h000; 
        10'b0010100110: data <= 9'h000; 
        10'b0010100111: data <= 9'h000; 
        10'b0010101000: data <= 9'h000; 
        10'b0010101001: data <= 9'h000; 
        10'b0010101010: data <= 9'h000; 
        10'b0010101011: data <= 9'h000; 
        10'b0010101100: data <= 9'h001; 
        10'b0010101101: data <= 9'h002; 
        10'b0010101110: data <= 9'h001; 
        10'b0010101111: data <= 9'h001; 
        10'b0010110000: data <= 9'h002; 
        10'b0010110001: data <= 9'h001; 
        10'b0010110010: data <= 9'h001; 
        10'b0010110011: data <= 9'h001; 
        10'b0010110100: data <= 9'h001; 
        10'b0010110101: data <= 9'h002; 
        10'b0010110110: data <= 9'h001; 
        10'b0010110111: data <= 9'h001; 
        10'b0010111000: data <= 9'h001; 
        10'b0010111001: data <= 9'h001; 
        10'b0010111010: data <= 9'h001; 
        10'b0010111011: data <= 9'h1ff; 
        10'b0010111100: data <= 9'h000; 
        10'b0010111101: data <= 9'h000; 
        10'b0010111110: data <= 9'h1fe; 
        10'b0010111111: data <= 9'h1fe; 
        10'b0011000000: data <= 9'h1ff; 
        10'b0011000001: data <= 9'h000; 
        10'b0011000010: data <= 9'h000; 
        10'b0011000011: data <= 9'h000; 
        10'b0011000100: data <= 9'h000; 
        10'b0011000101: data <= 9'h000; 
        10'b0011000110: data <= 9'h000; 
        10'b0011000111: data <= 9'h001; 
        10'b0011001000: data <= 9'h002; 
        10'b0011001001: data <= 9'h002; 
        10'b0011001010: data <= 9'h001; 
        10'b0011001011: data <= 9'h000; 
        10'b0011001100: data <= 9'h000; 
        10'b0011001101: data <= 9'h001; 
        10'b0011001110: data <= 9'h000; 
        10'b0011001111: data <= 9'h000; 
        10'b0011010000: data <= 9'h001; 
        10'b0011010001: data <= 9'h001; 
        10'b0011010010: data <= 9'h002; 
        10'b0011010011: data <= 9'h001; 
        10'b0011010100: data <= 9'h000; 
        10'b0011010101: data <= 9'h001; 
        10'b0011010110: data <= 9'h001; 
        10'b0011010111: data <= 9'h001; 
        10'b0011011000: data <= 9'h001; 
        10'b0011011001: data <= 9'h000; 
        10'b0011011010: data <= 9'h1ff; 
        10'b0011011011: data <= 9'h1fe; 
        10'b0011011100: data <= 9'h1ff; 
        10'b0011011101: data <= 9'h000; 
        10'b0011011110: data <= 9'h000; 
        10'b0011011111: data <= 9'h000; 
        10'b0011100000: data <= 9'h000; 
        10'b0011100001: data <= 9'h000; 
        10'b0011100010: data <= 9'h000; 
        10'b0011100011: data <= 9'h001; 
        10'b0011100100: data <= 9'h002; 
        10'b0011100101: data <= 9'h002; 
        10'b0011100110: data <= 9'h001; 
        10'b0011100111: data <= 9'h000; 
        10'b0011101000: data <= 9'h001; 
        10'b0011101001: data <= 9'h000; 
        10'b0011101010: data <= 9'h001; 
        10'b0011101011: data <= 9'h000; 
        10'b0011101100: data <= 9'h000; 
        10'b0011101101: data <= 9'h000; 
        10'b0011101110: data <= 9'h002; 
        10'b0011101111: data <= 9'h002; 
        10'b0011110000: data <= 9'h000; 
        10'b0011110001: data <= 9'h001; 
        10'b0011110010: data <= 9'h001; 
        10'b0011110011: data <= 9'h001; 
        10'b0011110100: data <= 9'h001; 
        10'b0011110101: data <= 9'h001; 
        10'b0011110110: data <= 9'h000; 
        10'b0011110111: data <= 9'h1fe; 
        10'b0011111000: data <= 9'h1ff; 
        10'b0011111001: data <= 9'h1ff; 
        10'b0011111010: data <= 9'h000; 
        10'b0011111011: data <= 9'h000; 
        10'b0011111100: data <= 9'h000; 
        10'b0011111101: data <= 9'h000; 
        10'b0011111110: data <= 9'h000; 
        10'b0011111111: data <= 9'h000; 
        10'b0100000000: data <= 9'h001; 
        10'b0100000001: data <= 9'h001; 
        10'b0100000010: data <= 9'h001; 
        10'b0100000011: data <= 9'h000; 
        10'b0100000100: data <= 9'h000; 
        10'b0100000101: data <= 9'h1ff; 
        10'b0100000110: data <= 9'h1fe; 
        10'b0100000111: data <= 9'h1fd; 
        10'b0100001000: data <= 9'h1fd; 
        10'b0100001001: data <= 9'h000; 
        10'b0100001010: data <= 9'h002; 
        10'b0100001011: data <= 9'h004; 
        10'b0100001100: data <= 9'h002; 
        10'b0100001101: data <= 9'h001; 
        10'b0100001110: data <= 9'h001; 
        10'b0100001111: data <= 9'h001; 
        10'b0100010000: data <= 9'h002; 
        10'b0100010001: data <= 9'h001; 
        10'b0100010010: data <= 9'h000; 
        10'b0100010011: data <= 9'h1fe; 
        10'b0100010100: data <= 9'h1ff; 
        10'b0100010101: data <= 9'h1ff; 
        10'b0100010110: data <= 9'h000; 
        10'b0100010111: data <= 9'h000; 
        10'b0100011000: data <= 9'h000; 
        10'b0100011001: data <= 9'h000; 
        10'b0100011010: data <= 9'h000; 
        10'b0100011011: data <= 9'h000; 
        10'b0100011100: data <= 9'h000; 
        10'b0100011101: data <= 9'h000; 
        10'b0100011110: data <= 9'h1ff; 
        10'b0100011111: data <= 9'h1ff; 
        10'b0100100000: data <= 9'h1fd; 
        10'b0100100001: data <= 9'h1fc; 
        10'b0100100010: data <= 9'h1fc; 
        10'b0100100011: data <= 9'h1fb; 
        10'b0100100100: data <= 9'h1fd; 
        10'b0100100101: data <= 9'h1ff; 
        10'b0100100110: data <= 9'h002; 
        10'b0100100111: data <= 9'h002; 
        10'b0100101000: data <= 9'h002; 
        10'b0100101001: data <= 9'h002; 
        10'b0100101010: data <= 9'h001; 
        10'b0100101011: data <= 9'h002; 
        10'b0100101100: data <= 9'h002; 
        10'b0100101101: data <= 9'h001; 
        10'b0100101110: data <= 9'h1ff; 
        10'b0100101111: data <= 9'h1ff; 
        10'b0100110000: data <= 9'h000; 
        10'b0100110001: data <= 9'h1ff; 
        10'b0100110010: data <= 9'h000; 
        10'b0100110011: data <= 9'h000; 
        10'b0100110100: data <= 9'h000; 
        10'b0100110101: data <= 9'h000; 
        10'b0100110110: data <= 9'h000; 
        10'b0100110111: data <= 9'h000; 
        10'b0100111000: data <= 9'h000; 
        10'b0100111001: data <= 9'h1ff; 
        10'b0100111010: data <= 9'h1fe; 
        10'b0100111011: data <= 9'h1fd; 
        10'b0100111100: data <= 9'h1fc; 
        10'b0100111101: data <= 9'h1fd; 
        10'b0100111110: data <= 9'h1fd; 
        10'b0100111111: data <= 9'h1ff; 
        10'b0101000000: data <= 9'h1ff; 
        10'b0101000001: data <= 9'h001; 
        10'b0101000010: data <= 9'h001; 
        10'b0101000011: data <= 9'h001; 
        10'b0101000100: data <= 9'h001; 
        10'b0101000101: data <= 9'h001; 
        10'b0101000110: data <= 9'h002; 
        10'b0101000111: data <= 9'h002; 
        10'b0101001000: data <= 9'h001; 
        10'b0101001001: data <= 9'h000; 
        10'b0101001010: data <= 9'h1ff; 
        10'b0101001011: data <= 9'h1ff; 
        10'b0101001100: data <= 9'h000; 
        10'b0101001101: data <= 9'h000; 
        10'b0101001110: data <= 9'h000; 
        10'b0101001111: data <= 9'h000; 
        10'b0101010000: data <= 9'h000; 
        10'b0101010001: data <= 9'h000; 
        10'b0101010010: data <= 9'h000; 
        10'b0101010011: data <= 9'h000; 
        10'b0101010100: data <= 9'h1ff; 
        10'b0101010101: data <= 9'h1ff; 
        10'b0101010110: data <= 9'h1fe; 
        10'b0101010111: data <= 9'h1fd; 
        10'b0101011000: data <= 9'h1fd; 
        10'b0101011001: data <= 9'h1ff; 
        10'b0101011010: data <= 9'h000; 
        10'b0101011011: data <= 9'h000; 
        10'b0101011100: data <= 9'h000; 
        10'b0101011101: data <= 9'h001; 
        10'b0101011110: data <= 9'h002; 
        10'b0101011111: data <= 9'h001; 
        10'b0101100000: data <= 9'h001; 
        10'b0101100001: data <= 9'h001; 
        10'b0101100010: data <= 9'h001; 
        10'b0101100011: data <= 9'h000; 
        10'b0101100100: data <= 9'h1ff; 
        10'b0101100101: data <= 9'h1fe; 
        10'b0101100110: data <= 9'h1fe; 
        10'b0101100111: data <= 9'h1ff; 
        10'b0101101000: data <= 9'h000; 
        10'b0101101001: data <= 9'h000; 
        10'b0101101010: data <= 9'h000; 
        10'b0101101011: data <= 9'h000; 
        10'b0101101100: data <= 9'h000; 
        10'b0101101101: data <= 9'h000; 
        10'b0101101110: data <= 9'h000; 
        10'b0101101111: data <= 9'h000; 
        10'b0101110000: data <= 9'h1ff; 
        10'b0101110001: data <= 9'h1ff; 
        10'b0101110010: data <= 9'h1fe; 
        10'b0101110011: data <= 9'h1fe; 
        10'b0101110100: data <= 9'h1fe; 
        10'b0101110101: data <= 9'h000; 
        10'b0101110110: data <= 9'h1ff; 
        10'b0101110111: data <= 9'h1ff; 
        10'b0101111000: data <= 9'h000; 
        10'b0101111001: data <= 9'h002; 
        10'b0101111010: data <= 9'h002; 
        10'b0101111011: data <= 9'h000; 
        10'b0101111100: data <= 9'h001; 
        10'b0101111101: data <= 9'h001; 
        10'b0101111110: data <= 9'h000; 
        10'b0101111111: data <= 9'h1ff; 
        10'b0110000000: data <= 9'h1fe; 
        10'b0110000001: data <= 9'h1fe; 
        10'b0110000010: data <= 9'h1ff; 
        10'b0110000011: data <= 9'h1ff; 
        10'b0110000100: data <= 9'h1ff; 
        10'b0110000101: data <= 9'h000; 
        10'b0110000110: data <= 9'h000; 
        10'b0110000111: data <= 9'h000; 
        10'b0110001000: data <= 9'h000; 
        10'b0110001001: data <= 9'h000; 
        10'b0110001010: data <= 9'h000; 
        10'b0110001011: data <= 9'h000; 
        10'b0110001100: data <= 9'h000; 
        10'b0110001101: data <= 9'h1ff; 
        10'b0110001110: data <= 9'h1fe; 
        10'b0110001111: data <= 9'h1fe; 
        10'b0110010000: data <= 9'h1ff; 
        10'b0110010001: data <= 9'h000; 
        10'b0110010010: data <= 9'h1ff; 
        10'b0110010011: data <= 9'h1ff; 
        10'b0110010100: data <= 9'h000; 
        10'b0110010101: data <= 9'h001; 
        10'b0110010110: data <= 9'h001; 
        10'b0110010111: data <= 9'h000; 
        10'b0110011000: data <= 9'h000; 
        10'b0110011001: data <= 9'h000; 
        10'b0110011010: data <= 9'h000; 
        10'b0110011011: data <= 9'h1ff; 
        10'b0110011100: data <= 9'h1ff; 
        10'b0110011101: data <= 9'h1ff; 
        10'b0110011110: data <= 9'h1ff; 
        10'b0110011111: data <= 9'h000; 
        10'b0110100000: data <= 9'h1ff; 
        10'b0110100001: data <= 9'h1ff; 
        10'b0110100010: data <= 9'h000; 
        10'b0110100011: data <= 9'h000; 
        10'b0110100100: data <= 9'h000; 
        10'b0110100101: data <= 9'h000; 
        10'b0110100110: data <= 9'h000; 
        10'b0110100111: data <= 9'h000; 
        10'b0110101000: data <= 9'h000; 
        10'b0110101001: data <= 9'h1ff; 
        10'b0110101010: data <= 9'h1fe; 
        10'b0110101011: data <= 9'h1fe; 
        10'b0110101100: data <= 9'h1ff; 
        10'b0110101101: data <= 9'h1ff; 
        10'b0110101110: data <= 9'h1ff; 
        10'b0110101111: data <= 9'h000; 
        10'b0110110000: data <= 9'h000; 
        10'b0110110001: data <= 9'h001; 
        10'b0110110010: data <= 9'h001; 
        10'b0110110011: data <= 9'h000; 
        10'b0110110100: data <= 9'h1ff; 
        10'b0110110101: data <= 9'h000; 
        10'b0110110110: data <= 9'h000; 
        10'b0110110111: data <= 9'h000; 
        10'b0110111000: data <= 9'h001; 
        10'b0110111001: data <= 9'h001; 
        10'b0110111010: data <= 9'h000; 
        10'b0110111011: data <= 9'h000; 
        10'b0110111100: data <= 9'h000; 
        10'b0110111101: data <= 9'h000; 
        10'b0110111110: data <= 9'h000; 
        10'b0110111111: data <= 9'h000; 
        10'b0111000000: data <= 9'h000; 
        10'b0111000001: data <= 9'h000; 
        10'b0111000010: data <= 9'h000; 
        10'b0111000011: data <= 9'h000; 
        10'b0111000100: data <= 9'h000; 
        10'b0111000101: data <= 9'h000; 
        10'b0111000110: data <= 9'h1ff; 
        10'b0111000111: data <= 9'h1ff; 
        10'b0111001000: data <= 9'h1fd; 
        10'b0111001001: data <= 9'h1fd; 
        10'b0111001010: data <= 9'h1fe; 
        10'b0111001011: data <= 9'h1ff; 
        10'b0111001100: data <= 9'h001; 
        10'b0111001101: data <= 9'h002; 
        10'b0111001110: data <= 9'h000; 
        10'b0111001111: data <= 9'h1ff; 
        10'b0111010000: data <= 9'h1ff; 
        10'b0111010001: data <= 9'h000; 
        10'b0111010010: data <= 9'h001; 
        10'b0111010011: data <= 9'h002; 
        10'b0111010100: data <= 9'h001; 
        10'b0111010101: data <= 9'h001; 
        10'b0111010110: data <= 9'h001; 
        10'b0111010111: data <= 9'h001; 
        10'b0111011000: data <= 9'h000; 
        10'b0111011001: data <= 9'h000; 
        10'b0111011010: data <= 9'h000; 
        10'b0111011011: data <= 9'h000; 
        10'b0111011100: data <= 9'h000; 
        10'b0111011101: data <= 9'h000; 
        10'b0111011110: data <= 9'h000; 
        10'b0111011111: data <= 9'h001; 
        10'b0111100000: data <= 9'h000; 
        10'b0111100001: data <= 9'h000; 
        10'b0111100010: data <= 9'h000; 
        10'b0111100011: data <= 9'h1fe; 
        10'b0111100100: data <= 9'h1fd; 
        10'b0111100101: data <= 9'h1fc; 
        10'b0111100110: data <= 9'h1fa; 
        10'b0111100111: data <= 9'h1fb; 
        10'b0111101000: data <= 9'h1fc; 
        10'b0111101001: data <= 9'h1fe; 
        10'b0111101010: data <= 9'h1fe; 
        10'b0111101011: data <= 9'h1fe; 
        10'b0111101100: data <= 9'h000; 
        10'b0111101101: data <= 9'h001; 
        10'b0111101110: data <= 9'h001; 
        10'b0111101111: data <= 9'h002; 
        10'b0111110000: data <= 9'h000; 
        10'b0111110001: data <= 9'h002; 
        10'b0111110010: data <= 9'h002; 
        10'b0111110011: data <= 9'h001; 
        10'b0111110100: data <= 9'h000; 
        10'b0111110101: data <= 9'h000; 
        10'b0111110110: data <= 9'h000; 
        10'b0111110111: data <= 9'h000; 
        10'b0111111000: data <= 9'h000; 
        10'b0111111001: data <= 9'h000; 
        10'b0111111010: data <= 9'h000; 
        10'b0111111011: data <= 9'h001; 
        10'b0111111100: data <= 9'h001; 
        10'b0111111101: data <= 9'h001; 
        10'b0111111110: data <= 9'h000; 
        10'b0111111111: data <= 9'h000; 
        10'b1000000000: data <= 9'h1ff; 
        10'b1000000001: data <= 9'h1fd; 
        10'b1000000010: data <= 9'h1fb; 
        10'b1000000011: data <= 9'h1fb; 
        10'b1000000100: data <= 9'h1fb; 
        10'b1000000101: data <= 9'h1fc; 
        10'b1000000110: data <= 9'h1fd; 
        10'b1000000111: data <= 9'h1ff; 
        10'b1000001000: data <= 9'h001; 
        10'b1000001001: data <= 9'h002; 
        10'b1000001010: data <= 9'h002; 
        10'b1000001011: data <= 9'h002; 
        10'b1000001100: data <= 9'h001; 
        10'b1000001101: data <= 9'h002; 
        10'b1000001110: data <= 9'h002; 
        10'b1000001111: data <= 9'h001; 
        10'b1000010000: data <= 9'h1ff; 
        10'b1000010001: data <= 9'h1ff; 
        10'b1000010010: data <= 9'h000; 
        10'b1000010011: data <= 9'h000; 
        10'b1000010100: data <= 9'h000; 
        10'b1000010101: data <= 9'h000; 
        10'b1000010110: data <= 9'h000; 
        10'b1000010111: data <= 9'h002; 
        10'b1000011000: data <= 9'h002; 
        10'b1000011001: data <= 9'h002; 
        10'b1000011010: data <= 9'h002; 
        10'b1000011011: data <= 9'h001; 
        10'b1000011100: data <= 9'h000; 
        10'b1000011101: data <= 9'h1ff; 
        10'b1000011110: data <= 9'h000; 
        10'b1000011111: data <= 9'h1fe; 
        10'b1000100000: data <= 9'h1fe; 
        10'b1000100001: data <= 9'h1fe; 
        10'b1000100010: data <= 9'h1fe; 
        10'b1000100011: data <= 9'h001; 
        10'b1000100100: data <= 9'h002; 
        10'b1000100101: data <= 9'h002; 
        10'b1000100110: data <= 9'h002; 
        10'b1000100111: data <= 9'h002; 
        10'b1000101000: data <= 9'h002; 
        10'b1000101001: data <= 9'h002; 
        10'b1000101010: data <= 9'h001; 
        10'b1000101011: data <= 9'h000; 
        10'b1000101100: data <= 9'h1ff; 
        10'b1000101101: data <= 9'h000; 
        10'b1000101110: data <= 9'h000; 
        10'b1000101111: data <= 9'h000; 
        10'b1000110000: data <= 9'h000; 
        10'b1000110001: data <= 9'h000; 
        10'b1000110010: data <= 9'h000; 
        10'b1000110011: data <= 9'h002; 
        10'b1000110100: data <= 9'h002; 
        10'b1000110101: data <= 9'h002; 
        10'b1000110110: data <= 9'h002; 
        10'b1000110111: data <= 9'h001; 
        10'b1000111000: data <= 9'h001; 
        10'b1000111001: data <= 9'h002; 
        10'b1000111010: data <= 9'h001; 
        10'b1000111011: data <= 9'h000; 
        10'b1000111100: data <= 9'h1ff; 
        10'b1000111101: data <= 9'h1ff; 
        10'b1000111110: data <= 9'h000; 
        10'b1000111111: data <= 9'h000; 
        10'b1001000000: data <= 9'h001; 
        10'b1001000001: data <= 9'h002; 
        10'b1001000010: data <= 9'h002; 
        10'b1001000011: data <= 9'h001; 
        10'b1001000100: data <= 9'h002; 
        10'b1001000101: data <= 9'h001; 
        10'b1001000110: data <= 9'h000; 
        10'b1001000111: data <= 9'h000; 
        10'b1001001000: data <= 9'h1ff; 
        10'b1001001001: data <= 9'h000; 
        10'b1001001010: data <= 9'h000; 
        10'b1001001011: data <= 9'h000; 
        10'b1001001100: data <= 9'h000; 
        10'b1001001101: data <= 9'h000; 
        10'b1001001110: data <= 9'h000; 
        10'b1001001111: data <= 9'h001; 
        10'b1001010000: data <= 9'h002; 
        10'b1001010001: data <= 9'h002; 
        10'b1001010010: data <= 9'h002; 
        10'b1001010011: data <= 9'h001; 
        10'b1001010100: data <= 9'h001; 
        10'b1001010101: data <= 9'h000; 
        10'b1001010110: data <= 9'h000; 
        10'b1001010111: data <= 9'h000; 
        10'b1001011000: data <= 9'h000; 
        10'b1001011001: data <= 9'h000; 
        10'b1001011010: data <= 9'h000; 
        10'b1001011011: data <= 9'h000; 
        10'b1001011100: data <= 9'h001; 
        10'b1001011101: data <= 9'h000; 
        10'b1001011110: data <= 9'h001; 
        10'b1001011111: data <= 9'h002; 
        10'b1001100000: data <= 9'h001; 
        10'b1001100001: data <= 9'h000; 
        10'b1001100010: data <= 9'h000; 
        10'b1001100011: data <= 9'h1ff; 
        10'b1001100100: data <= 9'h000; 
        10'b1001100101: data <= 9'h000; 
        10'b1001100110: data <= 9'h1ff; 
        10'b1001100111: data <= 9'h000; 
        10'b1001101000: data <= 9'h000; 
        10'b1001101001: data <= 9'h000; 
        10'b1001101010: data <= 9'h000; 
        10'b1001101011: data <= 9'h001; 
        10'b1001101100: data <= 9'h001; 
        10'b1001101101: data <= 9'h001; 
        10'b1001101110: data <= 9'h001; 
        10'b1001101111: data <= 9'h001; 
        10'b1001110000: data <= 9'h000; 
        10'b1001110001: data <= 9'h001; 
        10'b1001110010: data <= 9'h001; 
        10'b1001110011: data <= 9'h001; 
        10'b1001110100: data <= 9'h000; 
        10'b1001110101: data <= 9'h000; 
        10'b1001110110: data <= 9'h000; 
        10'b1001110111: data <= 9'h000; 
        10'b1001111000: data <= 9'h000; 
        10'b1001111001: data <= 9'h000; 
        10'b1001111010: data <= 9'h000; 
        10'b1001111011: data <= 9'h001; 
        10'b1001111100: data <= 9'h001; 
        10'b1001111101: data <= 9'h000; 
        10'b1001111110: data <= 9'h000; 
        10'b1001111111: data <= 9'h000; 
        10'b1010000000: data <= 9'h1ff; 
        10'b1010000001: data <= 9'h1ff; 
        10'b1010000010: data <= 9'h000; 
        10'b1010000011: data <= 9'h000; 
        10'b1010000100: data <= 9'h000; 
        10'b1010000101: data <= 9'h000; 
        10'b1010000110: data <= 9'h000; 
        10'b1010000111: data <= 9'h000; 
        10'b1010001000: data <= 9'h001; 
        10'b1010001001: data <= 9'h002; 
        10'b1010001010: data <= 9'h001; 
        10'b1010001011: data <= 9'h001; 
        10'b1010001100: data <= 9'h000; 
        10'b1010001101: data <= 9'h001; 
        10'b1010001110: data <= 9'h001; 
        10'b1010001111: data <= 9'h000; 
        10'b1010010000: data <= 9'h000; 
        10'b1010010001: data <= 9'h000; 
        10'b1010010010: data <= 9'h000; 
        10'b1010010011: data <= 9'h000; 
        10'b1010010100: data <= 9'h000; 
        10'b1010010101: data <= 9'h001; 
        10'b1010010110: data <= 9'h001; 
        10'b1010010111: data <= 9'h000; 
        10'b1010011000: data <= 9'h1ff; 
        10'b1010011001: data <= 9'h1ff; 
        10'b1010011010: data <= 9'h000; 
        10'b1010011011: data <= 9'h000; 
        10'b1010011100: data <= 9'h000; 
        10'b1010011101: data <= 9'h000; 
        10'b1010011110: data <= 9'h000; 
        10'b1010011111: data <= 9'h000; 
        10'b1010100000: data <= 9'h000; 
        10'b1010100001: data <= 9'h000; 
        10'b1010100010: data <= 9'h000; 
        10'b1010100011: data <= 9'h000; 
        10'b1010100100: data <= 9'h001; 
        10'b1010100101: data <= 9'h001; 
        10'b1010100110: data <= 9'h001; 
        10'b1010100111: data <= 9'h002; 
        10'b1010101000: data <= 9'h002; 
        10'b1010101001: data <= 9'h001; 
        10'b1010101010: data <= 9'h002; 
        10'b1010101011: data <= 9'h002; 
        10'b1010101100: data <= 9'h002; 
        10'b1010101101: data <= 9'h002; 
        10'b1010101110: data <= 9'h001; 
        10'b1010101111: data <= 9'h001; 
        10'b1010110000: data <= 9'h001; 
        10'b1010110001: data <= 9'h000; 
        10'b1010110010: data <= 9'h1ff; 
        10'b1010110011: data <= 9'h1ff; 
        10'b1010110100: data <= 9'h1ff; 
        10'b1010110101: data <= 9'h1ff; 
        10'b1010110110: data <= 9'h1ff; 
        10'b1010110111: data <= 9'h000; 
        10'b1010111000: data <= 9'h000; 
        10'b1010111001: data <= 9'h000; 
        10'b1010111010: data <= 9'h000; 
        10'b1010111011: data <= 9'h000; 
        10'b1010111100: data <= 9'h000; 
        10'b1010111101: data <= 9'h1ff; 
        10'b1010111110: data <= 9'h000; 
        10'b1010111111: data <= 9'h000; 
        10'b1011000000: data <= 9'h000; 
        10'b1011000001: data <= 9'h000; 
        10'b1011000010: data <= 9'h001; 
        10'b1011000011: data <= 9'h000; 
        10'b1011000100: data <= 9'h001; 
        10'b1011000101: data <= 9'h001; 
        10'b1011000110: data <= 9'h002; 
        10'b1011000111: data <= 9'h002; 
        10'b1011001000: data <= 9'h002; 
        10'b1011001001: data <= 9'h002; 
        10'b1011001010: data <= 9'h001; 
        10'b1011001011: data <= 9'h000; 
        10'b1011001100: data <= 9'h000; 
        10'b1011001101: data <= 9'h1ff; 
        10'b1011001110: data <= 9'h1ff; 
        10'b1011001111: data <= 9'h1ff; 
        10'b1011010000: data <= 9'h1ff; 
        10'b1011010001: data <= 9'h000; 
        10'b1011010010: data <= 9'h000; 
        10'b1011010011: data <= 9'h000; 
        10'b1011010100: data <= 9'h000; 
        10'b1011010101: data <= 9'h000; 
        10'b1011010110: data <= 9'h000; 
        10'b1011010111: data <= 9'h000; 
        10'b1011011000: data <= 9'h000; 
        10'b1011011001: data <= 9'h1ff; 
        10'b1011011010: data <= 9'h000; 
        10'b1011011011: data <= 9'h000; 
        10'b1011011100: data <= 9'h000; 
        10'b1011011101: data <= 9'h000; 
        10'b1011011110: data <= 9'h000; 
        10'b1011011111: data <= 9'h000; 
        10'b1011100000: data <= 9'h000; 
        10'b1011100001: data <= 9'h000; 
        10'b1011100010: data <= 9'h000; 
        10'b1011100011: data <= 9'h000; 
        10'b1011100100: data <= 9'h000; 
        10'b1011100101: data <= 9'h000; 
        10'b1011100110: data <= 9'h000; 
        10'b1011100111: data <= 9'h1ff; 
        10'b1011101000: data <= 9'h000; 
        10'b1011101001: data <= 9'h000; 
        10'b1011101010: data <= 9'h000; 
        10'b1011101011: data <= 9'h000; 
        10'b1011101100: data <= 9'h000; 
        10'b1011101101: data <= 9'h000; 
        10'b1011101110: data <= 9'h000; 
        10'b1011101111: data <= 9'h000; 
        10'b1011110000: data <= 9'h000; 
        10'b1011110001: data <= 9'h000; 
        10'b1011110010: data <= 9'h000; 
        10'b1011110011: data <= 9'h000; 
        10'b1011110100: data <= 9'h000; 
        10'b1011110101: data <= 9'h000; 
        10'b1011110110: data <= 9'h000; 
        10'b1011110111: data <= 9'h000; 
        10'b1011111000: data <= 9'h000; 
        10'b1011111001: data <= 9'h000; 
        10'b1011111010: data <= 9'h000; 
        10'b1011111011: data <= 9'h000; 
        10'b1011111100: data <= 9'h000; 
        10'b1011111101: data <= 9'h000; 
        10'b1011111110: data <= 9'h000; 
        10'b1011111111: data <= 9'h000; 
        10'b1100000000: data <= 9'h000; 
        10'b1100000001: data <= 9'h000; 
        10'b1100000010: data <= 9'h000; 
        10'b1100000011: data <= 9'h000; 
        10'b1100000100: data <= 9'h000; 
        10'b1100000101: data <= 9'h000; 
        10'b1100000110: data <= 9'h000; 
        10'b1100000111: data <= 9'h000; 
        10'b1100001000: data <= 9'h000; 
        10'b1100001001: data <= 9'h000; 
        10'b1100001010: data <= 9'h000; 
        10'b1100001011: data <= 9'h000; 
        10'b1100001100: data <= 9'h000; 
        10'b1100001101: data <= 9'h000; 
        10'b1100001110: data <= 9'h000; 
        10'b1100001111: data <= 9'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 4) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 10'h000; 
        10'b0000000001: data <= 10'h3ff; 
        10'b0000000010: data <= 10'h000; 
        10'b0000000011: data <= 10'h000; 
        10'b0000000100: data <= 10'h000; 
        10'b0000000101: data <= 10'h000; 
        10'b0000000110: data <= 10'h000; 
        10'b0000000111: data <= 10'h000; 
        10'b0000001000: data <= 10'h3ff; 
        10'b0000001001: data <= 10'h000; 
        10'b0000001010: data <= 10'h000; 
        10'b0000001011: data <= 10'h3ff; 
        10'b0000001100: data <= 10'h3ff; 
        10'b0000001101: data <= 10'h3ff; 
        10'b0000001110: data <= 10'h3ff; 
        10'b0000001111: data <= 10'h000; 
        10'b0000010000: data <= 10'h000; 
        10'b0000010001: data <= 10'h000; 
        10'b0000010010: data <= 10'h3ff; 
        10'b0000010011: data <= 10'h000; 
        10'b0000010100: data <= 10'h000; 
        10'b0000010101: data <= 10'h000; 
        10'b0000010110: data <= 10'h3ff; 
        10'b0000010111: data <= 10'h000; 
        10'b0000011000: data <= 10'h000; 
        10'b0000011001: data <= 10'h3ff; 
        10'b0000011010: data <= 10'h000; 
        10'b0000011011: data <= 10'h000; 
        10'b0000011100: data <= 10'h3ff; 
        10'b0000011101: data <= 10'h3ff; 
        10'b0000011110: data <= 10'h3ff; 
        10'b0000011111: data <= 10'h000; 
        10'b0000100000: data <= 10'h3ff; 
        10'b0000100001: data <= 10'h000; 
        10'b0000100010: data <= 10'h000; 
        10'b0000100011: data <= 10'h000; 
        10'b0000100100: data <= 10'h3ff; 
        10'b0000100101: data <= 10'h3ff; 
        10'b0000100110: data <= 10'h3ff; 
        10'b0000100111: data <= 10'h000; 
        10'b0000101000: data <= 10'h000; 
        10'b0000101001: data <= 10'h000; 
        10'b0000101010: data <= 10'h3ff; 
        10'b0000101011: data <= 10'h3ff; 
        10'b0000101100: data <= 10'h000; 
        10'b0000101101: data <= 10'h3ff; 
        10'b0000101110: data <= 10'h000; 
        10'b0000101111: data <= 10'h3ff; 
        10'b0000110000: data <= 10'h3ff; 
        10'b0000110001: data <= 10'h3ff; 
        10'b0000110010: data <= 10'h000; 
        10'b0000110011: data <= 10'h000; 
        10'b0000110100: data <= 10'h3ff; 
        10'b0000110101: data <= 10'h000; 
        10'b0000110110: data <= 10'h000; 
        10'b0000110111: data <= 10'h3ff; 
        10'b0000111000: data <= 10'h3ff; 
        10'b0000111001: data <= 10'h000; 
        10'b0000111010: data <= 10'h000; 
        10'b0000111011: data <= 10'h3ff; 
        10'b0000111100: data <= 10'h000; 
        10'b0000111101: data <= 10'h000; 
        10'b0000111110: data <= 10'h3ff; 
        10'b0000111111: data <= 10'h000; 
        10'b0001000000: data <= 10'h000; 
        10'b0001000001: data <= 10'h000; 
        10'b0001000010: data <= 10'h3ff; 
        10'b0001000011: data <= 10'h3ff; 
        10'b0001000100: data <= 10'h3ff; 
        10'b0001000101: data <= 10'h3ff; 
        10'b0001000110: data <= 10'h3ff; 
        10'b0001000111: data <= 10'h3ff; 
        10'b0001001000: data <= 10'h3ff; 
        10'b0001001001: data <= 10'h3ff; 
        10'b0001001010: data <= 10'h000; 
        10'b0001001011: data <= 10'h000; 
        10'b0001001100: data <= 10'h000; 
        10'b0001001101: data <= 10'h3ff; 
        10'b0001001110: data <= 10'h000; 
        10'b0001001111: data <= 10'h000; 
        10'b0001010000: data <= 10'h000; 
        10'b0001010001: data <= 10'h3ff; 
        10'b0001010010: data <= 10'h3ff; 
        10'b0001010011: data <= 10'h000; 
        10'b0001010100: data <= 10'h000; 
        10'b0001010101: data <= 10'h000; 
        10'b0001010110: data <= 10'h000; 
        10'b0001010111: data <= 10'h000; 
        10'b0001011000: data <= 10'h000; 
        10'b0001011001: data <= 10'h000; 
        10'b0001011010: data <= 10'h000; 
        10'b0001011011: data <= 10'h000; 
        10'b0001011100: data <= 10'h000; 
        10'b0001011101: data <= 10'h000; 
        10'b0001011110: data <= 10'h000; 
        10'b0001011111: data <= 10'h001; 
        10'b0001100000: data <= 10'h002; 
        10'b0001100001: data <= 10'h002; 
        10'b0001100010: data <= 10'h002; 
        10'b0001100011: data <= 10'h002; 
        10'b0001100100: data <= 10'h002; 
        10'b0001100101: data <= 10'h002; 
        10'b0001100110: data <= 10'h001; 
        10'b0001100111: data <= 10'h000; 
        10'b0001101000: data <= 10'h000; 
        10'b0001101001: data <= 10'h3fe; 
        10'b0001101010: data <= 10'h3ff; 
        10'b0001101011: data <= 10'h000; 
        10'b0001101100: data <= 10'h000; 
        10'b0001101101: data <= 10'h3ff; 
        10'b0001101110: data <= 10'h000; 
        10'b0001101111: data <= 10'h3ff; 
        10'b0001110000: data <= 10'h000; 
        10'b0001110001: data <= 10'h000; 
        10'b0001110010: data <= 10'h000; 
        10'b0001110011: data <= 10'h000; 
        10'b0001110100: data <= 10'h000; 
        10'b0001110101: data <= 10'h000; 
        10'b0001110110: data <= 10'h001; 
        10'b0001110111: data <= 10'h001; 
        10'b0001111000: data <= 10'h003; 
        10'b0001111001: data <= 10'h003; 
        10'b0001111010: data <= 10'h004; 
        10'b0001111011: data <= 10'h004; 
        10'b0001111100: data <= 10'h005; 
        10'b0001111101: data <= 10'h005; 
        10'b0001111110: data <= 10'h005; 
        10'b0001111111: data <= 10'h003; 
        10'b0010000000: data <= 10'h002; 
        10'b0010000001: data <= 10'h002; 
        10'b0010000010: data <= 10'h003; 
        10'b0010000011: data <= 10'h000; 
        10'b0010000100: data <= 10'h3fe; 
        10'b0010000101: data <= 10'h3fd; 
        10'b0010000110: data <= 10'h3fe; 
        10'b0010000111: data <= 10'h3fe; 
        10'b0010001000: data <= 10'h000; 
        10'b0010001001: data <= 10'h000; 
        10'b0010001010: data <= 10'h3ff; 
        10'b0010001011: data <= 10'h000; 
        10'b0010001100: data <= 10'h3ff; 
        10'b0010001101: data <= 10'h3ff; 
        10'b0010001110: data <= 10'h3ff; 
        10'b0010001111: data <= 10'h3ff; 
        10'b0010010000: data <= 10'h000; 
        10'b0010010001: data <= 10'h001; 
        10'b0010010010: data <= 10'h003; 
        10'b0010010011: data <= 10'h002; 
        10'b0010010100: data <= 10'h002; 
        10'b0010010101: data <= 10'h002; 
        10'b0010010110: data <= 10'h002; 
        10'b0010010111: data <= 10'h003; 
        10'b0010011000: data <= 10'h003; 
        10'b0010011001: data <= 10'h003; 
        10'b0010011010: data <= 10'h001; 
        10'b0010011011: data <= 10'h002; 
        10'b0010011100: data <= 10'h002; 
        10'b0010011101: data <= 10'h000; 
        10'b0010011110: data <= 10'h000; 
        10'b0010011111: data <= 10'h3ff; 
        10'b0010100000: data <= 10'h3fe; 
        10'b0010100001: data <= 10'h3fd; 
        10'b0010100010: data <= 10'h3fc; 
        10'b0010100011: data <= 10'h3fc; 
        10'b0010100100: data <= 10'h3ff; 
        10'b0010100101: data <= 10'h000; 
        10'b0010100110: data <= 10'h3ff; 
        10'b0010100111: data <= 10'h000; 
        10'b0010101000: data <= 10'h3ff; 
        10'b0010101001: data <= 10'h3ff; 
        10'b0010101010: data <= 10'h3ff; 
        10'b0010101011: data <= 10'h000; 
        10'b0010101100: data <= 10'h002; 
        10'b0010101101: data <= 10'h003; 
        10'b0010101110: data <= 10'h003; 
        10'b0010101111: data <= 10'h002; 
        10'b0010110000: data <= 10'h003; 
        10'b0010110001: data <= 10'h002; 
        10'b0010110010: data <= 10'h002; 
        10'b0010110011: data <= 10'h002; 
        10'b0010110100: data <= 10'h003; 
        10'b0010110101: data <= 10'h004; 
        10'b0010110110: data <= 10'h003; 
        10'b0010110111: data <= 10'h001; 
        10'b0010111000: data <= 10'h003; 
        10'b0010111001: data <= 10'h002; 
        10'b0010111010: data <= 10'h002; 
        10'b0010111011: data <= 10'h3ff; 
        10'b0010111100: data <= 10'h001; 
        10'b0010111101: data <= 10'h3ff; 
        10'b0010111110: data <= 10'h3fc; 
        10'b0010111111: data <= 10'h3fc; 
        10'b0011000000: data <= 10'h3fe; 
        10'b0011000001: data <= 10'h000; 
        10'b0011000010: data <= 10'h000; 
        10'b0011000011: data <= 10'h000; 
        10'b0011000100: data <= 10'h000; 
        10'b0011000101: data <= 10'h000; 
        10'b0011000110: data <= 10'h000; 
        10'b0011000111: data <= 10'h002; 
        10'b0011001000: data <= 10'h004; 
        10'b0011001001: data <= 10'h004; 
        10'b0011001010: data <= 10'h003; 
        10'b0011001011: data <= 10'h001; 
        10'b0011001100: data <= 10'h001; 
        10'b0011001101: data <= 10'h002; 
        10'b0011001110: data <= 10'h001; 
        10'b0011001111: data <= 10'h001; 
        10'b0011010000: data <= 10'h002; 
        10'b0011010001: data <= 10'h002; 
        10'b0011010010: data <= 10'h004; 
        10'b0011010011: data <= 10'h002; 
        10'b0011010100: data <= 10'h001; 
        10'b0011010101: data <= 10'h002; 
        10'b0011010110: data <= 10'h002; 
        10'b0011010111: data <= 10'h002; 
        10'b0011011000: data <= 10'h002; 
        10'b0011011001: data <= 10'h000; 
        10'b0011011010: data <= 10'h3fe; 
        10'b0011011011: data <= 10'h3fc; 
        10'b0011011100: data <= 10'h3fd; 
        10'b0011011101: data <= 10'h3ff; 
        10'b0011011110: data <= 10'h3ff; 
        10'b0011011111: data <= 10'h3ff; 
        10'b0011100000: data <= 10'h000; 
        10'b0011100001: data <= 10'h3ff; 
        10'b0011100010: data <= 10'h000; 
        10'b0011100011: data <= 10'h001; 
        10'b0011100100: data <= 10'h003; 
        10'b0011100101: data <= 10'h003; 
        10'b0011100110: data <= 10'h002; 
        10'b0011100111: data <= 10'h001; 
        10'b0011101000: data <= 10'h002; 
        10'b0011101001: data <= 10'h001; 
        10'b0011101010: data <= 10'h002; 
        10'b0011101011: data <= 10'h001; 
        10'b0011101100: data <= 10'h001; 
        10'b0011101101: data <= 10'h001; 
        10'b0011101110: data <= 10'h004; 
        10'b0011101111: data <= 10'h003; 
        10'b0011110000: data <= 10'h001; 
        10'b0011110001: data <= 10'h002; 
        10'b0011110010: data <= 10'h003; 
        10'b0011110011: data <= 10'h002; 
        10'b0011110100: data <= 10'h003; 
        10'b0011110101: data <= 10'h001; 
        10'b0011110110: data <= 10'h3ff; 
        10'b0011110111: data <= 10'h3fc; 
        10'b0011111000: data <= 10'h3fd; 
        10'b0011111001: data <= 10'h3ff; 
        10'b0011111010: data <= 10'h3ff; 
        10'b0011111011: data <= 10'h3ff; 
        10'b0011111100: data <= 10'h000; 
        10'b0011111101: data <= 10'h3ff; 
        10'b0011111110: data <= 10'h000; 
        10'b0011111111: data <= 10'h001; 
        10'b0100000000: data <= 10'h002; 
        10'b0100000001: data <= 10'h002; 
        10'b0100000010: data <= 10'h002; 
        10'b0100000011: data <= 10'h000; 
        10'b0100000100: data <= 10'h000; 
        10'b0100000101: data <= 10'h3fe; 
        10'b0100000110: data <= 10'h3fd; 
        10'b0100000111: data <= 10'h3fa; 
        10'b0100001000: data <= 10'h3fb; 
        10'b0100001001: data <= 10'h3ff; 
        10'b0100001010: data <= 10'h005; 
        10'b0100001011: data <= 10'h007; 
        10'b0100001100: data <= 10'h004; 
        10'b0100001101: data <= 10'h003; 
        10'b0100001110: data <= 10'h003; 
        10'b0100001111: data <= 10'h003; 
        10'b0100010000: data <= 10'h004; 
        10'b0100010001: data <= 10'h002; 
        10'b0100010010: data <= 10'h3ff; 
        10'b0100010011: data <= 10'h3fc; 
        10'b0100010100: data <= 10'h3fe; 
        10'b0100010101: data <= 10'h3ff; 
        10'b0100010110: data <= 10'h3ff; 
        10'b0100010111: data <= 10'h3ff; 
        10'b0100011000: data <= 10'h000; 
        10'b0100011001: data <= 10'h000; 
        10'b0100011010: data <= 10'h000; 
        10'b0100011011: data <= 10'h001; 
        10'b0100011100: data <= 10'h001; 
        10'b0100011101: data <= 10'h000; 
        10'b0100011110: data <= 10'h3ff; 
        10'b0100011111: data <= 10'h3fd; 
        10'b0100100000: data <= 10'h3fb; 
        10'b0100100001: data <= 10'h3f9; 
        10'b0100100010: data <= 10'h3f7; 
        10'b0100100011: data <= 10'h3f7; 
        10'b0100100100: data <= 10'h3f9; 
        10'b0100100101: data <= 10'h3fe; 
        10'b0100100110: data <= 10'h004; 
        10'b0100100111: data <= 10'h005; 
        10'b0100101000: data <= 10'h004; 
        10'b0100101001: data <= 10'h004; 
        10'b0100101010: data <= 10'h002; 
        10'b0100101011: data <= 10'h004; 
        10'b0100101100: data <= 10'h004; 
        10'b0100101101: data <= 10'h001; 
        10'b0100101110: data <= 10'h3ff; 
        10'b0100101111: data <= 10'h3fe; 
        10'b0100110000: data <= 10'h3ff; 
        10'b0100110001: data <= 10'h3ff; 
        10'b0100110010: data <= 10'h000; 
        10'b0100110011: data <= 10'h000; 
        10'b0100110100: data <= 10'h000; 
        10'b0100110101: data <= 10'h000; 
        10'b0100110110: data <= 10'h3ff; 
        10'b0100110111: data <= 10'h001; 
        10'b0100111000: data <= 10'h3ff; 
        10'b0100111001: data <= 10'h3fd; 
        10'b0100111010: data <= 10'h3fc; 
        10'b0100111011: data <= 10'h3fa; 
        10'b0100111100: data <= 10'h3f8; 
        10'b0100111101: data <= 10'h3f9; 
        10'b0100111110: data <= 10'h3fb; 
        10'b0100111111: data <= 10'h3fe; 
        10'b0101000000: data <= 10'h3ff; 
        10'b0101000001: data <= 10'h002; 
        10'b0101000010: data <= 10'h003; 
        10'b0101000011: data <= 10'h003; 
        10'b0101000100: data <= 10'h001; 
        10'b0101000101: data <= 10'h003; 
        10'b0101000110: data <= 10'h003; 
        10'b0101000111: data <= 10'h003; 
        10'b0101001000: data <= 10'h003; 
        10'b0101001001: data <= 10'h000; 
        10'b0101001010: data <= 10'h3ff; 
        10'b0101001011: data <= 10'h3ff; 
        10'b0101001100: data <= 10'h3ff; 
        10'b0101001101: data <= 10'h3ff; 
        10'b0101001110: data <= 10'h3ff; 
        10'b0101001111: data <= 10'h3ff; 
        10'b0101010000: data <= 10'h000; 
        10'b0101010001: data <= 10'h3ff; 
        10'b0101010010: data <= 10'h000; 
        10'b0101010011: data <= 10'h000; 
        10'b0101010100: data <= 10'h3ff; 
        10'b0101010101: data <= 10'h3fd; 
        10'b0101010110: data <= 10'h3fb; 
        10'b0101010111: data <= 10'h3fa; 
        10'b0101011000: data <= 10'h3fa; 
        10'b0101011001: data <= 10'h3fd; 
        10'b0101011010: data <= 10'h000; 
        10'b0101011011: data <= 10'h000; 
        10'b0101011100: data <= 10'h001; 
        10'b0101011101: data <= 10'h002; 
        10'b0101011110: data <= 10'h004; 
        10'b0101011111: data <= 10'h002; 
        10'b0101100000: data <= 10'h002; 
        10'b0101100001: data <= 10'h002; 
        10'b0101100010: data <= 10'h002; 
        10'b0101100011: data <= 10'h000; 
        10'b0101100100: data <= 10'h3fe; 
        10'b0101100101: data <= 10'h3fd; 
        10'b0101100110: data <= 10'h3fd; 
        10'b0101100111: data <= 10'h3fe; 
        10'b0101101000: data <= 10'h000; 
        10'b0101101001: data <= 10'h3ff; 
        10'b0101101010: data <= 10'h000; 
        10'b0101101011: data <= 10'h000; 
        10'b0101101100: data <= 10'h000; 
        10'b0101101101: data <= 10'h3ff; 
        10'b0101101110: data <= 10'h000; 
        10'b0101101111: data <= 10'h000; 
        10'b0101110000: data <= 10'h3ff; 
        10'b0101110001: data <= 10'h3fe; 
        10'b0101110010: data <= 10'h3fc; 
        10'b0101110011: data <= 10'h3fb; 
        10'b0101110100: data <= 10'h3fd; 
        10'b0101110101: data <= 10'h3ff; 
        10'b0101110110: data <= 10'h3ff; 
        10'b0101110111: data <= 10'h3fd; 
        10'b0101111000: data <= 10'h000; 
        10'b0101111001: data <= 10'h004; 
        10'b0101111010: data <= 10'h004; 
        10'b0101111011: data <= 10'h001; 
        10'b0101111100: data <= 10'h002; 
        10'b0101111101: data <= 10'h002; 
        10'b0101111110: data <= 10'h001; 
        10'b0101111111: data <= 10'h3ff; 
        10'b0110000000: data <= 10'h3fc; 
        10'b0110000001: data <= 10'h3fc; 
        10'b0110000010: data <= 10'h3fd; 
        10'b0110000011: data <= 10'h3fe; 
        10'b0110000100: data <= 10'h3ff; 
        10'b0110000101: data <= 10'h000; 
        10'b0110000110: data <= 10'h000; 
        10'b0110000111: data <= 10'h3ff; 
        10'b0110001000: data <= 10'h000; 
        10'b0110001001: data <= 10'h3ff; 
        10'b0110001010: data <= 10'h000; 
        10'b0110001011: data <= 10'h000; 
        10'b0110001100: data <= 10'h000; 
        10'b0110001101: data <= 10'h3fe; 
        10'b0110001110: data <= 10'h3fc; 
        10'b0110001111: data <= 10'h3fd; 
        10'b0110010000: data <= 10'h3fe; 
        10'b0110010001: data <= 10'h000; 
        10'b0110010010: data <= 10'h3fe; 
        10'b0110010011: data <= 10'h3fe; 
        10'b0110010100: data <= 10'h001; 
        10'b0110010101: data <= 10'h002; 
        10'b0110010110: data <= 10'h002; 
        10'b0110010111: data <= 10'h000; 
        10'b0110011000: data <= 10'h3ff; 
        10'b0110011001: data <= 10'h3ff; 
        10'b0110011010: data <= 10'h000; 
        10'b0110011011: data <= 10'h3fe; 
        10'b0110011100: data <= 10'h3fe; 
        10'b0110011101: data <= 10'h3ff; 
        10'b0110011110: data <= 10'h3ff; 
        10'b0110011111: data <= 10'h3ff; 
        10'b0110100000: data <= 10'h3ff; 
        10'b0110100001: data <= 10'h3ff; 
        10'b0110100010: data <= 10'h000; 
        10'b0110100011: data <= 10'h000; 
        10'b0110100100: data <= 10'h000; 
        10'b0110100101: data <= 10'h3ff; 
        10'b0110100110: data <= 10'h000; 
        10'b0110100111: data <= 10'h000; 
        10'b0110101000: data <= 10'h000; 
        10'b0110101001: data <= 10'h3fe; 
        10'b0110101010: data <= 10'h3fd; 
        10'b0110101011: data <= 10'h3fc; 
        10'b0110101100: data <= 10'h3fd; 
        10'b0110101101: data <= 10'h3fe; 
        10'b0110101110: data <= 10'h3fe; 
        10'b0110101111: data <= 10'h3ff; 
        10'b0110110000: data <= 10'h001; 
        10'b0110110001: data <= 10'h003; 
        10'b0110110010: data <= 10'h002; 
        10'b0110110011: data <= 10'h000; 
        10'b0110110100: data <= 10'h3fe; 
        10'b0110110101: data <= 10'h3ff; 
        10'b0110110110: data <= 10'h000; 
        10'b0110110111: data <= 10'h001; 
        10'b0110111000: data <= 10'h002; 
        10'b0110111001: data <= 10'h002; 
        10'b0110111010: data <= 10'h001; 
        10'b0110111011: data <= 10'h000; 
        10'b0110111100: data <= 10'h3ff; 
        10'b0110111101: data <= 10'h000; 
        10'b0110111110: data <= 10'h000; 
        10'b0110111111: data <= 10'h3ff; 
        10'b0111000000: data <= 10'h000; 
        10'b0111000001: data <= 10'h000; 
        10'b0111000010: data <= 10'h001; 
        10'b0111000011: data <= 10'h000; 
        10'b0111000100: data <= 10'h001; 
        10'b0111000101: data <= 10'h3ff; 
        10'b0111000110: data <= 10'h3ff; 
        10'b0111000111: data <= 10'h3fe; 
        10'b0111001000: data <= 10'h3fb; 
        10'b0111001001: data <= 10'h3fb; 
        10'b0111001010: data <= 10'h3fb; 
        10'b0111001011: data <= 10'h3ff; 
        10'b0111001100: data <= 10'h001; 
        10'b0111001101: data <= 10'h004; 
        10'b0111001110: data <= 10'h000; 
        10'b0111001111: data <= 10'h3fd; 
        10'b0111010000: data <= 10'h3fd; 
        10'b0111010001: data <= 10'h3ff; 
        10'b0111010010: data <= 10'h001; 
        10'b0111010011: data <= 10'h003; 
        10'b0111010100: data <= 10'h002; 
        10'b0111010101: data <= 10'h003; 
        10'b0111010110: data <= 10'h003; 
        10'b0111010111: data <= 10'h001; 
        10'b0111011000: data <= 10'h000; 
        10'b0111011001: data <= 10'h000; 
        10'b0111011010: data <= 10'h000; 
        10'b0111011011: data <= 10'h000; 
        10'b0111011100: data <= 10'h000; 
        10'b0111011101: data <= 10'h000; 
        10'b0111011110: data <= 10'h000; 
        10'b0111011111: data <= 10'h002; 
        10'b0111100000: data <= 10'h001; 
        10'b0111100001: data <= 10'h000; 
        10'b0111100010: data <= 10'h3ff; 
        10'b0111100011: data <= 10'h3fd; 
        10'b0111100100: data <= 10'h3fa; 
        10'b0111100101: data <= 10'h3f7; 
        10'b0111100110: data <= 10'h3f5; 
        10'b0111100111: data <= 10'h3f6; 
        10'b0111101000: data <= 10'h3f8; 
        10'b0111101001: data <= 10'h3fc; 
        10'b0111101010: data <= 10'h3fc; 
        10'b0111101011: data <= 10'h3fc; 
        10'b0111101100: data <= 10'h000; 
        10'b0111101101: data <= 10'h001; 
        10'b0111101110: data <= 10'h002; 
        10'b0111101111: data <= 10'h003; 
        10'b0111110000: data <= 10'h001; 
        10'b0111110001: data <= 10'h004; 
        10'b0111110010: data <= 10'h004; 
        10'b0111110011: data <= 10'h001; 
        10'b0111110100: data <= 10'h3ff; 
        10'b0111110101: data <= 10'h3ff; 
        10'b0111110110: data <= 10'h3ff; 
        10'b0111110111: data <= 10'h3ff; 
        10'b0111111000: data <= 10'h000; 
        10'b0111111001: data <= 10'h000; 
        10'b0111111010: data <= 10'h000; 
        10'b0111111011: data <= 10'h003; 
        10'b0111111100: data <= 10'h002; 
        10'b0111111101: data <= 10'h001; 
        10'b0111111110: data <= 10'h001; 
        10'b0111111111: data <= 10'h3ff; 
        10'b1000000000: data <= 10'h3fe; 
        10'b1000000001: data <= 10'h3fa; 
        10'b1000000010: data <= 10'h3f6; 
        10'b1000000011: data <= 10'h3f7; 
        10'b1000000100: data <= 10'h3f5; 
        10'b1000000101: data <= 10'h3f7; 
        10'b1000000110: data <= 10'h3fa; 
        10'b1000000111: data <= 10'h3ff; 
        10'b1000001000: data <= 10'h002; 
        10'b1000001001: data <= 10'h003; 
        10'b1000001010: data <= 10'h003; 
        10'b1000001011: data <= 10'h003; 
        10'b1000001100: data <= 10'h002; 
        10'b1000001101: data <= 10'h005; 
        10'b1000001110: data <= 10'h004; 
        10'b1000001111: data <= 10'h002; 
        10'b1000010000: data <= 10'h3ff; 
        10'b1000010001: data <= 10'h3ff; 
        10'b1000010010: data <= 10'h3ff; 
        10'b1000010011: data <= 10'h000; 
        10'b1000010100: data <= 10'h000; 
        10'b1000010101: data <= 10'h3ff; 
        10'b1000010110: data <= 10'h000; 
        10'b1000010111: data <= 10'h003; 
        10'b1000011000: data <= 10'h003; 
        10'b1000011001: data <= 10'h004; 
        10'b1000011010: data <= 10'h003; 
        10'b1000011011: data <= 10'h001; 
        10'b1000011100: data <= 10'h000; 
        10'b1000011101: data <= 10'h3ff; 
        10'b1000011110: data <= 10'h3ff; 
        10'b1000011111: data <= 10'h3fd; 
        10'b1000100000: data <= 10'h3fc; 
        10'b1000100001: data <= 10'h3fb; 
        10'b1000100010: data <= 10'h3fd; 
        10'b1000100011: data <= 10'h001; 
        10'b1000100100: data <= 10'h003; 
        10'b1000100101: data <= 10'h004; 
        10'b1000100110: data <= 10'h004; 
        10'b1000100111: data <= 10'h004; 
        10'b1000101000: data <= 10'h003; 
        10'b1000101001: data <= 10'h004; 
        10'b1000101010: data <= 10'h002; 
        10'b1000101011: data <= 10'h000; 
        10'b1000101100: data <= 10'h3ff; 
        10'b1000101101: data <= 10'h000; 
        10'b1000101110: data <= 10'h000; 
        10'b1000101111: data <= 10'h000; 
        10'b1000110000: data <= 10'h000; 
        10'b1000110001: data <= 10'h3ff; 
        10'b1000110010: data <= 10'h001; 
        10'b1000110011: data <= 10'h003; 
        10'b1000110100: data <= 10'h004; 
        10'b1000110101: data <= 10'h005; 
        10'b1000110110: data <= 10'h005; 
        10'b1000110111: data <= 10'h002; 
        10'b1000111000: data <= 10'h003; 
        10'b1000111001: data <= 10'h003; 
        10'b1000111010: data <= 10'h001; 
        10'b1000111011: data <= 10'h000; 
        10'b1000111100: data <= 10'h3ff; 
        10'b1000111101: data <= 10'h3fe; 
        10'b1000111110: data <= 10'h001; 
        10'b1000111111: data <= 10'h001; 
        10'b1001000000: data <= 10'h002; 
        10'b1001000001: data <= 10'h003; 
        10'b1001000010: data <= 10'h003; 
        10'b1001000011: data <= 10'h002; 
        10'b1001000100: data <= 10'h004; 
        10'b1001000101: data <= 10'h002; 
        10'b1001000110: data <= 10'h000; 
        10'b1001000111: data <= 10'h3ff; 
        10'b1001001000: data <= 10'h3ff; 
        10'b1001001001: data <= 10'h000; 
        10'b1001001010: data <= 10'h000; 
        10'b1001001011: data <= 10'h000; 
        10'b1001001100: data <= 10'h3ff; 
        10'b1001001101: data <= 10'h000; 
        10'b1001001110: data <= 10'h000; 
        10'b1001001111: data <= 10'h002; 
        10'b1001010000: data <= 10'h004; 
        10'b1001010001: data <= 10'h004; 
        10'b1001010010: data <= 10'h004; 
        10'b1001010011: data <= 10'h002; 
        10'b1001010100: data <= 10'h002; 
        10'b1001010101: data <= 10'h001; 
        10'b1001010110: data <= 10'h000; 
        10'b1001010111: data <= 10'h3ff; 
        10'b1001011000: data <= 10'h000; 
        10'b1001011001: data <= 10'h000; 
        10'b1001011010: data <= 10'h000; 
        10'b1001011011: data <= 10'h000; 
        10'b1001011100: data <= 10'h001; 
        10'b1001011101: data <= 10'h000; 
        10'b1001011110: data <= 10'h002; 
        10'b1001011111: data <= 10'h003; 
        10'b1001100000: data <= 10'h002; 
        10'b1001100001: data <= 10'h001; 
        10'b1001100010: data <= 10'h3ff; 
        10'b1001100011: data <= 10'h3fe; 
        10'b1001100100: data <= 10'h3ff; 
        10'b1001100101: data <= 10'h3ff; 
        10'b1001100110: data <= 10'h3ff; 
        10'b1001100111: data <= 10'h3ff; 
        10'b1001101000: data <= 10'h000; 
        10'b1001101001: data <= 10'h000; 
        10'b1001101010: data <= 10'h000; 
        10'b1001101011: data <= 10'h001; 
        10'b1001101100: data <= 10'h002; 
        10'b1001101101: data <= 10'h003; 
        10'b1001101110: data <= 10'h003; 
        10'b1001101111: data <= 10'h001; 
        10'b1001110000: data <= 10'h000; 
        10'b1001110001: data <= 10'h001; 
        10'b1001110010: data <= 10'h001; 
        10'b1001110011: data <= 10'h002; 
        10'b1001110100: data <= 10'h000; 
        10'b1001110101: data <= 10'h3ff; 
        10'b1001110110: data <= 10'h3ff; 
        10'b1001110111: data <= 10'h3ff; 
        10'b1001111000: data <= 10'h001; 
        10'b1001111001: data <= 10'h000; 
        10'b1001111010: data <= 10'h000; 
        10'b1001111011: data <= 10'h002; 
        10'b1001111100: data <= 10'h001; 
        10'b1001111101: data <= 10'h000; 
        10'b1001111110: data <= 10'h000; 
        10'b1001111111: data <= 10'h3ff; 
        10'b1010000000: data <= 10'h3ff; 
        10'b1010000001: data <= 10'h3ff; 
        10'b1010000010: data <= 10'h000; 
        10'b1010000011: data <= 10'h000; 
        10'b1010000100: data <= 10'h000; 
        10'b1010000101: data <= 10'h3ff; 
        10'b1010000110: data <= 10'h3ff; 
        10'b1010000111: data <= 10'h001; 
        10'b1010001000: data <= 10'h002; 
        10'b1010001001: data <= 10'h003; 
        10'b1010001010: data <= 10'h003; 
        10'b1010001011: data <= 10'h003; 
        10'b1010001100: data <= 10'h001; 
        10'b1010001101: data <= 10'h002; 
        10'b1010001110: data <= 10'h001; 
        10'b1010001111: data <= 10'h000; 
        10'b1010010000: data <= 10'h3ff; 
        10'b1010010001: data <= 10'h000; 
        10'b1010010010: data <= 10'h000; 
        10'b1010010011: data <= 10'h001; 
        10'b1010010100: data <= 10'h001; 
        10'b1010010101: data <= 10'h001; 
        10'b1010010110: data <= 10'h002; 
        10'b1010010111: data <= 10'h000; 
        10'b1010011000: data <= 10'h3ff; 
        10'b1010011001: data <= 10'h3ff; 
        10'b1010011010: data <= 10'h3ff; 
        10'b1010011011: data <= 10'h3ff; 
        10'b1010011100: data <= 10'h000; 
        10'b1010011101: data <= 10'h000; 
        10'b1010011110: data <= 10'h3ff; 
        10'b1010011111: data <= 10'h3ff; 
        10'b1010100000: data <= 10'h3ff; 
        10'b1010100001: data <= 10'h000; 
        10'b1010100010: data <= 10'h000; 
        10'b1010100011: data <= 10'h000; 
        10'b1010100100: data <= 10'h001; 
        10'b1010100101: data <= 10'h002; 
        10'b1010100110: data <= 10'h003; 
        10'b1010100111: data <= 10'h003; 
        10'b1010101000: data <= 10'h003; 
        10'b1010101001: data <= 10'h003; 
        10'b1010101010: data <= 10'h004; 
        10'b1010101011: data <= 10'h004; 
        10'b1010101100: data <= 10'h004; 
        10'b1010101101: data <= 10'h003; 
        10'b1010101110: data <= 10'h003; 
        10'b1010101111: data <= 10'h002; 
        10'b1010110000: data <= 10'h002; 
        10'b1010110001: data <= 10'h000; 
        10'b1010110010: data <= 10'h3fe; 
        10'b1010110011: data <= 10'h3fe; 
        10'b1010110100: data <= 10'h3fe; 
        10'b1010110101: data <= 10'h3ff; 
        10'b1010110110: data <= 10'h3ff; 
        10'b1010110111: data <= 10'h000; 
        10'b1010111000: data <= 10'h3ff; 
        10'b1010111001: data <= 10'h000; 
        10'b1010111010: data <= 10'h3ff; 
        10'b1010111011: data <= 10'h000; 
        10'b1010111100: data <= 10'h000; 
        10'b1010111101: data <= 10'h3ff; 
        10'b1010111110: data <= 10'h000; 
        10'b1010111111: data <= 10'h000; 
        10'b1011000000: data <= 10'h000; 
        10'b1011000001: data <= 10'h001; 
        10'b1011000010: data <= 10'h001; 
        10'b1011000011: data <= 10'h001; 
        10'b1011000100: data <= 10'h002; 
        10'b1011000101: data <= 10'h002; 
        10'b1011000110: data <= 10'h003; 
        10'b1011000111: data <= 10'h004; 
        10'b1011001000: data <= 10'h004; 
        10'b1011001001: data <= 10'h003; 
        10'b1011001010: data <= 10'h002; 
        10'b1011001011: data <= 10'h001; 
        10'b1011001100: data <= 10'h000; 
        10'b1011001101: data <= 10'h3fe; 
        10'b1011001110: data <= 10'h3fe; 
        10'b1011001111: data <= 10'h3ff; 
        10'b1011010000: data <= 10'h3ff; 
        10'b1011010001: data <= 10'h3ff; 
        10'b1011010010: data <= 10'h3ff; 
        10'b1011010011: data <= 10'h000; 
        10'b1011010100: data <= 10'h3ff; 
        10'b1011010101: data <= 10'h000; 
        10'b1011010110: data <= 10'h3ff; 
        10'b1011010111: data <= 10'h000; 
        10'b1011011000: data <= 10'h3ff; 
        10'b1011011001: data <= 10'h3ff; 
        10'b1011011010: data <= 10'h3ff; 
        10'b1011011011: data <= 10'h000; 
        10'b1011011100: data <= 10'h000; 
        10'b1011011101: data <= 10'h3ff; 
        10'b1011011110: data <= 10'h3ff; 
        10'b1011011111: data <= 10'h000; 
        10'b1011100000: data <= 10'h000; 
        10'b1011100001: data <= 10'h000; 
        10'b1011100010: data <= 10'h000; 
        10'b1011100011: data <= 10'h000; 
        10'b1011100100: data <= 10'h3ff; 
        10'b1011100101: data <= 10'h000; 
        10'b1011100110: data <= 10'h3ff; 
        10'b1011100111: data <= 10'h3ff; 
        10'b1011101000: data <= 10'h3ff; 
        10'b1011101001: data <= 10'h000; 
        10'b1011101010: data <= 10'h000; 
        10'b1011101011: data <= 10'h000; 
        10'b1011101100: data <= 10'h3ff; 
        10'b1011101101: data <= 10'h3ff; 
        10'b1011101110: data <= 10'h000; 
        10'b1011101111: data <= 10'h3ff; 
        10'b1011110000: data <= 10'h000; 
        10'b1011110001: data <= 10'h3ff; 
        10'b1011110010: data <= 10'h000; 
        10'b1011110011: data <= 10'h000; 
        10'b1011110100: data <= 10'h000; 
        10'b1011110101: data <= 10'h3ff; 
        10'b1011110110: data <= 10'h000; 
        10'b1011110111: data <= 10'h3ff; 
        10'b1011111000: data <= 10'h000; 
        10'b1011111001: data <= 10'h000; 
        10'b1011111010: data <= 10'h000; 
        10'b1011111011: data <= 10'h000; 
        10'b1011111100: data <= 10'h000; 
        10'b1011111101: data <= 10'h3ff; 
        10'b1011111110: data <= 10'h3ff; 
        10'b1011111111: data <= 10'h000; 
        10'b1100000000: data <= 10'h3ff; 
        10'b1100000001: data <= 10'h000; 
        10'b1100000010: data <= 10'h3ff; 
        10'b1100000011: data <= 10'h000; 
        10'b1100000100: data <= 10'h3ff; 
        10'b1100000101: data <= 10'h000; 
        10'b1100000110: data <= 10'h3ff; 
        10'b1100000111: data <= 10'h3ff; 
        10'b1100001000: data <= 10'h000; 
        10'b1100001001: data <= 10'h000; 
        10'b1100001010: data <= 10'h3ff; 
        10'b1100001011: data <= 10'h000; 
        10'b1100001100: data <= 10'h3ff; 
        10'b1100001101: data <= 10'h3ff; 
        10'b1100001110: data <= 10'h000; 
        10'b1100001111: data <= 10'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 5) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 11'h7ff; 
        10'b0000000001: data <= 11'h7fe; 
        10'b0000000010: data <= 11'h000; 
        10'b0000000011: data <= 11'h000; 
        10'b0000000100: data <= 11'h000; 
        10'b0000000101: data <= 11'h000; 
        10'b0000000110: data <= 11'h7ff; 
        10'b0000000111: data <= 11'h000; 
        10'b0000001000: data <= 11'h7ff; 
        10'b0000001001: data <= 11'h000; 
        10'b0000001010: data <= 11'h000; 
        10'b0000001011: data <= 11'h7ff; 
        10'b0000001100: data <= 11'h7ff; 
        10'b0000001101: data <= 11'h7ff; 
        10'b0000001110: data <= 11'h7ff; 
        10'b0000001111: data <= 11'h7ff; 
        10'b0000010000: data <= 11'h000; 
        10'b0000010001: data <= 11'h000; 
        10'b0000010010: data <= 11'h7fe; 
        10'b0000010011: data <= 11'h000; 
        10'b0000010100: data <= 11'h7ff; 
        10'b0000010101: data <= 11'h000; 
        10'b0000010110: data <= 11'h7fe; 
        10'b0000010111: data <= 11'h000; 
        10'b0000011000: data <= 11'h000; 
        10'b0000011001: data <= 11'h7fe; 
        10'b0000011010: data <= 11'h7ff; 
        10'b0000011011: data <= 11'h000; 
        10'b0000011100: data <= 11'h7fe; 
        10'b0000011101: data <= 11'h7ff; 
        10'b0000011110: data <= 11'h7fe; 
        10'b0000011111: data <= 11'h7ff; 
        10'b0000100000: data <= 11'h7fe; 
        10'b0000100001: data <= 11'h7ff; 
        10'b0000100010: data <= 11'h000; 
        10'b0000100011: data <= 11'h000; 
        10'b0000100100: data <= 11'h7fe; 
        10'b0000100101: data <= 11'h7fe; 
        10'b0000100110: data <= 11'h7fe; 
        10'b0000100111: data <= 11'h7ff; 
        10'b0000101000: data <= 11'h000; 
        10'b0000101001: data <= 11'h7ff; 
        10'b0000101010: data <= 11'h7ff; 
        10'b0000101011: data <= 11'h7ff; 
        10'b0000101100: data <= 11'h000; 
        10'b0000101101: data <= 11'h7fe; 
        10'b0000101110: data <= 11'h000; 
        10'b0000101111: data <= 11'h7ff; 
        10'b0000110000: data <= 11'h7ff; 
        10'b0000110001: data <= 11'h7fe; 
        10'b0000110010: data <= 11'h7ff; 
        10'b0000110011: data <= 11'h000; 
        10'b0000110100: data <= 11'h7fe; 
        10'b0000110101: data <= 11'h000; 
        10'b0000110110: data <= 11'h7ff; 
        10'b0000110111: data <= 11'h7fe; 
        10'b0000111000: data <= 11'h7ff; 
        10'b0000111001: data <= 11'h7ff; 
        10'b0000111010: data <= 11'h7ff; 
        10'b0000111011: data <= 11'h7fe; 
        10'b0000111100: data <= 11'h000; 
        10'b0000111101: data <= 11'h000; 
        10'b0000111110: data <= 11'h7ff; 
        10'b0000111111: data <= 11'h000; 
        10'b0001000000: data <= 11'h000; 
        10'b0001000001: data <= 11'h7ff; 
        10'b0001000010: data <= 11'h7fe; 
        10'b0001000011: data <= 11'h7fe; 
        10'b0001000100: data <= 11'h7fe; 
        10'b0001000101: data <= 11'h7fe; 
        10'b0001000110: data <= 11'h7ff; 
        10'b0001000111: data <= 11'h7ff; 
        10'b0001001000: data <= 11'h7ff; 
        10'b0001001001: data <= 11'h7ff; 
        10'b0001001010: data <= 11'h000; 
        10'b0001001011: data <= 11'h000; 
        10'b0001001100: data <= 11'h7ff; 
        10'b0001001101: data <= 11'h7fe; 
        10'b0001001110: data <= 11'h000; 
        10'b0001001111: data <= 11'h000; 
        10'b0001010000: data <= 11'h000; 
        10'b0001010001: data <= 11'h7ff; 
        10'b0001010010: data <= 11'h7fe; 
        10'b0001010011: data <= 11'h7ff; 
        10'b0001010100: data <= 11'h000; 
        10'b0001010101: data <= 11'h000; 
        10'b0001010110: data <= 11'h7ff; 
        10'b0001010111: data <= 11'h000; 
        10'b0001011000: data <= 11'h000; 
        10'b0001011001: data <= 11'h000; 
        10'b0001011010: data <= 11'h7ff; 
        10'b0001011011: data <= 11'h000; 
        10'b0001011100: data <= 11'h000; 
        10'b0001011101: data <= 11'h7ff; 
        10'b0001011110: data <= 11'h001; 
        10'b0001011111: data <= 11'h002; 
        10'b0001100000: data <= 11'h005; 
        10'b0001100001: data <= 11'h004; 
        10'b0001100010: data <= 11'h004; 
        10'b0001100011: data <= 11'h005; 
        10'b0001100100: data <= 11'h003; 
        10'b0001100101: data <= 11'h004; 
        10'b0001100110: data <= 11'h003; 
        10'b0001100111: data <= 11'h000; 
        10'b0001101000: data <= 11'h000; 
        10'b0001101001: data <= 11'h7fd; 
        10'b0001101010: data <= 11'h7fe; 
        10'b0001101011: data <= 11'h000; 
        10'b0001101100: data <= 11'h000; 
        10'b0001101101: data <= 11'h7ff; 
        10'b0001101110: data <= 11'h7ff; 
        10'b0001101111: data <= 11'h7ff; 
        10'b0001110000: data <= 11'h7ff; 
        10'b0001110001: data <= 11'h000; 
        10'b0001110010: data <= 11'h7ff; 
        10'b0001110011: data <= 11'h000; 
        10'b0001110100: data <= 11'h001; 
        10'b0001110101: data <= 11'h000; 
        10'b0001110110: data <= 11'h003; 
        10'b0001110111: data <= 11'h002; 
        10'b0001111000: data <= 11'h007; 
        10'b0001111001: data <= 11'h006; 
        10'b0001111010: data <= 11'h007; 
        10'b0001111011: data <= 11'h008; 
        10'b0001111100: data <= 11'h00a; 
        10'b0001111101: data <= 11'h00b; 
        10'b0001111110: data <= 11'h009; 
        10'b0001111111: data <= 11'h007; 
        10'b0010000000: data <= 11'h004; 
        10'b0010000001: data <= 11'h003; 
        10'b0010000010: data <= 11'h005; 
        10'b0010000011: data <= 11'h001; 
        10'b0010000100: data <= 11'h7fc; 
        10'b0010000101: data <= 11'h7fb; 
        10'b0010000110: data <= 11'h7fb; 
        10'b0010000111: data <= 11'h7fb; 
        10'b0010001000: data <= 11'h7ff; 
        10'b0010001001: data <= 11'h7ff; 
        10'b0010001010: data <= 11'h7ff; 
        10'b0010001011: data <= 11'h000; 
        10'b0010001100: data <= 11'h7fe; 
        10'b0010001101: data <= 11'h7fe; 
        10'b0010001110: data <= 11'h7ff; 
        10'b0010001111: data <= 11'h7ff; 
        10'b0010010000: data <= 11'h000; 
        10'b0010010001: data <= 11'h003; 
        10'b0010010010: data <= 11'h005; 
        10'b0010010011: data <= 11'h004; 
        10'b0010010100: data <= 11'h005; 
        10'b0010010101: data <= 11'h004; 
        10'b0010010110: data <= 11'h004; 
        10'b0010010111: data <= 11'h005; 
        10'b0010011000: data <= 11'h005; 
        10'b0010011001: data <= 11'h006; 
        10'b0010011010: data <= 11'h001; 
        10'b0010011011: data <= 11'h004; 
        10'b0010011100: data <= 11'h005; 
        10'b0010011101: data <= 11'h000; 
        10'b0010011110: data <= 11'h000; 
        10'b0010011111: data <= 11'h7fe; 
        10'b0010100000: data <= 11'h7fd; 
        10'b0010100001: data <= 11'h7f9; 
        10'b0010100010: data <= 11'h7f8; 
        10'b0010100011: data <= 11'h7f9; 
        10'b0010100100: data <= 11'h7fe; 
        10'b0010100101: data <= 11'h000; 
        10'b0010100110: data <= 11'h7ff; 
        10'b0010100111: data <= 11'h7ff; 
        10'b0010101000: data <= 11'h7fe; 
        10'b0010101001: data <= 11'h7ff; 
        10'b0010101010: data <= 11'h7ff; 
        10'b0010101011: data <= 11'h001; 
        10'b0010101100: data <= 11'h004; 
        10'b0010101101: data <= 11'h007; 
        10'b0010101110: data <= 11'h005; 
        10'b0010101111: data <= 11'h004; 
        10'b0010110000: data <= 11'h006; 
        10'b0010110001: data <= 11'h005; 
        10'b0010110010: data <= 11'h004; 
        10'b0010110011: data <= 11'h004; 
        10'b0010110100: data <= 11'h006; 
        10'b0010110101: data <= 11'h008; 
        10'b0010110110: data <= 11'h006; 
        10'b0010110111: data <= 11'h002; 
        10'b0010111000: data <= 11'h005; 
        10'b0010111001: data <= 11'h005; 
        10'b0010111010: data <= 11'h005; 
        10'b0010111011: data <= 11'h7fe; 
        10'b0010111100: data <= 11'h002; 
        10'b0010111101: data <= 11'h7fe; 
        10'b0010111110: data <= 11'h7f9; 
        10'b0010111111: data <= 11'h7f9; 
        10'b0011000000: data <= 11'h7fc; 
        10'b0011000001: data <= 11'h7ff; 
        10'b0011000010: data <= 11'h000; 
        10'b0011000011: data <= 11'h7ff; 
        10'b0011000100: data <= 11'h000; 
        10'b0011000101: data <= 11'h000; 
        10'b0011000110: data <= 11'h000; 
        10'b0011000111: data <= 11'h003; 
        10'b0011001000: data <= 11'h008; 
        10'b0011001001: data <= 11'h008; 
        10'b0011001010: data <= 11'h006; 
        10'b0011001011: data <= 11'h002; 
        10'b0011001100: data <= 11'h002; 
        10'b0011001101: data <= 11'h004; 
        10'b0011001110: data <= 11'h001; 
        10'b0011001111: data <= 11'h002; 
        10'b0011010000: data <= 11'h005; 
        10'b0011010001: data <= 11'h005; 
        10'b0011010010: data <= 11'h007; 
        10'b0011010011: data <= 11'h004; 
        10'b0011010100: data <= 11'h001; 
        10'b0011010101: data <= 11'h004; 
        10'b0011010110: data <= 11'h003; 
        10'b0011010111: data <= 11'h003; 
        10'b0011011000: data <= 11'h003; 
        10'b0011011001: data <= 11'h000; 
        10'b0011011010: data <= 11'h7fd; 
        10'b0011011011: data <= 11'h7f8; 
        10'b0011011100: data <= 11'h7fa; 
        10'b0011011101: data <= 11'h7fe; 
        10'b0011011110: data <= 11'h7fe; 
        10'b0011011111: data <= 11'h7ff; 
        10'b0011100000: data <= 11'h7ff; 
        10'b0011100001: data <= 11'h7ff; 
        10'b0011100010: data <= 11'h000; 
        10'b0011100011: data <= 11'h003; 
        10'b0011100100: data <= 11'h007; 
        10'b0011100101: data <= 11'h006; 
        10'b0011100110: data <= 11'h005; 
        10'b0011100111: data <= 11'h002; 
        10'b0011101000: data <= 11'h003; 
        10'b0011101001: data <= 11'h002; 
        10'b0011101010: data <= 11'h004; 
        10'b0011101011: data <= 11'h001; 
        10'b0011101100: data <= 11'h001; 
        10'b0011101101: data <= 11'h002; 
        10'b0011101110: data <= 11'h008; 
        10'b0011101111: data <= 11'h007; 
        10'b0011110000: data <= 11'h002; 
        10'b0011110001: data <= 11'h004; 
        10'b0011110010: data <= 11'h005; 
        10'b0011110011: data <= 11'h004; 
        10'b0011110100: data <= 11'h005; 
        10'b0011110101: data <= 11'h003; 
        10'b0011110110: data <= 11'h7ff; 
        10'b0011110111: data <= 11'h7f9; 
        10'b0011111000: data <= 11'h7fa; 
        10'b0011111001: data <= 11'h7fe; 
        10'b0011111010: data <= 11'h7fe; 
        10'b0011111011: data <= 11'h7ff; 
        10'b0011111100: data <= 11'h7ff; 
        10'b0011111101: data <= 11'h7fe; 
        10'b0011111110: data <= 11'h7ff; 
        10'b0011111111: data <= 11'h001; 
        10'b0100000000: data <= 11'h003; 
        10'b0100000001: data <= 11'h005; 
        10'b0100000010: data <= 11'h004; 
        10'b0100000011: data <= 11'h001; 
        10'b0100000100: data <= 11'h000; 
        10'b0100000101: data <= 11'h7fc; 
        10'b0100000110: data <= 11'h7f9; 
        10'b0100000111: data <= 11'h7f4; 
        10'b0100001000: data <= 11'h7f6; 
        10'b0100001001: data <= 11'h7ff; 
        10'b0100001010: data <= 11'h00a; 
        10'b0100001011: data <= 11'h00f; 
        10'b0100001100: data <= 11'h009; 
        10'b0100001101: data <= 11'h005; 
        10'b0100001110: data <= 11'h005; 
        10'b0100001111: data <= 11'h005; 
        10'b0100010000: data <= 11'h008; 
        10'b0100010001: data <= 11'h005; 
        10'b0100010010: data <= 11'h7ff; 
        10'b0100010011: data <= 11'h7f9; 
        10'b0100010100: data <= 11'h7fc; 
        10'b0100010101: data <= 11'h7fe; 
        10'b0100010110: data <= 11'h7fe; 
        10'b0100010111: data <= 11'h7ff; 
        10'b0100011000: data <= 11'h000; 
        10'b0100011001: data <= 11'h000; 
        10'b0100011010: data <= 11'h000; 
        10'b0100011011: data <= 11'h002; 
        10'b0100011100: data <= 11'h002; 
        10'b0100011101: data <= 11'h001; 
        10'b0100011110: data <= 11'h7fe; 
        10'b0100011111: data <= 11'h7fb; 
        10'b0100100000: data <= 11'h7f6; 
        10'b0100100001: data <= 11'h7f2; 
        10'b0100100010: data <= 11'h7ee; 
        10'b0100100011: data <= 11'h7ee; 
        10'b0100100100: data <= 11'h7f3; 
        10'b0100100101: data <= 11'h7fd; 
        10'b0100100110: data <= 11'h008; 
        10'b0100100111: data <= 11'h009; 
        10'b0100101000: data <= 11'h008; 
        10'b0100101001: data <= 11'h007; 
        10'b0100101010: data <= 11'h004; 
        10'b0100101011: data <= 11'h008; 
        10'b0100101100: data <= 11'h007; 
        10'b0100101101: data <= 11'h003; 
        10'b0100101110: data <= 11'h7fd; 
        10'b0100101111: data <= 11'h7fb; 
        10'b0100110000: data <= 11'h7fe; 
        10'b0100110001: data <= 11'h7fe; 
        10'b0100110010: data <= 11'h7ff; 
        10'b0100110011: data <= 11'h000; 
        10'b0100110100: data <= 11'h000; 
        10'b0100110101: data <= 11'h000; 
        10'b0100110110: data <= 11'h7fe; 
        10'b0100110111: data <= 11'h002; 
        10'b0100111000: data <= 11'h7ff; 
        10'b0100111001: data <= 11'h7fa; 
        10'b0100111010: data <= 11'h7f8; 
        10'b0100111011: data <= 11'h7f4; 
        10'b0100111100: data <= 11'h7f1; 
        10'b0100111101: data <= 11'h7f3; 
        10'b0100111110: data <= 11'h7f6; 
        10'b0100111111: data <= 11'h7fb; 
        10'b0101000000: data <= 11'h7fd; 
        10'b0101000001: data <= 11'h003; 
        10'b0101000010: data <= 11'h005; 
        10'b0101000011: data <= 11'h005; 
        10'b0101000100: data <= 11'h002; 
        10'b0101000101: data <= 11'h005; 
        10'b0101000110: data <= 11'h007; 
        10'b0101000111: data <= 11'h007; 
        10'b0101001000: data <= 11'h006; 
        10'b0101001001: data <= 11'h000; 
        10'b0101001010: data <= 11'h7fd; 
        10'b0101001011: data <= 11'h7fe; 
        10'b0101001100: data <= 11'h7fe; 
        10'b0101001101: data <= 11'h7ff; 
        10'b0101001110: data <= 11'h7fe; 
        10'b0101001111: data <= 11'h7fe; 
        10'b0101010000: data <= 11'h000; 
        10'b0101010001: data <= 11'h7ff; 
        10'b0101010010: data <= 11'h000; 
        10'b0101010011: data <= 11'h000; 
        10'b0101010100: data <= 11'h7fe; 
        10'b0101010101: data <= 11'h7fa; 
        10'b0101010110: data <= 11'h7f6; 
        10'b0101010111: data <= 11'h7f4; 
        10'b0101011000: data <= 11'h7f5; 
        10'b0101011001: data <= 11'h7fa; 
        10'b0101011010: data <= 11'h000; 
        10'b0101011011: data <= 11'h001; 
        10'b0101011100: data <= 11'h002; 
        10'b0101011101: data <= 11'h004; 
        10'b0101011110: data <= 11'h009; 
        10'b0101011111: data <= 11'h005; 
        10'b0101100000: data <= 11'h003; 
        10'b0101100001: data <= 11'h004; 
        10'b0101100010: data <= 11'h004; 
        10'b0101100011: data <= 11'h000; 
        10'b0101100100: data <= 11'h7fb; 
        10'b0101100101: data <= 11'h7fa; 
        10'b0101100110: data <= 11'h7f9; 
        10'b0101100111: data <= 11'h7fc; 
        10'b0101101000: data <= 11'h7ff; 
        10'b0101101001: data <= 11'h7ff; 
        10'b0101101010: data <= 11'h7ff; 
        10'b0101101011: data <= 11'h000; 
        10'b0101101100: data <= 11'h7ff; 
        10'b0101101101: data <= 11'h7ff; 
        10'b0101101110: data <= 11'h7ff; 
        10'b0101101111: data <= 11'h7ff; 
        10'b0101110000: data <= 11'h7fd; 
        10'b0101110001: data <= 11'h7fc; 
        10'b0101110010: data <= 11'h7f8; 
        10'b0101110011: data <= 11'h7f7; 
        10'b0101110100: data <= 11'h7fa; 
        10'b0101110101: data <= 11'h7ff; 
        10'b0101110110: data <= 11'h7fe; 
        10'b0101110111: data <= 11'h7fb; 
        10'b0101111000: data <= 11'h000; 
        10'b0101111001: data <= 11'h008; 
        10'b0101111010: data <= 11'h008; 
        10'b0101111011: data <= 11'h001; 
        10'b0101111100: data <= 11'h003; 
        10'b0101111101: data <= 11'h004; 
        10'b0101111110: data <= 11'h002; 
        10'b0101111111: data <= 11'h7fd; 
        10'b0110000000: data <= 11'h7f9; 
        10'b0110000001: data <= 11'h7f9; 
        10'b0110000010: data <= 11'h7fa; 
        10'b0110000011: data <= 11'h7fc; 
        10'b0110000100: data <= 11'h7fe; 
        10'b0110000101: data <= 11'h000; 
        10'b0110000110: data <= 11'h000; 
        10'b0110000111: data <= 11'h7ff; 
        10'b0110001000: data <= 11'h000; 
        10'b0110001001: data <= 11'h7fe; 
        10'b0110001010: data <= 11'h7ff; 
        10'b0110001011: data <= 11'h7ff; 
        10'b0110001100: data <= 11'h000; 
        10'b0110001101: data <= 11'h7fd; 
        10'b0110001110: data <= 11'h7f9; 
        10'b0110001111: data <= 11'h7f9; 
        10'b0110010000: data <= 11'h7fc; 
        10'b0110010001: data <= 11'h7ff; 
        10'b0110010010: data <= 11'h7fb; 
        10'b0110010011: data <= 11'h7fb; 
        10'b0110010100: data <= 11'h001; 
        10'b0110010101: data <= 11'h004; 
        10'b0110010110: data <= 11'h004; 
        10'b0110010111: data <= 11'h7ff; 
        10'b0110011000: data <= 11'h7fe; 
        10'b0110011001: data <= 11'h7ff; 
        10'b0110011010: data <= 11'h001; 
        10'b0110011011: data <= 11'h7fd; 
        10'b0110011100: data <= 11'h7fc; 
        10'b0110011101: data <= 11'h7fe; 
        10'b0110011110: data <= 11'h7fd; 
        10'b0110011111: data <= 11'h7fe; 
        10'b0110100000: data <= 11'h7fd; 
        10'b0110100001: data <= 11'h7fe; 
        10'b0110100010: data <= 11'h000; 
        10'b0110100011: data <= 11'h000; 
        10'b0110100100: data <= 11'h000; 
        10'b0110100101: data <= 11'h7fe; 
        10'b0110100110: data <= 11'h000; 
        10'b0110100111: data <= 11'h001; 
        10'b0110101000: data <= 11'h7ff; 
        10'b0110101001: data <= 11'h7fc; 
        10'b0110101010: data <= 11'h7f9; 
        10'b0110101011: data <= 11'h7f9; 
        10'b0110101100: data <= 11'h7fb; 
        10'b0110101101: data <= 11'h7fd; 
        10'b0110101110: data <= 11'h7fd; 
        10'b0110101111: data <= 11'h7ff; 
        10'b0110110000: data <= 11'h001; 
        10'b0110110001: data <= 11'h006; 
        10'b0110110010: data <= 11'h003; 
        10'b0110110011: data <= 11'h000; 
        10'b0110110100: data <= 11'h7fb; 
        10'b0110110101: data <= 11'h7ff; 
        10'b0110110110: data <= 11'h000; 
        10'b0110110111: data <= 11'h001; 
        10'b0110111000: data <= 11'h003; 
        10'b0110111001: data <= 11'h003; 
        10'b0110111010: data <= 11'h001; 
        10'b0110111011: data <= 11'h000; 
        10'b0110111100: data <= 11'h7fe; 
        10'b0110111101: data <= 11'h000; 
        10'b0110111110: data <= 11'h7ff; 
        10'b0110111111: data <= 11'h7fe; 
        10'b0111000000: data <= 11'h7ff; 
        10'b0111000001: data <= 11'h000; 
        10'b0111000010: data <= 11'h001; 
        10'b0111000011: data <= 11'h000; 
        10'b0111000100: data <= 11'h001; 
        10'b0111000101: data <= 11'h7fe; 
        10'b0111000110: data <= 11'h7fd; 
        10'b0111000111: data <= 11'h7fb; 
        10'b0111001000: data <= 11'h7f6; 
        10'b0111001001: data <= 11'h7f5; 
        10'b0111001010: data <= 11'h7f6; 
        10'b0111001011: data <= 11'h7fe; 
        10'b0111001100: data <= 11'h003; 
        10'b0111001101: data <= 11'h007; 
        10'b0111001110: data <= 11'h7ff; 
        10'b0111001111: data <= 11'h7fb; 
        10'b0111010000: data <= 11'h7fa; 
        10'b0111010001: data <= 11'h7fe; 
        10'b0111010010: data <= 11'h002; 
        10'b0111010011: data <= 11'h006; 
        10'b0111010100: data <= 11'h004; 
        10'b0111010101: data <= 11'h006; 
        10'b0111010110: data <= 11'h005; 
        10'b0111010111: data <= 11'h002; 
        10'b0111011000: data <= 11'h7ff; 
        10'b0111011001: data <= 11'h000; 
        10'b0111011010: data <= 11'h000; 
        10'b0111011011: data <= 11'h000; 
        10'b0111011100: data <= 11'h000; 
        10'b0111011101: data <= 11'h000; 
        10'b0111011110: data <= 11'h000; 
        10'b0111011111: data <= 11'h003; 
        10'b0111100000: data <= 11'h002; 
        10'b0111100001: data <= 11'h001; 
        10'b0111100010: data <= 11'h7fe; 
        10'b0111100011: data <= 11'h7fa; 
        10'b0111100100: data <= 11'h7f5; 
        10'b0111100101: data <= 11'h7ee; 
        10'b0111100110: data <= 11'h7ea; 
        10'b0111100111: data <= 11'h7ec; 
        10'b0111101000: data <= 11'h7f1; 
        10'b0111101001: data <= 11'h7f7; 
        10'b0111101010: data <= 11'h7f8; 
        10'b0111101011: data <= 11'h7f9; 
        10'b0111101100: data <= 11'h000; 
        10'b0111101101: data <= 11'h002; 
        10'b0111101110: data <= 11'h004; 
        10'b0111101111: data <= 11'h006; 
        10'b0111110000: data <= 11'h001; 
        10'b0111110001: data <= 11'h008; 
        10'b0111110010: data <= 11'h008; 
        10'b0111110011: data <= 11'h002; 
        10'b0111110100: data <= 11'h7ff; 
        10'b0111110101: data <= 11'h7fe; 
        10'b0111110110: data <= 11'h7fe; 
        10'b0111110111: data <= 11'h7ff; 
        10'b0111111000: data <= 11'h7ff; 
        10'b0111111001: data <= 11'h7ff; 
        10'b0111111010: data <= 11'h001; 
        10'b0111111011: data <= 11'h005; 
        10'b0111111100: data <= 11'h004; 
        10'b0111111101: data <= 11'h002; 
        10'b0111111110: data <= 11'h001; 
        10'b0111111111: data <= 11'h7ff; 
        10'b1000000000: data <= 11'h7fc; 
        10'b1000000001: data <= 11'h7f3; 
        10'b1000000010: data <= 11'h7ed; 
        10'b1000000011: data <= 11'h7ee; 
        10'b1000000100: data <= 11'h7ea; 
        10'b1000000101: data <= 11'h7ee; 
        10'b1000000110: data <= 11'h7f5; 
        10'b1000000111: data <= 11'h7fd; 
        10'b1000001000: data <= 11'h005; 
        10'b1000001001: data <= 11'h006; 
        10'b1000001010: data <= 11'h007; 
        10'b1000001011: data <= 11'h007; 
        10'b1000001100: data <= 11'h005; 
        10'b1000001101: data <= 11'h009; 
        10'b1000001110: data <= 11'h009; 
        10'b1000001111: data <= 11'h003; 
        10'b1000010000: data <= 11'h7fd; 
        10'b1000010001: data <= 11'h7fe; 
        10'b1000010010: data <= 11'h7ff; 
        10'b1000010011: data <= 11'h000; 
        10'b1000010100: data <= 11'h000; 
        10'b1000010101: data <= 11'h7ff; 
        10'b1000010110: data <= 11'h7ff; 
        10'b1000010111: data <= 11'h006; 
        10'b1000011000: data <= 11'h007; 
        10'b1000011001: data <= 11'h008; 
        10'b1000011010: data <= 11'h007; 
        10'b1000011011: data <= 11'h002; 
        10'b1000011100: data <= 11'h001; 
        10'b1000011101: data <= 11'h7fd; 
        10'b1000011110: data <= 11'h7fe; 
        10'b1000011111: data <= 11'h7fa; 
        10'b1000100000: data <= 11'h7f7; 
        10'b1000100001: data <= 11'h7f6; 
        10'b1000100010: data <= 11'h7f9; 
        10'b1000100011: data <= 11'h002; 
        10'b1000100100: data <= 11'h006; 
        10'b1000100101: data <= 11'h008; 
        10'b1000100110: data <= 11'h009; 
        10'b1000100111: data <= 11'h008; 
        10'b1000101000: data <= 11'h007; 
        10'b1000101001: data <= 11'h008; 
        10'b1000101010: data <= 11'h003; 
        10'b1000101011: data <= 11'h000; 
        10'b1000101100: data <= 11'h7fd; 
        10'b1000101101: data <= 11'h000; 
        10'b1000101110: data <= 11'h000; 
        10'b1000101111: data <= 11'h7ff; 
        10'b1000110000: data <= 11'h000; 
        10'b1000110001: data <= 11'h7fe; 
        10'b1000110010: data <= 11'h001; 
        10'b1000110011: data <= 11'h007; 
        10'b1000110100: data <= 11'h009; 
        10'b1000110101: data <= 11'h009; 
        10'b1000110110: data <= 11'h00a; 
        10'b1000110111: data <= 11'h005; 
        10'b1000111000: data <= 11'h006; 
        10'b1000111001: data <= 11'h007; 
        10'b1000111010: data <= 11'h002; 
        10'b1000111011: data <= 11'h7ff; 
        10'b1000111100: data <= 11'h7fe; 
        10'b1000111101: data <= 11'h7fd; 
        10'b1000111110: data <= 11'h001; 
        10'b1000111111: data <= 11'h002; 
        10'b1001000000: data <= 11'h003; 
        10'b1001000001: data <= 11'h006; 
        10'b1001000010: data <= 11'h006; 
        10'b1001000011: data <= 11'h004; 
        10'b1001000100: data <= 11'h008; 
        10'b1001000101: data <= 11'h004; 
        10'b1001000110: data <= 11'h7ff; 
        10'b1001000111: data <= 11'h7fe; 
        10'b1001001000: data <= 11'h7fe; 
        10'b1001001001: data <= 11'h7ff; 
        10'b1001001010: data <= 11'h7ff; 
        10'b1001001011: data <= 11'h7ff; 
        10'b1001001100: data <= 11'h7ff; 
        10'b1001001101: data <= 11'h000; 
        10'b1001001110: data <= 11'h000; 
        10'b1001001111: data <= 11'h003; 
        10'b1001010000: data <= 11'h008; 
        10'b1001010001: data <= 11'h008; 
        10'b1001010010: data <= 11'h007; 
        10'b1001010011: data <= 11'h004; 
        10'b1001010100: data <= 11'h004; 
        10'b1001010101: data <= 11'h001; 
        10'b1001010110: data <= 11'h7ff; 
        10'b1001010111: data <= 11'h7fe; 
        10'b1001011000: data <= 11'h001; 
        10'b1001011001: data <= 11'h000; 
        10'b1001011010: data <= 11'h7ff; 
        10'b1001011011: data <= 11'h7ff; 
        10'b1001011100: data <= 11'h002; 
        10'b1001011101: data <= 11'h001; 
        10'b1001011110: data <= 11'h004; 
        10'b1001011111: data <= 11'h006; 
        10'b1001100000: data <= 11'h004; 
        10'b1001100001: data <= 11'h001; 
        10'b1001100010: data <= 11'h7ff; 
        10'b1001100011: data <= 11'h7fc; 
        10'b1001100100: data <= 11'h7ff; 
        10'b1001100101: data <= 11'h7fe; 
        10'b1001100110: data <= 11'h7fe; 
        10'b1001100111: data <= 11'h7fe; 
        10'b1001101000: data <= 11'h7ff; 
        10'b1001101001: data <= 11'h7ff; 
        10'b1001101010: data <= 11'h000; 
        10'b1001101011: data <= 11'h002; 
        10'b1001101100: data <= 11'h004; 
        10'b1001101101: data <= 11'h006; 
        10'b1001101110: data <= 11'h005; 
        10'b1001101111: data <= 11'h003; 
        10'b1001110000: data <= 11'h000; 
        10'b1001110001: data <= 11'h002; 
        10'b1001110010: data <= 11'h003; 
        10'b1001110011: data <= 11'h003; 
        10'b1001110100: data <= 11'h001; 
        10'b1001110101: data <= 11'h7ff; 
        10'b1001110110: data <= 11'h7ff; 
        10'b1001110111: data <= 11'h7fe; 
        10'b1001111000: data <= 11'h001; 
        10'b1001111001: data <= 11'h001; 
        10'b1001111010: data <= 11'h001; 
        10'b1001111011: data <= 11'h004; 
        10'b1001111100: data <= 11'h002; 
        10'b1001111101: data <= 11'h7ff; 
        10'b1001111110: data <= 11'h7ff; 
        10'b1001111111: data <= 11'h7ff; 
        10'b1010000000: data <= 11'h7fd; 
        10'b1010000001: data <= 11'h7fe; 
        10'b1010000010: data <= 11'h000; 
        10'b1010000011: data <= 11'h000; 
        10'b1010000100: data <= 11'h7ff; 
        10'b1010000101: data <= 11'h7fe; 
        10'b1010000110: data <= 11'h7ff; 
        10'b1010000111: data <= 11'h001; 
        10'b1010001000: data <= 11'h005; 
        10'b1010001001: data <= 11'h007; 
        10'b1010001010: data <= 11'h005; 
        10'b1010001011: data <= 11'h005; 
        10'b1010001100: data <= 11'h001; 
        10'b1010001101: data <= 11'h003; 
        10'b1010001110: data <= 11'h002; 
        10'b1010001111: data <= 11'h000; 
        10'b1010010000: data <= 11'h7fe; 
        10'b1010010001: data <= 11'h000; 
        10'b1010010010: data <= 11'h001; 
        10'b1010010011: data <= 11'h002; 
        10'b1010010100: data <= 11'h001; 
        10'b1010010101: data <= 11'h003; 
        10'b1010010110: data <= 11'h004; 
        10'b1010010111: data <= 11'h7ff; 
        10'b1010011000: data <= 11'h7fd; 
        10'b1010011001: data <= 11'h7fd; 
        10'b1010011010: data <= 11'h7ff; 
        10'b1010011011: data <= 11'h7fe; 
        10'b1010011100: data <= 11'h000; 
        10'b1010011101: data <= 11'h000; 
        10'b1010011110: data <= 11'h7fe; 
        10'b1010011111: data <= 11'h7fe; 
        10'b1010100000: data <= 11'h7ff; 
        10'b1010100001: data <= 11'h000; 
        10'b1010100010: data <= 11'h000; 
        10'b1010100011: data <= 11'h000; 
        10'b1010100100: data <= 11'h003; 
        10'b1010100101: data <= 11'h005; 
        10'b1010100110: data <= 11'h006; 
        10'b1010100111: data <= 11'h007; 
        10'b1010101000: data <= 11'h007; 
        10'b1010101001: data <= 11'h005; 
        10'b1010101010: data <= 11'h008; 
        10'b1010101011: data <= 11'h008; 
        10'b1010101100: data <= 11'h009; 
        10'b1010101101: data <= 11'h007; 
        10'b1010101110: data <= 11'h006; 
        10'b1010101111: data <= 11'h004; 
        10'b1010110000: data <= 11'h004; 
        10'b1010110001: data <= 11'h000; 
        10'b1010110010: data <= 11'h7fd; 
        10'b1010110011: data <= 11'h7fb; 
        10'b1010110100: data <= 11'h7fc; 
        10'b1010110101: data <= 11'h7fd; 
        10'b1010110110: data <= 11'h7fe; 
        10'b1010110111: data <= 11'h7ff; 
        10'b1010111000: data <= 11'h7ff; 
        10'b1010111001: data <= 11'h000; 
        10'b1010111010: data <= 11'h7ff; 
        10'b1010111011: data <= 11'h000; 
        10'b1010111100: data <= 11'h000; 
        10'b1010111101: data <= 11'h7fe; 
        10'b1010111110: data <= 11'h000; 
        10'b1010111111: data <= 11'h000; 
        10'b1011000000: data <= 11'h7ff; 
        10'b1011000001: data <= 11'h002; 
        10'b1011000010: data <= 11'h003; 
        10'b1011000011: data <= 11'h002; 
        10'b1011000100: data <= 11'h004; 
        10'b1011000101: data <= 11'h004; 
        10'b1011000110: data <= 11'h007; 
        10'b1011000111: data <= 11'h008; 
        10'b1011001000: data <= 11'h009; 
        10'b1011001001: data <= 11'h007; 
        10'b1011001010: data <= 11'h005; 
        10'b1011001011: data <= 11'h002; 
        10'b1011001100: data <= 11'h7ff; 
        10'b1011001101: data <= 11'h7fd; 
        10'b1011001110: data <= 11'h7fd; 
        10'b1011001111: data <= 11'h7fe; 
        10'b1011010000: data <= 11'h7fe; 
        10'b1011010001: data <= 11'h7ff; 
        10'b1011010010: data <= 11'h7ff; 
        10'b1011010011: data <= 11'h000; 
        10'b1011010100: data <= 11'h7fe; 
        10'b1011010101: data <= 11'h000; 
        10'b1011010110: data <= 11'h7fe; 
        10'b1011010111: data <= 11'h000; 
        10'b1011011000: data <= 11'h7ff; 
        10'b1011011001: data <= 11'h7fe; 
        10'b1011011010: data <= 11'h7fe; 
        10'b1011011011: data <= 11'h000; 
        10'b1011011100: data <= 11'h000; 
        10'b1011011101: data <= 11'h7ff; 
        10'b1011011110: data <= 11'h7fe; 
        10'b1011011111: data <= 11'h7ff; 
        10'b1011100000: data <= 11'h000; 
        10'b1011100001: data <= 11'h7ff; 
        10'b1011100010: data <= 11'h7ff; 
        10'b1011100011: data <= 11'h7ff; 
        10'b1011100100: data <= 11'h7ff; 
        10'b1011100101: data <= 11'h7ff; 
        10'b1011100110: data <= 11'h7ff; 
        10'b1011100111: data <= 11'h7fe; 
        10'b1011101000: data <= 11'h7ff; 
        10'b1011101001: data <= 11'h7ff; 
        10'b1011101010: data <= 11'h7ff; 
        10'b1011101011: data <= 11'h7ff; 
        10'b1011101100: data <= 11'h7fe; 
        10'b1011101101: data <= 11'h7fe; 
        10'b1011101110: data <= 11'h000; 
        10'b1011101111: data <= 11'h7ff; 
        10'b1011110000: data <= 11'h000; 
        10'b1011110001: data <= 11'h7ff; 
        10'b1011110010: data <= 11'h000; 
        10'b1011110011: data <= 11'h000; 
        10'b1011110100: data <= 11'h7ff; 
        10'b1011110101: data <= 11'h7fe; 
        10'b1011110110: data <= 11'h7ff; 
        10'b1011110111: data <= 11'h7fe; 
        10'b1011111000: data <= 11'h000; 
        10'b1011111001: data <= 11'h7ff; 
        10'b1011111010: data <= 11'h000; 
        10'b1011111011: data <= 11'h7ff; 
        10'b1011111100: data <= 11'h000; 
        10'b1011111101: data <= 11'h7fe; 
        10'b1011111110: data <= 11'h7fe; 
        10'b1011111111: data <= 11'h000; 
        10'b1100000000: data <= 11'h7fe; 
        10'b1100000001: data <= 11'h000; 
        10'b1100000010: data <= 11'h7ff; 
        10'b1100000011: data <= 11'h7ff; 
        10'b1100000100: data <= 11'h7ff; 
        10'b1100000101: data <= 11'h000; 
        10'b1100000110: data <= 11'h7fe; 
        10'b1100000111: data <= 11'h7fe; 
        10'b1100001000: data <= 11'h000; 
        10'b1100001001: data <= 11'h7ff; 
        10'b1100001010: data <= 11'h7fe; 
        10'b1100001011: data <= 11'h000; 
        10'b1100001100: data <= 11'h7fe; 
        10'b1100001101: data <= 11'h7fe; 
        10'b1100001110: data <= 11'h000; 
        10'b1100001111: data <= 11'h7ff; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 6) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 12'hfff; 
        10'b0000000001: data <= 12'hffd; 
        10'b0000000010: data <= 12'h000; 
        10'b0000000011: data <= 12'h000; 
        10'b0000000100: data <= 12'h000; 
        10'b0000000101: data <= 12'h000; 
        10'b0000000110: data <= 12'hfff; 
        10'b0000000111: data <= 12'h000; 
        10'b0000001000: data <= 12'hffd; 
        10'b0000001001: data <= 12'h000; 
        10'b0000001010: data <= 12'h000; 
        10'b0000001011: data <= 12'hffe; 
        10'b0000001100: data <= 12'hffe; 
        10'b0000001101: data <= 12'hffe; 
        10'b0000001110: data <= 12'hffe; 
        10'b0000001111: data <= 12'hffe; 
        10'b0000010000: data <= 12'h000; 
        10'b0000010001: data <= 12'h000; 
        10'b0000010010: data <= 12'hffd; 
        10'b0000010011: data <= 12'h000; 
        10'b0000010100: data <= 12'hfff; 
        10'b0000010101: data <= 12'hfff; 
        10'b0000010110: data <= 12'hffc; 
        10'b0000010111: data <= 12'h000; 
        10'b0000011000: data <= 12'h000; 
        10'b0000011001: data <= 12'hffc; 
        10'b0000011010: data <= 12'hffe; 
        10'b0000011011: data <= 12'h000; 
        10'b0000011100: data <= 12'hffd; 
        10'b0000011101: data <= 12'hffe; 
        10'b0000011110: data <= 12'hffd; 
        10'b0000011111: data <= 12'hfff; 
        10'b0000100000: data <= 12'hffc; 
        10'b0000100001: data <= 12'hffe; 
        10'b0000100010: data <= 12'h000; 
        10'b0000100011: data <= 12'h000; 
        10'b0000100100: data <= 12'hffc; 
        10'b0000100101: data <= 12'hffc; 
        10'b0000100110: data <= 12'hffc; 
        10'b0000100111: data <= 12'hfff; 
        10'b0000101000: data <= 12'hfff; 
        10'b0000101001: data <= 12'hffe; 
        10'b0000101010: data <= 12'hffe; 
        10'b0000101011: data <= 12'hffd; 
        10'b0000101100: data <= 12'h000; 
        10'b0000101101: data <= 12'hffd; 
        10'b0000101110: data <= 12'hfff; 
        10'b0000101111: data <= 12'hffe; 
        10'b0000110000: data <= 12'hffe; 
        10'b0000110001: data <= 12'hffc; 
        10'b0000110010: data <= 12'hffe; 
        10'b0000110011: data <= 12'h000; 
        10'b0000110100: data <= 12'hffd; 
        10'b0000110101: data <= 12'h000; 
        10'b0000110110: data <= 12'hfff; 
        10'b0000110111: data <= 12'hffd; 
        10'b0000111000: data <= 12'hffd; 
        10'b0000111001: data <= 12'hffe; 
        10'b0000111010: data <= 12'hffe; 
        10'b0000111011: data <= 12'hffd; 
        10'b0000111100: data <= 12'hfff; 
        10'b0000111101: data <= 12'hfff; 
        10'b0000111110: data <= 12'hffd; 
        10'b0000111111: data <= 12'hfff; 
        10'b0001000000: data <= 12'h000; 
        10'b0001000001: data <= 12'hffe; 
        10'b0001000010: data <= 12'hffd; 
        10'b0001000011: data <= 12'hffd; 
        10'b0001000100: data <= 12'hffc; 
        10'b0001000101: data <= 12'hffd; 
        10'b0001000110: data <= 12'hffe; 
        10'b0001000111: data <= 12'hffe; 
        10'b0001001000: data <= 12'hffd; 
        10'b0001001001: data <= 12'hffd; 
        10'b0001001010: data <= 12'hfff; 
        10'b0001001011: data <= 12'h000; 
        10'b0001001100: data <= 12'hffe; 
        10'b0001001101: data <= 12'hffd; 
        10'b0001001110: data <= 12'h000; 
        10'b0001001111: data <= 12'h000; 
        10'b0001010000: data <= 12'h000; 
        10'b0001010001: data <= 12'hffe; 
        10'b0001010010: data <= 12'hffc; 
        10'b0001010011: data <= 12'hffe; 
        10'b0001010100: data <= 12'h000; 
        10'b0001010101: data <= 12'hfff; 
        10'b0001010110: data <= 12'hffe; 
        10'b0001010111: data <= 12'h000; 
        10'b0001011000: data <= 12'hfff; 
        10'b0001011001: data <= 12'h000; 
        10'b0001011010: data <= 12'hfff; 
        10'b0001011011: data <= 12'h000; 
        10'b0001011100: data <= 12'h000; 
        10'b0001011101: data <= 12'hfff; 
        10'b0001011110: data <= 12'h001; 
        10'b0001011111: data <= 12'h005; 
        10'b0001100000: data <= 12'h00a; 
        10'b0001100001: data <= 12'h008; 
        10'b0001100010: data <= 12'h008; 
        10'b0001100011: data <= 12'h009; 
        10'b0001100100: data <= 12'h006; 
        10'b0001100101: data <= 12'h007; 
        10'b0001100110: data <= 12'h006; 
        10'b0001100111: data <= 12'h000; 
        10'b0001101000: data <= 12'hfff; 
        10'b0001101001: data <= 12'hff9; 
        10'b0001101010: data <= 12'hffc; 
        10'b0001101011: data <= 12'h000; 
        10'b0001101100: data <= 12'h000; 
        10'b0001101101: data <= 12'hffd; 
        10'b0001101110: data <= 12'hfff; 
        10'b0001101111: data <= 12'hffd; 
        10'b0001110000: data <= 12'hfff; 
        10'b0001110001: data <= 12'h000; 
        10'b0001110010: data <= 12'hfff; 
        10'b0001110011: data <= 12'h000; 
        10'b0001110100: data <= 12'h001; 
        10'b0001110101: data <= 12'h000; 
        10'b0001110110: data <= 12'h006; 
        10'b0001110111: data <= 12'h005; 
        10'b0001111000: data <= 12'h00d; 
        10'b0001111001: data <= 12'h00b; 
        10'b0001111010: data <= 12'h00e; 
        10'b0001111011: data <= 12'h011; 
        10'b0001111100: data <= 12'h014; 
        10'b0001111101: data <= 12'h015; 
        10'b0001111110: data <= 12'h013; 
        10'b0001111111: data <= 12'h00e; 
        10'b0010000000: data <= 12'h008; 
        10'b0010000001: data <= 12'h006; 
        10'b0010000010: data <= 12'h00a; 
        10'b0010000011: data <= 12'h001; 
        10'b0010000100: data <= 12'hff9; 
        10'b0010000101: data <= 12'hff5; 
        10'b0010000110: data <= 12'hff7; 
        10'b0010000111: data <= 12'hff7; 
        10'b0010001000: data <= 12'hfff; 
        10'b0010001001: data <= 12'hffe; 
        10'b0010001010: data <= 12'hffe; 
        10'b0010001011: data <= 12'hfff; 
        10'b0010001100: data <= 12'hffd; 
        10'b0010001101: data <= 12'hffc; 
        10'b0010001110: data <= 12'hffd; 
        10'b0010001111: data <= 12'hffd; 
        10'b0010010000: data <= 12'h001; 
        10'b0010010001: data <= 12'h006; 
        10'b0010010010: data <= 12'h00b; 
        10'b0010010011: data <= 12'h009; 
        10'b0010010100: data <= 12'h00a; 
        10'b0010010101: data <= 12'h009; 
        10'b0010010110: data <= 12'h008; 
        10'b0010010111: data <= 12'h00a; 
        10'b0010011000: data <= 12'h00b; 
        10'b0010011001: data <= 12'h00d; 
        10'b0010011010: data <= 12'h002; 
        10'b0010011011: data <= 12'h008; 
        10'b0010011100: data <= 12'h00a; 
        10'b0010011101: data <= 12'hfff; 
        10'b0010011110: data <= 12'hfff; 
        10'b0010011111: data <= 12'hffc; 
        10'b0010100000: data <= 12'hffa; 
        10'b0010100001: data <= 12'hff3; 
        10'b0010100010: data <= 12'hfef; 
        10'b0010100011: data <= 12'hff2; 
        10'b0010100100: data <= 12'hffc; 
        10'b0010100101: data <= 12'h000; 
        10'b0010100110: data <= 12'hffd; 
        10'b0010100111: data <= 12'hffe; 
        10'b0010101000: data <= 12'hffd; 
        10'b0010101001: data <= 12'hffe; 
        10'b0010101010: data <= 12'hffd; 
        10'b0010101011: data <= 12'h001; 
        10'b0010101100: data <= 12'h007; 
        10'b0010101101: data <= 12'h00e; 
        10'b0010101110: data <= 12'h00b; 
        10'b0010101111: data <= 12'h008; 
        10'b0010110000: data <= 12'h00c; 
        10'b0010110001: data <= 12'h00a; 
        10'b0010110010: data <= 12'h009; 
        10'b0010110011: data <= 12'h008; 
        10'b0010110100: data <= 12'h00b; 
        10'b0010110101: data <= 12'h010; 
        10'b0010110110: data <= 12'h00b; 
        10'b0010110111: data <= 12'h004; 
        10'b0010111000: data <= 12'h00b; 
        10'b0010111001: data <= 12'h00a; 
        10'b0010111010: data <= 12'h009; 
        10'b0010111011: data <= 12'hffc; 
        10'b0010111100: data <= 12'h004; 
        10'b0010111101: data <= 12'hffc; 
        10'b0010111110: data <= 12'hff2; 
        10'b0010111111: data <= 12'hff2; 
        10'b0011000000: data <= 12'hff7; 
        10'b0011000001: data <= 12'hffe; 
        10'b0011000010: data <= 12'h000; 
        10'b0011000011: data <= 12'hfff; 
        10'b0011000100: data <= 12'h000; 
        10'b0011000101: data <= 12'h000; 
        10'b0011000110: data <= 12'h001; 
        10'b0011000111: data <= 12'h006; 
        10'b0011001000: data <= 12'h010; 
        10'b0011001001: data <= 12'h010; 
        10'b0011001010: data <= 12'h00b; 
        10'b0011001011: data <= 12'h003; 
        10'b0011001100: data <= 12'h003; 
        10'b0011001101: data <= 12'h007; 
        10'b0011001110: data <= 12'h002; 
        10'b0011001111: data <= 12'h003; 
        10'b0011010000: data <= 12'h00a; 
        10'b0011010001: data <= 12'h009; 
        10'b0011010010: data <= 12'h00f; 
        10'b0011010011: data <= 12'h009; 
        10'b0011010100: data <= 12'h003; 
        10'b0011010101: data <= 12'h008; 
        10'b0011010110: data <= 12'h006; 
        10'b0011010111: data <= 12'h007; 
        10'b0011011000: data <= 12'h007; 
        10'b0011011001: data <= 12'h001; 
        10'b0011011010: data <= 12'hff9; 
        10'b0011011011: data <= 12'hff0; 
        10'b0011011100: data <= 12'hff5; 
        10'b0011011101: data <= 12'hffd; 
        10'b0011011110: data <= 12'hffc; 
        10'b0011011111: data <= 12'hffe; 
        10'b0011100000: data <= 12'hffe; 
        10'b0011100001: data <= 12'hffe; 
        10'b0011100010: data <= 12'h001; 
        10'b0011100011: data <= 12'h006; 
        10'b0011100100: data <= 12'h00d; 
        10'b0011100101: data <= 12'h00d; 
        10'b0011100110: data <= 12'h00a; 
        10'b0011100111: data <= 12'h004; 
        10'b0011101000: data <= 12'h006; 
        10'b0011101001: data <= 12'h003; 
        10'b0011101010: data <= 12'h008; 
        10'b0011101011: data <= 12'h003; 
        10'b0011101100: data <= 12'h002; 
        10'b0011101101: data <= 12'h004; 
        10'b0011101110: data <= 12'h010; 
        10'b0011101111: data <= 12'h00d; 
        10'b0011110000: data <= 12'h003; 
        10'b0011110001: data <= 12'h007; 
        10'b0011110010: data <= 12'h00b; 
        10'b0011110011: data <= 12'h007; 
        10'b0011110100: data <= 12'h00a; 
        10'b0011110101: data <= 12'h005; 
        10'b0011110110: data <= 12'hffd; 
        10'b0011110111: data <= 12'hff1; 
        10'b0011111000: data <= 12'hff5; 
        10'b0011111001: data <= 12'hffc; 
        10'b0011111010: data <= 12'hffd; 
        10'b0011111011: data <= 12'hffe; 
        10'b0011111100: data <= 12'hffe; 
        10'b0011111101: data <= 12'hffc; 
        10'b0011111110: data <= 12'hfff; 
        10'b0011111111: data <= 12'h002; 
        10'b0100000000: data <= 12'h007; 
        10'b0100000001: data <= 12'h009; 
        10'b0100000010: data <= 12'h008; 
        10'b0100000011: data <= 12'h002; 
        10'b0100000100: data <= 12'hfff; 
        10'b0100000101: data <= 12'hff9; 
        10'b0100000110: data <= 12'hff2; 
        10'b0100000111: data <= 12'hfe7; 
        10'b0100001000: data <= 12'hfec; 
        10'b0100001001: data <= 12'hffd; 
        10'b0100001010: data <= 12'h013; 
        10'b0100001011: data <= 12'h01e; 
        10'b0100001100: data <= 12'h011; 
        10'b0100001101: data <= 12'h00a; 
        10'b0100001110: data <= 12'h00b; 
        10'b0100001111: data <= 12'h00a; 
        10'b0100010000: data <= 12'h00f; 
        10'b0100010001: data <= 12'h00a; 
        10'b0100010010: data <= 12'hffd; 
        10'b0100010011: data <= 12'hff1; 
        10'b0100010100: data <= 12'hff9; 
        10'b0100010101: data <= 12'hffc; 
        10'b0100010110: data <= 12'hffd; 
        10'b0100010111: data <= 12'hffd; 
        10'b0100011000: data <= 12'h000; 
        10'b0100011001: data <= 12'hfff; 
        10'b0100011010: data <= 12'h000; 
        10'b0100011011: data <= 12'h004; 
        10'b0100011100: data <= 12'h003; 
        10'b0100011101: data <= 12'h001; 
        10'b0100011110: data <= 12'hffc; 
        10'b0100011111: data <= 12'hff5; 
        10'b0100100000: data <= 12'hfec; 
        10'b0100100001: data <= 12'hfe3; 
        10'b0100100010: data <= 12'hfdd; 
        10'b0100100011: data <= 12'hfdc; 
        10'b0100100100: data <= 12'hfe5; 
        10'b0100100101: data <= 12'hff9; 
        10'b0100100110: data <= 12'h010; 
        10'b0100100111: data <= 12'h012; 
        10'b0100101000: data <= 12'h010; 
        10'b0100101001: data <= 12'h00f; 
        10'b0100101010: data <= 12'h009; 
        10'b0100101011: data <= 12'h010; 
        10'b0100101100: data <= 12'h00e; 
        10'b0100101101: data <= 12'h006; 
        10'b0100101110: data <= 12'hffb; 
        10'b0100101111: data <= 12'hff6; 
        10'b0100110000: data <= 12'hffc; 
        10'b0100110001: data <= 12'hffc; 
        10'b0100110010: data <= 12'hffe; 
        10'b0100110011: data <= 12'h000; 
        10'b0100110100: data <= 12'h000; 
        10'b0100110101: data <= 12'h000; 
        10'b0100110110: data <= 12'hffd; 
        10'b0100110111: data <= 12'h004; 
        10'b0100111000: data <= 12'hffe; 
        10'b0100111001: data <= 12'hff5; 
        10'b0100111010: data <= 12'hfef; 
        10'b0100111011: data <= 12'hfe7; 
        10'b0100111100: data <= 12'hfe1; 
        10'b0100111101: data <= 12'hfe5; 
        10'b0100111110: data <= 12'hfec; 
        10'b0100111111: data <= 12'hff6; 
        10'b0101000000: data <= 12'hffb; 
        10'b0101000001: data <= 12'h007; 
        10'b0101000010: data <= 12'h00b; 
        10'b0101000011: data <= 12'h00b; 
        10'b0101000100: data <= 12'h005; 
        10'b0101000101: data <= 12'h00b; 
        10'b0101000110: data <= 12'h00e; 
        10'b0101000111: data <= 12'h00d; 
        10'b0101001000: data <= 12'h00c; 
        10'b0101001001: data <= 12'h000; 
        10'b0101001010: data <= 12'hffb; 
        10'b0101001011: data <= 12'hffc; 
        10'b0101001100: data <= 12'hffc; 
        10'b0101001101: data <= 12'hffe; 
        10'b0101001110: data <= 12'hffd; 
        10'b0101001111: data <= 12'hffd; 
        10'b0101010000: data <= 12'h000; 
        10'b0101010001: data <= 12'hffd; 
        10'b0101010010: data <= 12'hfff; 
        10'b0101010011: data <= 12'h000; 
        10'b0101010100: data <= 12'hffc; 
        10'b0101010101: data <= 12'hff5; 
        10'b0101010110: data <= 12'hfec; 
        10'b0101010111: data <= 12'hfe7; 
        10'b0101011000: data <= 12'hfea; 
        10'b0101011001: data <= 12'hff4; 
        10'b0101011010: data <= 12'h000; 
        10'b0101011011: data <= 12'h002; 
        10'b0101011100: data <= 12'h003; 
        10'b0101011101: data <= 12'h007; 
        10'b0101011110: data <= 12'h012; 
        10'b0101011111: data <= 12'h009; 
        10'b0101100000: data <= 12'h006; 
        10'b0101100001: data <= 12'h009; 
        10'b0101100010: data <= 12'h007; 
        10'b0101100011: data <= 12'hfff; 
        10'b0101100100: data <= 12'hff7; 
        10'b0101100101: data <= 12'hff3; 
        10'b0101100110: data <= 12'hff3; 
        10'b0101100111: data <= 12'hff8; 
        10'b0101101000: data <= 12'hfff; 
        10'b0101101001: data <= 12'hffd; 
        10'b0101101010: data <= 12'hfff; 
        10'b0101101011: data <= 12'hfff; 
        10'b0101101100: data <= 12'hffe; 
        10'b0101101101: data <= 12'hffd; 
        10'b0101101110: data <= 12'hffe; 
        10'b0101101111: data <= 12'hfff; 
        10'b0101110000: data <= 12'hffb; 
        10'b0101110001: data <= 12'hff8; 
        10'b0101110010: data <= 12'hff0; 
        10'b0101110011: data <= 12'hfed; 
        10'b0101110100: data <= 12'hff3; 
        10'b0101110101: data <= 12'hffe; 
        10'b0101110110: data <= 12'hffc; 
        10'b0101110111: data <= 12'hff5; 
        10'b0101111000: data <= 12'h001; 
        10'b0101111001: data <= 12'h00f; 
        10'b0101111010: data <= 12'h00f; 
        10'b0101111011: data <= 12'h003; 
        10'b0101111100: data <= 12'h007; 
        10'b0101111101: data <= 12'h007; 
        10'b0101111110: data <= 12'h004; 
        10'b0101111111: data <= 12'hffb; 
        10'b0110000000: data <= 12'hff2; 
        10'b0110000001: data <= 12'hff2; 
        10'b0110000010: data <= 12'hff5; 
        10'b0110000011: data <= 12'hff8; 
        10'b0110000100: data <= 12'hffc; 
        10'b0110000101: data <= 12'h000; 
        10'b0110000110: data <= 12'hfff; 
        10'b0110000111: data <= 12'hffe; 
        10'b0110001000: data <= 12'h000; 
        10'b0110001001: data <= 12'hffd; 
        10'b0110001010: data <= 12'hffe; 
        10'b0110001011: data <= 12'hfff; 
        10'b0110001100: data <= 12'hfff; 
        10'b0110001101: data <= 12'hffa; 
        10'b0110001110: data <= 12'hff2; 
        10'b0110001111: data <= 12'hff3; 
        10'b0110010000: data <= 12'hff7; 
        10'b0110010001: data <= 12'hfff; 
        10'b0110010010: data <= 12'hff7; 
        10'b0110010011: data <= 12'hff6; 
        10'b0110010100: data <= 12'h003; 
        10'b0110010101: data <= 12'h007; 
        10'b0110010110: data <= 12'h008; 
        10'b0110010111: data <= 12'hfff; 
        10'b0110011000: data <= 12'hffd; 
        10'b0110011001: data <= 12'hffe; 
        10'b0110011010: data <= 12'h001; 
        10'b0110011011: data <= 12'hffa; 
        10'b0110011100: data <= 12'hff8; 
        10'b0110011101: data <= 12'hffc; 
        10'b0110011110: data <= 12'hffa; 
        10'b0110011111: data <= 12'hffc; 
        10'b0110100000: data <= 12'hffb; 
        10'b0110100001: data <= 12'hffb; 
        10'b0110100010: data <= 12'h000; 
        10'b0110100011: data <= 12'h000; 
        10'b0110100100: data <= 12'h000; 
        10'b0110100101: data <= 12'hffd; 
        10'b0110100110: data <= 12'h000; 
        10'b0110100111: data <= 12'h001; 
        10'b0110101000: data <= 12'hfff; 
        10'b0110101001: data <= 12'hff9; 
        10'b0110101010: data <= 12'hff3; 
        10'b0110101011: data <= 12'hff2; 
        10'b0110101100: data <= 12'hff5; 
        10'b0110101101: data <= 12'hffa; 
        10'b0110101110: data <= 12'hff9; 
        10'b0110101111: data <= 12'hffe; 
        10'b0110110000: data <= 12'h003; 
        10'b0110110001: data <= 12'h00c; 
        10'b0110110010: data <= 12'h007; 
        10'b0110110011: data <= 12'hfff; 
        10'b0110110100: data <= 12'hff6; 
        10'b0110110101: data <= 12'hffd; 
        10'b0110110110: data <= 12'hfff; 
        10'b0110110111: data <= 12'h003; 
        10'b0110111000: data <= 12'h006; 
        10'b0110111001: data <= 12'h006; 
        10'b0110111010: data <= 12'h002; 
        10'b0110111011: data <= 12'h001; 
        10'b0110111100: data <= 12'hffc; 
        10'b0110111101: data <= 12'hfff; 
        10'b0110111110: data <= 12'hfff; 
        10'b0110111111: data <= 12'hffd; 
        10'b0111000000: data <= 12'hfff; 
        10'b0111000001: data <= 12'hfff; 
        10'b0111000010: data <= 12'h003; 
        10'b0111000011: data <= 12'h000; 
        10'b0111000100: data <= 12'h002; 
        10'b0111000101: data <= 12'hffd; 
        10'b0111000110: data <= 12'hffb; 
        10'b0111000111: data <= 12'hff6; 
        10'b0111001000: data <= 12'hfeb; 
        10'b0111001001: data <= 12'hfea; 
        10'b0111001010: data <= 12'hfed; 
        10'b0111001011: data <= 12'hffb; 
        10'b0111001100: data <= 12'h006; 
        10'b0111001101: data <= 12'h00f; 
        10'b0111001110: data <= 12'hffe; 
        10'b0111001111: data <= 12'hff5; 
        10'b0111010000: data <= 12'hff4; 
        10'b0111010001: data <= 12'hffc; 
        10'b0111010010: data <= 12'h005; 
        10'b0111010011: data <= 12'h00d; 
        10'b0111010100: data <= 12'h009; 
        10'b0111010101: data <= 12'h00b; 
        10'b0111010110: data <= 12'h00b; 
        10'b0111010111: data <= 12'h005; 
        10'b0111011000: data <= 12'hfff; 
        10'b0111011001: data <= 12'hfff; 
        10'b0111011010: data <= 12'h000; 
        10'b0111011011: data <= 12'h000; 
        10'b0111011100: data <= 12'h000; 
        10'b0111011101: data <= 12'h000; 
        10'b0111011110: data <= 12'h000; 
        10'b0111011111: data <= 12'h007; 
        10'b0111100000: data <= 12'h004; 
        10'b0111100001: data <= 12'h001; 
        10'b0111100010: data <= 12'hffc; 
        10'b0111100011: data <= 12'hff3; 
        10'b0111100100: data <= 12'hfea; 
        10'b0111100101: data <= 12'hfdd; 
        10'b0111100110: data <= 12'hfd4; 
        10'b0111100111: data <= 12'hfd8; 
        10'b0111101000: data <= 12'hfe1; 
        10'b0111101001: data <= 12'hfef; 
        10'b0111101010: data <= 12'hff0; 
        10'b0111101011: data <= 12'hff2; 
        10'b0111101100: data <= 12'hfff; 
        10'b0111101101: data <= 12'h004; 
        10'b0111101110: data <= 12'h008; 
        10'b0111101111: data <= 12'h00d; 
        10'b0111110000: data <= 12'h003; 
        10'b0111110001: data <= 12'h010; 
        10'b0111110010: data <= 12'h010; 
        10'b0111110011: data <= 12'h005; 
        10'b0111110100: data <= 12'hffe; 
        10'b0111110101: data <= 12'hffd; 
        10'b0111110110: data <= 12'hffd; 
        10'b0111110111: data <= 12'hffd; 
        10'b0111111000: data <= 12'hffe; 
        10'b0111111001: data <= 12'hffe; 
        10'b0111111010: data <= 12'h001; 
        10'b0111111011: data <= 12'h00a; 
        10'b0111111100: data <= 12'h007; 
        10'b0111111101: data <= 12'h004; 
        10'b0111111110: data <= 12'h002; 
        10'b0111111111: data <= 12'hffd; 
        10'b1000000000: data <= 12'hff8; 
        10'b1000000001: data <= 12'hfe6; 
        10'b1000000010: data <= 12'hfda; 
        10'b1000000011: data <= 12'hfdc; 
        10'b1000000100: data <= 12'hfd4; 
        10'b1000000101: data <= 12'hfdc; 
        10'b1000000110: data <= 12'hfe9; 
        10'b1000000111: data <= 12'hffb; 
        10'b1000001000: data <= 12'h009; 
        10'b1000001001: data <= 12'h00c; 
        10'b1000001010: data <= 12'h00d; 
        10'b1000001011: data <= 12'h00d; 
        10'b1000001100: data <= 12'h009; 
        10'b1000001101: data <= 12'h012; 
        10'b1000001110: data <= 12'h011; 
        10'b1000001111: data <= 12'h007; 
        10'b1000010000: data <= 12'hffa; 
        10'b1000010001: data <= 12'hffc; 
        10'b1000010010: data <= 12'hffd; 
        10'b1000010011: data <= 12'h000; 
        10'b1000010100: data <= 12'h000; 
        10'b1000010101: data <= 12'hffd; 
        10'b1000010110: data <= 12'hffe; 
        10'b1000010111: data <= 12'h00d; 
        10'b1000011000: data <= 12'h00d; 
        10'b1000011001: data <= 12'h010; 
        10'b1000011010: data <= 12'h00d; 
        10'b1000011011: data <= 12'h005; 
        10'b1000011100: data <= 12'h001; 
        10'b1000011101: data <= 12'hffb; 
        10'b1000011110: data <= 12'hffc; 
        10'b1000011111: data <= 12'hff4; 
        10'b1000100000: data <= 12'hfee; 
        10'b1000100001: data <= 12'hfed; 
        10'b1000100010: data <= 12'hff3; 
        10'b1000100011: data <= 12'h005; 
        10'b1000100100: data <= 12'h00c; 
        10'b1000100101: data <= 12'h00f; 
        10'b1000100110: data <= 12'h011; 
        10'b1000100111: data <= 12'h00f; 
        10'b1000101000: data <= 12'h00e; 
        10'b1000101001: data <= 12'h010; 
        10'b1000101010: data <= 12'h006; 
        10'b1000101011: data <= 12'h001; 
        10'b1000101100: data <= 12'hffb; 
        10'b1000101101: data <= 12'hfff; 
        10'b1000101110: data <= 12'hfff; 
        10'b1000101111: data <= 12'hfff; 
        10'b1000110000: data <= 12'hfff; 
        10'b1000110001: data <= 12'hffc; 
        10'b1000110010: data <= 12'h002; 
        10'b1000110011: data <= 12'h00e; 
        10'b1000110100: data <= 12'h011; 
        10'b1000110101: data <= 12'h012; 
        10'b1000110110: data <= 12'h014; 
        10'b1000110111: data <= 12'h00a; 
        10'b1000111000: data <= 12'h00c; 
        10'b1000111001: data <= 12'h00d; 
        10'b1000111010: data <= 12'h005; 
        10'b1000111011: data <= 12'hfff; 
        10'b1000111100: data <= 12'hffc; 
        10'b1000111101: data <= 12'hff9; 
        10'b1000111110: data <= 12'h002; 
        10'b1000111111: data <= 12'h004; 
        10'b1001000000: data <= 12'h007; 
        10'b1001000001: data <= 12'h00c; 
        10'b1001000010: data <= 12'h00d; 
        10'b1001000011: data <= 12'h009; 
        10'b1001000100: data <= 12'h00f; 
        10'b1001000101: data <= 12'h009; 
        10'b1001000110: data <= 12'hffe; 
        10'b1001000111: data <= 12'hffd; 
        10'b1001001000: data <= 12'hffc; 
        10'b1001001001: data <= 12'hfff; 
        10'b1001001010: data <= 12'hfff; 
        10'b1001001011: data <= 12'hfff; 
        10'b1001001100: data <= 12'hffd; 
        10'b1001001101: data <= 12'h000; 
        10'b1001001110: data <= 12'hfff; 
        10'b1001001111: data <= 12'h007; 
        10'b1001010000: data <= 12'h010; 
        10'b1001010001: data <= 12'h010; 
        10'b1001010010: data <= 12'h00e; 
        10'b1001010011: data <= 12'h008; 
        10'b1001010100: data <= 12'h009; 
        10'b1001010101: data <= 12'h003; 
        10'b1001010110: data <= 12'hfff; 
        10'b1001010111: data <= 12'hffc; 
        10'b1001011000: data <= 12'h001; 
        10'b1001011001: data <= 12'hfff; 
        10'b1001011010: data <= 12'hfff; 
        10'b1001011011: data <= 12'hffe; 
        10'b1001011100: data <= 12'h004; 
        10'b1001011101: data <= 12'h001; 
        10'b1001011110: data <= 12'h008; 
        10'b1001011111: data <= 12'h00d; 
        10'b1001100000: data <= 12'h007; 
        10'b1001100001: data <= 12'h003; 
        10'b1001100010: data <= 12'hffd; 
        10'b1001100011: data <= 12'hff9; 
        10'b1001100100: data <= 12'hffe; 
        10'b1001100101: data <= 12'hffd; 
        10'b1001100110: data <= 12'hffc; 
        10'b1001100111: data <= 12'hffc; 
        10'b1001101000: data <= 12'hffe; 
        10'b1001101001: data <= 12'hfff; 
        10'b1001101010: data <= 12'hfff; 
        10'b1001101011: data <= 12'h004; 
        10'b1001101100: data <= 12'h008; 
        10'b1001101101: data <= 12'h00b; 
        10'b1001101110: data <= 12'h00a; 
        10'b1001101111: data <= 12'h006; 
        10'b1001110000: data <= 12'h000; 
        10'b1001110001: data <= 12'h004; 
        10'b1001110010: data <= 12'h005; 
        10'b1001110011: data <= 12'h006; 
        10'b1001110100: data <= 12'h002; 
        10'b1001110101: data <= 12'hffe; 
        10'b1001110110: data <= 12'hffe; 
        10'b1001110111: data <= 12'hffd; 
        10'b1001111000: data <= 12'h003; 
        10'b1001111001: data <= 12'h002; 
        10'b1001111010: data <= 12'h002; 
        10'b1001111011: data <= 12'h009; 
        10'b1001111100: data <= 12'h004; 
        10'b1001111101: data <= 12'hffe; 
        10'b1001111110: data <= 12'hffe; 
        10'b1001111111: data <= 12'hffd; 
        10'b1010000000: data <= 12'hffa; 
        10'b1010000001: data <= 12'hffc; 
        10'b1010000010: data <= 12'hfff; 
        10'b1010000011: data <= 12'h000; 
        10'b1010000100: data <= 12'hfff; 
        10'b1010000101: data <= 12'hffd; 
        10'b1010000110: data <= 12'hffd; 
        10'b1010000111: data <= 12'h003; 
        10'b1010001000: data <= 12'h009; 
        10'b1010001001: data <= 12'h00e; 
        10'b1010001010: data <= 12'h00a; 
        10'b1010001011: data <= 12'h00b; 
        10'b1010001100: data <= 12'h003; 
        10'b1010001101: data <= 12'h007; 
        10'b1010001110: data <= 12'h004; 
        10'b1010001111: data <= 12'h000; 
        10'b1010010000: data <= 12'hffd; 
        10'b1010010001: data <= 12'h001; 
        10'b1010010010: data <= 12'h001; 
        10'b1010010011: data <= 12'h003; 
        10'b1010010100: data <= 12'h003; 
        10'b1010010101: data <= 12'h005; 
        10'b1010010110: data <= 12'h008; 
        10'b1010010111: data <= 12'hfff; 
        10'b1010011000: data <= 12'hffa; 
        10'b1010011001: data <= 12'hffa; 
        10'b1010011010: data <= 12'hffd; 
        10'b1010011011: data <= 12'hffc; 
        10'b1010011100: data <= 12'h000; 
        10'b1010011101: data <= 12'hfff; 
        10'b1010011110: data <= 12'hffc; 
        10'b1010011111: data <= 12'hffd; 
        10'b1010100000: data <= 12'hffd; 
        10'b1010100001: data <= 12'h000; 
        10'b1010100010: data <= 12'h000; 
        10'b1010100011: data <= 12'h000; 
        10'b1010100100: data <= 12'h006; 
        10'b1010100101: data <= 12'h009; 
        10'b1010100110: data <= 12'h00b; 
        10'b1010100111: data <= 12'h00d; 
        10'b1010101000: data <= 12'h00d; 
        10'b1010101001: data <= 12'h00b; 
        10'b1010101010: data <= 12'h010; 
        10'b1010101011: data <= 12'h011; 
        10'b1010101100: data <= 12'h011; 
        10'b1010101101: data <= 12'h00d; 
        10'b1010101110: data <= 12'h00c; 
        10'b1010101111: data <= 12'h009; 
        10'b1010110000: data <= 12'h008; 
        10'b1010110001: data <= 12'hfff; 
        10'b1010110010: data <= 12'hff9; 
        10'b1010110011: data <= 12'hff7; 
        10'b1010110100: data <= 12'hff8; 
        10'b1010110101: data <= 12'hffb; 
        10'b1010110110: data <= 12'hffb; 
        10'b1010110111: data <= 12'hfff; 
        10'b1010111000: data <= 12'hffe; 
        10'b1010111001: data <= 12'h000; 
        10'b1010111010: data <= 12'hffe; 
        10'b1010111011: data <= 12'h000; 
        10'b1010111100: data <= 12'h000; 
        10'b1010111101: data <= 12'hffc; 
        10'b1010111110: data <= 12'h000; 
        10'b1010111111: data <= 12'h001; 
        10'b1011000000: data <= 12'hfff; 
        10'b1011000001: data <= 12'h004; 
        10'b1011000010: data <= 12'h005; 
        10'b1011000011: data <= 12'h003; 
        10'b1011000100: data <= 12'h007; 
        10'b1011000101: data <= 12'h007; 
        10'b1011000110: data <= 12'h00e; 
        10'b1011000111: data <= 12'h010; 
        10'b1011001000: data <= 12'h011; 
        10'b1011001001: data <= 12'h00d; 
        10'b1011001010: data <= 12'h00a; 
        10'b1011001011: data <= 12'h004; 
        10'b1011001100: data <= 12'hffe; 
        10'b1011001101: data <= 12'hffa; 
        10'b1011001110: data <= 12'hffa; 
        10'b1011001111: data <= 12'hffb; 
        10'b1011010000: data <= 12'hffb; 
        10'b1011010001: data <= 12'hffe; 
        10'b1011010010: data <= 12'hffe; 
        10'b1011010011: data <= 12'h000; 
        10'b1011010100: data <= 12'hffd; 
        10'b1011010101: data <= 12'h000; 
        10'b1011010110: data <= 12'hffc; 
        10'b1011010111: data <= 12'hfff; 
        10'b1011011000: data <= 12'hffd; 
        10'b1011011001: data <= 12'hffc; 
        10'b1011011010: data <= 12'hffc; 
        10'b1011011011: data <= 12'hfff; 
        10'b1011011100: data <= 12'hfff; 
        10'b1011011101: data <= 12'hffd; 
        10'b1011011110: data <= 12'hffd; 
        10'b1011011111: data <= 12'hfff; 
        10'b1011100000: data <= 12'hfff; 
        10'b1011100001: data <= 12'hfff; 
        10'b1011100010: data <= 12'hffe; 
        10'b1011100011: data <= 12'hffe; 
        10'b1011100100: data <= 12'hffe; 
        10'b1011100101: data <= 12'hfff; 
        10'b1011100110: data <= 12'hffe; 
        10'b1011100111: data <= 12'hffc; 
        10'b1011101000: data <= 12'hffd; 
        10'b1011101001: data <= 12'hfff; 
        10'b1011101010: data <= 12'hffe; 
        10'b1011101011: data <= 12'hfff; 
        10'b1011101100: data <= 12'hffc; 
        10'b1011101101: data <= 12'hffc; 
        10'b1011101110: data <= 12'hfff; 
        10'b1011101111: data <= 12'hffe; 
        10'b1011110000: data <= 12'h000; 
        10'b1011110001: data <= 12'hffd; 
        10'b1011110010: data <= 12'h000; 
        10'b1011110011: data <= 12'h000; 
        10'b1011110100: data <= 12'hffe; 
        10'b1011110101: data <= 12'hffd; 
        10'b1011110110: data <= 12'hfff; 
        10'b1011110111: data <= 12'hffc; 
        10'b1011111000: data <= 12'h000; 
        10'b1011111001: data <= 12'hfff; 
        10'b1011111010: data <= 12'h000; 
        10'b1011111011: data <= 12'hfff; 
        10'b1011111100: data <= 12'hfff; 
        10'b1011111101: data <= 12'hffc; 
        10'b1011111110: data <= 12'hffd; 
        10'b1011111111: data <= 12'hfff; 
        10'b1100000000: data <= 12'hffd; 
        10'b1100000001: data <= 12'hfff; 
        10'b1100000010: data <= 12'hffe; 
        10'b1100000011: data <= 12'hfff; 
        10'b1100000100: data <= 12'hffe; 
        10'b1100000101: data <= 12'h000; 
        10'b1100000110: data <= 12'hffc; 
        10'b1100000111: data <= 12'hffd; 
        10'b1100001000: data <= 12'h000; 
        10'b1100001001: data <= 12'hfff; 
        10'b1100001010: data <= 12'hffd; 
        10'b1100001011: data <= 12'hfff; 
        10'b1100001100: data <= 12'hffc; 
        10'b1100001101: data <= 12'hffc; 
        10'b1100001110: data <= 12'h000; 
        10'b1100001111: data <= 12'hffe; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 7) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 13'h1ffd; 
        10'b0000000001: data <= 13'h1ffa; 
        10'b0000000010: data <= 13'h0000; 
        10'b0000000011: data <= 13'h0000; 
        10'b0000000100: data <= 13'h0001; 
        10'b0000000101: data <= 13'h1fff; 
        10'b0000000110: data <= 13'h1ffe; 
        10'b0000000111: data <= 13'h0001; 
        10'b0000001000: data <= 13'h1ffb; 
        10'b0000001001: data <= 13'h0000; 
        10'b0000001010: data <= 13'h0000; 
        10'b0000001011: data <= 13'h1ffc; 
        10'b0000001100: data <= 13'h1ffc; 
        10'b0000001101: data <= 13'h1ffb; 
        10'b0000001110: data <= 13'h1ffc; 
        10'b0000001111: data <= 13'h1ffc; 
        10'b0000010000: data <= 13'h0000; 
        10'b0000010001: data <= 13'h0000; 
        10'b0000010010: data <= 13'h1ffa; 
        10'b0000010011: data <= 13'h0001; 
        10'b0000010100: data <= 13'h1ffe; 
        10'b0000010101: data <= 13'h1ffe; 
        10'b0000010110: data <= 13'h1ff8; 
        10'b0000010111: data <= 13'h0000; 
        10'b0000011000: data <= 13'h0000; 
        10'b0000011001: data <= 13'h1ff8; 
        10'b0000011010: data <= 13'h1ffc; 
        10'b0000011011: data <= 13'h0000; 
        10'b0000011100: data <= 13'h1ffa; 
        10'b0000011101: data <= 13'h1ffc; 
        10'b0000011110: data <= 13'h1ffa; 
        10'b0000011111: data <= 13'h1ffe; 
        10'b0000100000: data <= 13'h1ff9; 
        10'b0000100001: data <= 13'h1ffd; 
        10'b0000100010: data <= 13'h0001; 
        10'b0000100011: data <= 13'h0000; 
        10'b0000100100: data <= 13'h1ff8; 
        10'b0000100101: data <= 13'h1ff8; 
        10'b0000100110: data <= 13'h1ff9; 
        10'b0000100111: data <= 13'h1ffe; 
        10'b0000101000: data <= 13'h1ffe; 
        10'b0000101001: data <= 13'h1ffc; 
        10'b0000101010: data <= 13'h1ffc; 
        10'b0000101011: data <= 13'h1ffa; 
        10'b0000101100: data <= 13'h0001; 
        10'b0000101101: data <= 13'h1ffa; 
        10'b0000101110: data <= 13'h1fff; 
        10'b0000101111: data <= 13'h1ffb; 
        10'b0000110000: data <= 13'h1ffb; 
        10'b0000110001: data <= 13'h1ff8; 
        10'b0000110010: data <= 13'h1ffd; 
        10'b0000110011: data <= 13'h1fff; 
        10'b0000110100: data <= 13'h1ff9; 
        10'b0000110101: data <= 13'h0000; 
        10'b0000110110: data <= 13'h1ffd; 
        10'b0000110111: data <= 13'h1ff9; 
        10'b0000111000: data <= 13'h1ffa; 
        10'b0000111001: data <= 13'h1ffd; 
        10'b0000111010: data <= 13'h1ffd; 
        10'b0000111011: data <= 13'h1ffa; 
        10'b0000111100: data <= 13'h1ffe; 
        10'b0000111101: data <= 13'h1fff; 
        10'b0000111110: data <= 13'h1ffb; 
        10'b0000111111: data <= 13'h1fff; 
        10'b0001000000: data <= 13'h1fff; 
        10'b0001000001: data <= 13'h1ffc; 
        10'b0001000010: data <= 13'h1ff9; 
        10'b0001000011: data <= 13'h1ff9; 
        10'b0001000100: data <= 13'h1ff8; 
        10'b0001000101: data <= 13'h1ff9; 
        10'b0001000110: data <= 13'h1ffc; 
        10'b0001000111: data <= 13'h1ffb; 
        10'b0001001000: data <= 13'h1ffb; 
        10'b0001001001: data <= 13'h1ffa; 
        10'b0001001010: data <= 13'h1fff; 
        10'b0001001011: data <= 13'h0000; 
        10'b0001001100: data <= 13'h1ffc; 
        10'b0001001101: data <= 13'h1ffa; 
        10'b0001001110: data <= 13'h0001; 
        10'b0001001111: data <= 13'h1fff; 
        10'b0001010000: data <= 13'h0000; 
        10'b0001010001: data <= 13'h1ffb; 
        10'b0001010010: data <= 13'h1ff8; 
        10'b0001010011: data <= 13'h1ffc; 
        10'b0001010100: data <= 13'h0001; 
        10'b0001010101: data <= 13'h1fff; 
        10'b0001010110: data <= 13'h1ffc; 
        10'b0001010111: data <= 13'h1fff; 
        10'b0001011000: data <= 13'h1ffe; 
        10'b0001011001: data <= 13'h0000; 
        10'b0001011010: data <= 13'h1ffe; 
        10'b0001011011: data <= 13'h0000; 
        10'b0001011100: data <= 13'h1fff; 
        10'b0001011101: data <= 13'h1ffd; 
        10'b0001011110: data <= 13'h0003; 
        10'b0001011111: data <= 13'h0009; 
        10'b0001100000: data <= 13'h0014; 
        10'b0001100001: data <= 13'h0010; 
        10'b0001100010: data <= 13'h0011; 
        10'b0001100011: data <= 13'h0012; 
        10'b0001100100: data <= 13'h000d; 
        10'b0001100101: data <= 13'h000e; 
        10'b0001100110: data <= 13'h000b; 
        10'b0001100111: data <= 13'h0001; 
        10'b0001101000: data <= 13'h1fff; 
        10'b0001101001: data <= 13'h1ff2; 
        10'b0001101010: data <= 13'h1ff8; 
        10'b0001101011: data <= 13'h1fff; 
        10'b0001101100: data <= 13'h0000; 
        10'b0001101101: data <= 13'h1ffa; 
        10'b0001101110: data <= 13'h1ffd; 
        10'b0001101111: data <= 13'h1ffb; 
        10'b0001110000: data <= 13'h1ffd; 
        10'b0001110001: data <= 13'h0000; 
        10'b0001110010: data <= 13'h1ffe; 
        10'b0001110011: data <= 13'h0000; 
        10'b0001110100: data <= 13'h0003; 
        10'b0001110101: data <= 13'h0000; 
        10'b0001110110: data <= 13'h000b; 
        10'b0001110111: data <= 13'h000a; 
        10'b0001111000: data <= 13'h001a; 
        10'b0001111001: data <= 13'h0017; 
        10'b0001111010: data <= 13'h001c; 
        10'b0001111011: data <= 13'h0022; 
        10'b0001111100: data <= 13'h0027; 
        10'b0001111101: data <= 13'h002a; 
        10'b0001111110: data <= 13'h0026; 
        10'b0001111111: data <= 13'h001c; 
        10'b0010000000: data <= 13'h0010; 
        10'b0010000001: data <= 13'h000d; 
        10'b0010000010: data <= 13'h0014; 
        10'b0010000011: data <= 13'h0003; 
        10'b0010000100: data <= 13'h1ff2; 
        10'b0010000101: data <= 13'h1fea; 
        10'b0010000110: data <= 13'h1fed; 
        10'b0010000111: data <= 13'h1fee; 
        10'b0010001000: data <= 13'h1ffe; 
        10'b0010001001: data <= 13'h1ffd; 
        10'b0010001010: data <= 13'h1ffb; 
        10'b0010001011: data <= 13'h1fff; 
        10'b0010001100: data <= 13'h1ff9; 
        10'b0010001101: data <= 13'h1ff8; 
        10'b0010001110: data <= 13'h1ffa; 
        10'b0010001111: data <= 13'h1ffa; 
        10'b0010010000: data <= 13'h0001; 
        10'b0010010001: data <= 13'h000c; 
        10'b0010010010: data <= 13'h0016; 
        10'b0010010011: data <= 13'h0011; 
        10'b0010010100: data <= 13'h0014; 
        10'b0010010101: data <= 13'h0012; 
        10'b0010010110: data <= 13'h0010; 
        10'b0010010111: data <= 13'h0015; 
        10'b0010011000: data <= 13'h0015; 
        10'b0010011001: data <= 13'h0019; 
        10'b0010011010: data <= 13'h0004; 
        10'b0010011011: data <= 13'h0011; 
        10'b0010011100: data <= 13'h0013; 
        10'b0010011101: data <= 13'h1fff; 
        10'b0010011110: data <= 13'h1fff; 
        10'b0010011111: data <= 13'h1ff7; 
        10'b0010100000: data <= 13'h1ff4; 
        10'b0010100001: data <= 13'h1fe6; 
        10'b0010100010: data <= 13'h1fdf; 
        10'b0010100011: data <= 13'h1fe4; 
        10'b0010100100: data <= 13'h1ff8; 
        10'b0010100101: data <= 13'h0000; 
        10'b0010100110: data <= 13'h1ffa; 
        10'b0010100111: data <= 13'h1ffd; 
        10'b0010101000: data <= 13'h1ffa; 
        10'b0010101001: data <= 13'h1ffb; 
        10'b0010101010: data <= 13'h1ffb; 
        10'b0010101011: data <= 13'h0003; 
        10'b0010101100: data <= 13'h000f; 
        10'b0010101101: data <= 13'h001c; 
        10'b0010101110: data <= 13'h0015; 
        10'b0010101111: data <= 13'h0010; 
        10'b0010110000: data <= 13'h0018; 
        10'b0010110001: data <= 13'h0014; 
        10'b0010110010: data <= 13'h0012; 
        10'b0010110011: data <= 13'h0011; 
        10'b0010110100: data <= 13'h0017; 
        10'b0010110101: data <= 13'h0020; 
        10'b0010110110: data <= 13'h0017; 
        10'b0010110111: data <= 13'h0008; 
        10'b0010111000: data <= 13'h0015; 
        10'b0010111001: data <= 13'h0014; 
        10'b0010111010: data <= 13'h0013; 
        10'b0010111011: data <= 13'h1ff8; 
        10'b0010111100: data <= 13'h0008; 
        10'b0010111101: data <= 13'h1ff8; 
        10'b0010111110: data <= 13'h1fe3; 
        10'b0010111111: data <= 13'h1fe3; 
        10'b0011000000: data <= 13'h1fef; 
        10'b0011000001: data <= 13'h1ffc; 
        10'b0011000010: data <= 13'h1fff; 
        10'b0011000011: data <= 13'h1ffd; 
        10'b0011000100: data <= 13'h0000; 
        10'b0011000101: data <= 13'h1fff; 
        10'b0011000110: data <= 13'h0002; 
        10'b0011000111: data <= 13'h000c; 
        10'b0011001000: data <= 13'h0020; 
        10'b0011001001: data <= 13'h0020; 
        10'b0011001010: data <= 13'h0017; 
        10'b0011001011: data <= 13'h0006; 
        10'b0011001100: data <= 13'h0007; 
        10'b0011001101: data <= 13'h000e; 
        10'b0011001110: data <= 13'h0004; 
        10'b0011001111: data <= 13'h0007; 
        10'b0011010000: data <= 13'h0013; 
        10'b0011010001: data <= 13'h0012; 
        10'b0011010010: data <= 13'h001e; 
        10'b0011010011: data <= 13'h0012; 
        10'b0011010100: data <= 13'h0005; 
        10'b0011010101: data <= 13'h000f; 
        10'b0011010110: data <= 13'h000c; 
        10'b0011010111: data <= 13'h000e; 
        10'b0011011000: data <= 13'h000e; 
        10'b0011011001: data <= 13'h0002; 
        10'b0011011010: data <= 13'h1ff2; 
        10'b0011011011: data <= 13'h1fe0; 
        10'b0011011100: data <= 13'h1fe9; 
        10'b0011011101: data <= 13'h1ffa; 
        10'b0011011110: data <= 13'h1ff8; 
        10'b0011011111: data <= 13'h1ffc; 
        10'b0011100000: data <= 13'h1ffd; 
        10'b0011100001: data <= 13'h1ffb; 
        10'b0011100010: data <= 13'h0001; 
        10'b0011100011: data <= 13'h000c; 
        10'b0011100100: data <= 13'h001b; 
        10'b0011100101: data <= 13'h0019; 
        10'b0011100110: data <= 13'h0013; 
        10'b0011100111: data <= 13'h0008; 
        10'b0011101000: data <= 13'h000d; 
        10'b0011101001: data <= 13'h0006; 
        10'b0011101010: data <= 13'h0010; 
        10'b0011101011: data <= 13'h0005; 
        10'b0011101100: data <= 13'h0004; 
        10'b0011101101: data <= 13'h0008; 
        10'b0011101110: data <= 13'h0020; 
        10'b0011101111: data <= 13'h001b; 
        10'b0011110000: data <= 13'h0006; 
        10'b0011110001: data <= 13'h000f; 
        10'b0011110010: data <= 13'h0016; 
        10'b0011110011: data <= 13'h000e; 
        10'b0011110100: data <= 13'h0015; 
        10'b0011110101: data <= 13'h000b; 
        10'b0011110110: data <= 13'h1ffb; 
        10'b0011110111: data <= 13'h1fe2; 
        10'b0011111000: data <= 13'h1fea; 
        10'b0011111001: data <= 13'h1ff8; 
        10'b0011111010: data <= 13'h1ff9; 
        10'b0011111011: data <= 13'h1ffb; 
        10'b0011111100: data <= 13'h1ffc; 
        10'b0011111101: data <= 13'h1ff8; 
        10'b0011111110: data <= 13'h1ffe; 
        10'b0011111111: data <= 13'h0005; 
        10'b0100000000: data <= 13'h000e; 
        10'b0100000001: data <= 13'h0012; 
        10'b0100000010: data <= 13'h000f; 
        10'b0100000011: data <= 13'h0004; 
        10'b0100000100: data <= 13'h1ffe; 
        10'b0100000101: data <= 13'h1ff2; 
        10'b0100000110: data <= 13'h1fe5; 
        10'b0100000111: data <= 13'h1fce; 
        10'b0100001000: data <= 13'h1fd8; 
        10'b0100001001: data <= 13'h1ffb; 
        10'b0100001010: data <= 13'h0027; 
        10'b0100001011: data <= 13'h003b; 
        10'b0100001100: data <= 13'h0022; 
        10'b0100001101: data <= 13'h0014; 
        10'b0100001110: data <= 13'h0016; 
        10'b0100001111: data <= 13'h0014; 
        10'b0100010000: data <= 13'h001e; 
        10'b0100010001: data <= 13'h0013; 
        10'b0100010010: data <= 13'h1ffa; 
        10'b0100010011: data <= 13'h1fe2; 
        10'b0100010100: data <= 13'h1ff1; 
        10'b0100010101: data <= 13'h1ff8; 
        10'b0100010110: data <= 13'h1ffa; 
        10'b0100010111: data <= 13'h1ffb; 
        10'b0100011000: data <= 13'h1fff; 
        10'b0100011001: data <= 13'h1fff; 
        10'b0100011010: data <= 13'h0000; 
        10'b0100011011: data <= 13'h0007; 
        10'b0100011100: data <= 13'h0007; 
        10'b0100011101: data <= 13'h0003; 
        10'b0100011110: data <= 13'h1ff7; 
        10'b0100011111: data <= 13'h1fea; 
        10'b0100100000: data <= 13'h1fd8; 
        10'b0100100001: data <= 13'h1fc7; 
        10'b0100100010: data <= 13'h1fba; 
        10'b0100100011: data <= 13'h1fb8; 
        10'b0100100100: data <= 13'h1fcb; 
        10'b0100100101: data <= 13'h1ff3; 
        10'b0100100110: data <= 13'h0020; 
        10'b0100100111: data <= 13'h0025; 
        10'b0100101000: data <= 13'h001f; 
        10'b0100101001: data <= 13'h001d; 
        10'b0100101010: data <= 13'h0012; 
        10'b0100101011: data <= 13'h001f; 
        10'b0100101100: data <= 13'h001d; 
        10'b0100101101: data <= 13'h000c; 
        10'b0100101110: data <= 13'h1ff6; 
        10'b0100101111: data <= 13'h1fed; 
        10'b0100110000: data <= 13'h1ff9; 
        10'b0100110001: data <= 13'h1ff8; 
        10'b0100110010: data <= 13'h1ffd; 
        10'b0100110011: data <= 13'h1fff; 
        10'b0100110100: data <= 13'h0001; 
        10'b0100110101: data <= 13'h1fff; 
        10'b0100110110: data <= 13'h1ff9; 
        10'b0100110111: data <= 13'h0007; 
        10'b0100111000: data <= 13'h1ffc; 
        10'b0100111001: data <= 13'h1fea; 
        10'b0100111010: data <= 13'h1fde; 
        10'b0100111011: data <= 13'h1fce; 
        10'b0100111100: data <= 13'h1fc2; 
        10'b0100111101: data <= 13'h1fca; 
        10'b0100111110: data <= 13'h1fd7; 
        10'b0100111111: data <= 13'h1fed; 
        10'b0101000000: data <= 13'h1ff6; 
        10'b0101000001: data <= 13'h000d; 
        10'b0101000010: data <= 13'h0015; 
        10'b0101000011: data <= 13'h0015; 
        10'b0101000100: data <= 13'h000a; 
        10'b0101000101: data <= 13'h0016; 
        10'b0101000110: data <= 13'h001b; 
        10'b0101000111: data <= 13'h001b; 
        10'b0101001000: data <= 13'h0017; 
        10'b0101001001: data <= 13'h0000; 
        10'b0101001010: data <= 13'h1ff6; 
        10'b0101001011: data <= 13'h1ff7; 
        10'b0101001100: data <= 13'h1ff8; 
        10'b0101001101: data <= 13'h1ffc; 
        10'b0101001110: data <= 13'h1ffa; 
        10'b0101001111: data <= 13'h1ff9; 
        10'b0101010000: data <= 13'h0000; 
        10'b0101010001: data <= 13'h1ffb; 
        10'b0101010010: data <= 13'h1fff; 
        10'b0101010011: data <= 13'h0000; 
        10'b0101010100: data <= 13'h1ff8; 
        10'b0101010101: data <= 13'h1fe9; 
        10'b0101010110: data <= 13'h1fd9; 
        10'b0101010111: data <= 13'h1fcf; 
        10'b0101011000: data <= 13'h1fd3; 
        10'b0101011001: data <= 13'h1fe8; 
        10'b0101011010: data <= 13'h0000; 
        10'b0101011011: data <= 13'h0004; 
        10'b0101011100: data <= 13'h0006; 
        10'b0101011101: data <= 13'h000e; 
        10'b0101011110: data <= 13'h0023; 
        10'b0101011111: data <= 13'h0012; 
        10'b0101100000: data <= 13'h000c; 
        10'b0101100001: data <= 13'h0012; 
        10'b0101100010: data <= 13'h000e; 
        10'b0101100011: data <= 13'h1fff; 
        10'b0101100100: data <= 13'h1fee; 
        10'b0101100101: data <= 13'h1fe7; 
        10'b0101100110: data <= 13'h1fe6; 
        10'b0101100111: data <= 13'h1fef; 
        10'b0101101000: data <= 13'h1ffd; 
        10'b0101101001: data <= 13'h1ffb; 
        10'b0101101010: data <= 13'h1ffd; 
        10'b0101101011: data <= 13'h1ffe; 
        10'b0101101100: data <= 13'h1ffc; 
        10'b0101101101: data <= 13'h1ffb; 
        10'b0101101110: data <= 13'h1ffd; 
        10'b0101101111: data <= 13'h1ffe; 
        10'b0101110000: data <= 13'h1ff6; 
        10'b0101110001: data <= 13'h1ff1; 
        10'b0101110010: data <= 13'h1fe0; 
        10'b0101110011: data <= 13'h1fdb; 
        10'b0101110100: data <= 13'h1fe7; 
        10'b0101110101: data <= 13'h1ffb; 
        10'b0101110110: data <= 13'h1ff8; 
        10'b0101110111: data <= 13'h1feb; 
        10'b0101111000: data <= 13'h0002; 
        10'b0101111001: data <= 13'h001e; 
        10'b0101111010: data <= 13'h001f; 
        10'b0101111011: data <= 13'h0006; 
        10'b0101111100: data <= 13'h000e; 
        10'b0101111101: data <= 13'h000f; 
        10'b0101111110: data <= 13'h0008; 
        10'b0101111111: data <= 13'h1ff6; 
        10'b0110000000: data <= 13'h1fe4; 
        10'b0110000001: data <= 13'h1fe4; 
        10'b0110000010: data <= 13'h1fea; 
        10'b0110000011: data <= 13'h1ff0; 
        10'b0110000100: data <= 13'h1ff7; 
        10'b0110000101: data <= 13'h0000; 
        10'b0110000110: data <= 13'h1ffe; 
        10'b0110000111: data <= 13'h1ffb; 
        10'b0110001000: data <= 13'h0001; 
        10'b0110001001: data <= 13'h1ffa; 
        10'b0110001010: data <= 13'h1ffc; 
        10'b0110001011: data <= 13'h1ffd; 
        10'b0110001100: data <= 13'h1ffe; 
        10'b0110001101: data <= 13'h1ff3; 
        10'b0110001110: data <= 13'h1fe3; 
        10'b0110001111: data <= 13'h1fe6; 
        10'b0110010000: data <= 13'h1fee; 
        10'b0110010001: data <= 13'h1ffe; 
        10'b0110010010: data <= 13'h1fed; 
        10'b0110010011: data <= 13'h1fec; 
        10'b0110010100: data <= 13'h0006; 
        10'b0110010101: data <= 13'h000f; 
        10'b0110010110: data <= 13'h0010; 
        10'b0110010111: data <= 13'h1ffe; 
        10'b0110011000: data <= 13'h1ffa; 
        10'b0110011001: data <= 13'h1ffb; 
        10'b0110011010: data <= 13'h0002; 
        10'b0110011011: data <= 13'h1ff4; 
        10'b0110011100: data <= 13'h1fef; 
        10'b0110011101: data <= 13'h1ff8; 
        10'b0110011110: data <= 13'h1ff5; 
        10'b0110011111: data <= 13'h1ff8; 
        10'b0110100000: data <= 13'h1ff6; 
        10'b0110100001: data <= 13'h1ff7; 
        10'b0110100010: data <= 13'h0000; 
        10'b0110100011: data <= 13'h0000; 
        10'b0110100100: data <= 13'h0001; 
        10'b0110100101: data <= 13'h1ffa; 
        10'b0110100110: data <= 13'h0001; 
        10'b0110100111: data <= 13'h0002; 
        10'b0110101000: data <= 13'h1ffd; 
        10'b0110101001: data <= 13'h1ff2; 
        10'b0110101010: data <= 13'h1fe5; 
        10'b0110101011: data <= 13'h1fe3; 
        10'b0110101100: data <= 13'h1fea; 
        10'b0110101101: data <= 13'h1ff3; 
        10'b0110101110: data <= 13'h1ff2; 
        10'b0110101111: data <= 13'h1ffb; 
        10'b0110110000: data <= 13'h0006; 
        10'b0110110001: data <= 13'h0018; 
        10'b0110110010: data <= 13'h000e; 
        10'b0110110011: data <= 13'h1fff; 
        10'b0110110100: data <= 13'h1fec; 
        10'b0110110101: data <= 13'h1ffa; 
        10'b0110110110: data <= 13'h1ffe; 
        10'b0110110111: data <= 13'h0005; 
        10'b0110111000: data <= 13'h000c; 
        10'b0110111001: data <= 13'h000c; 
        10'b0110111010: data <= 13'h0004; 
        10'b0110111011: data <= 13'h0002; 
        10'b0110111100: data <= 13'h1ff8; 
        10'b0110111101: data <= 13'h1ffe; 
        10'b0110111110: data <= 13'h1ffe; 
        10'b0110111111: data <= 13'h1ffa; 
        10'b0111000000: data <= 13'h1ffe; 
        10'b0111000001: data <= 13'h1fff; 
        10'b0111000010: data <= 13'h0006; 
        10'b0111000011: data <= 13'h0001; 
        10'b0111000100: data <= 13'h0004; 
        10'b0111000101: data <= 13'h1ff9; 
        10'b0111000110: data <= 13'h1ff5; 
        10'b0111000111: data <= 13'h1fed; 
        10'b0111001000: data <= 13'h1fd7; 
        10'b0111001001: data <= 13'h1fd4; 
        10'b0111001010: data <= 13'h1fd9; 
        10'b0111001011: data <= 13'h1ff6; 
        10'b0111001100: data <= 13'h000c; 
        10'b0111001101: data <= 13'h001e; 
        10'b0111001110: data <= 13'h1ffd; 
        10'b0111001111: data <= 13'h1fea; 
        10'b0111010000: data <= 13'h1fe9; 
        10'b0111010001: data <= 13'h1ff8; 
        10'b0111010010: data <= 13'h000a; 
        10'b0111010011: data <= 13'h0019; 
        10'b0111010100: data <= 13'h0012; 
        10'b0111010101: data <= 13'h0017; 
        10'b0111010110: data <= 13'h0016; 
        10'b0111010111: data <= 13'h000a; 
        10'b0111011000: data <= 13'h1ffd; 
        10'b0111011001: data <= 13'h1ffe; 
        10'b0111011010: data <= 13'h0000; 
        10'b0111011011: data <= 13'h1fff; 
        10'b0111011100: data <= 13'h1fff; 
        10'b0111011101: data <= 13'h0001; 
        10'b0111011110: data <= 13'h0000; 
        10'b0111011111: data <= 13'h000e; 
        10'b0111100000: data <= 13'h0008; 
        10'b0111100001: data <= 13'h0002; 
        10'b0111100010: data <= 13'h1ff9; 
        10'b0111100011: data <= 13'h1fe7; 
        10'b0111100100: data <= 13'h1fd3; 
        10'b0111100101: data <= 13'h1fb9; 
        10'b0111100110: data <= 13'h1fa8; 
        10'b0111100111: data <= 13'h1faf; 
        10'b0111101000: data <= 13'h1fc3; 
        10'b0111101001: data <= 13'h1fdd; 
        10'b0111101010: data <= 13'h1fe0; 
        10'b0111101011: data <= 13'h1fe3; 
        10'b0111101100: data <= 13'h1fff; 
        10'b0111101101: data <= 13'h0009; 
        10'b0111101110: data <= 13'h0010; 
        10'b0111101111: data <= 13'h001a; 
        10'b0111110000: data <= 13'h0005; 
        10'b0111110001: data <= 13'h001f; 
        10'b0111110010: data <= 13'h001f; 
        10'b0111110011: data <= 13'h0009; 
        10'b0111110100: data <= 13'h1ffb; 
        10'b0111110101: data <= 13'h1ff9; 
        10'b0111110110: data <= 13'h1ffa; 
        10'b0111110111: data <= 13'h1ffa; 
        10'b0111111000: data <= 13'h1ffd; 
        10'b0111111001: data <= 13'h1ffd; 
        10'b0111111010: data <= 13'h0003; 
        10'b0111111011: data <= 13'h0015; 
        10'b0111111100: data <= 13'h000f; 
        10'b0111111101: data <= 13'h0009; 
        10'b0111111110: data <= 13'h0005; 
        10'b0111111111: data <= 13'h1ffb; 
        10'b1000000000: data <= 13'h1ff0; 
        10'b1000000001: data <= 13'h1fcc; 
        10'b1000000010: data <= 13'h1fb4; 
        10'b1000000011: data <= 13'h1fb8; 
        10'b1000000100: data <= 13'h1fa9; 
        10'b1000000101: data <= 13'h1fb9; 
        10'b1000000110: data <= 13'h1fd3; 
        10'b1000000111: data <= 13'h1ff6; 
        10'b1000001000: data <= 13'h0012; 
        10'b1000001001: data <= 13'h0019; 
        10'b1000001010: data <= 13'h001a; 
        10'b1000001011: data <= 13'h001a; 
        10'b1000001100: data <= 13'h0012; 
        10'b1000001101: data <= 13'h0024; 
        10'b1000001110: data <= 13'h0022; 
        10'b1000001111: data <= 13'h000d; 
        10'b1000010000: data <= 13'h1ff4; 
        10'b1000010001: data <= 13'h1ff8; 
        10'b1000010010: data <= 13'h1ffa; 
        10'b1000010011: data <= 13'h1fff; 
        10'b1000010100: data <= 13'h1fff; 
        10'b1000010101: data <= 13'h1ffa; 
        10'b1000010110: data <= 13'h1ffc; 
        10'b1000010111: data <= 13'h001a; 
        10'b1000011000: data <= 13'h001a; 
        10'b1000011001: data <= 13'h001f; 
        10'b1000011010: data <= 13'h001b; 
        10'b1000011011: data <= 13'h000a; 
        10'b1000011100: data <= 13'h0003; 
        10'b1000011101: data <= 13'h1ff5; 
        10'b1000011110: data <= 13'h1ff8; 
        10'b1000011111: data <= 13'h1fe7; 
        10'b1000100000: data <= 13'h1fdc; 
        10'b1000100001: data <= 13'h1fda; 
        10'b1000100010: data <= 13'h1fe6; 
        10'b1000100011: data <= 13'h0009; 
        10'b1000100100: data <= 13'h0019; 
        10'b1000100101: data <= 13'h001f; 
        10'b1000100110: data <= 13'h0023; 
        10'b1000100111: data <= 13'h001f; 
        10'b1000101000: data <= 13'h001b; 
        10'b1000101001: data <= 13'h0020; 
        10'b1000101010: data <= 13'h000c; 
        10'b1000101011: data <= 13'h0001; 
        10'b1000101100: data <= 13'h1ff6; 
        10'b1000101101: data <= 13'h1ffe; 
        10'b1000101110: data <= 13'h1fff; 
        10'b1000101111: data <= 13'h1ffe; 
        10'b1000110000: data <= 13'h1fff; 
        10'b1000110001: data <= 13'h1ff8; 
        10'b1000110010: data <= 13'h0005; 
        10'b1000110011: data <= 13'h001c; 
        10'b1000110100: data <= 13'h0022; 
        10'b1000110101: data <= 13'h0025; 
        10'b1000110110: data <= 13'h0027; 
        10'b1000110111: data <= 13'h0014; 
        10'b1000111000: data <= 13'h0017; 
        10'b1000111001: data <= 13'h001a; 
        10'b1000111010: data <= 13'h000a; 
        10'b1000111011: data <= 13'h1ffd; 
        10'b1000111100: data <= 13'h1ff7; 
        10'b1000111101: data <= 13'h1ff2; 
        10'b1000111110: data <= 13'h0004; 
        10'b1000111111: data <= 13'h0007; 
        10'b1001000000: data <= 13'h000e; 
        10'b1001000001: data <= 13'h0019; 
        10'b1001000010: data <= 13'h001a; 
        10'b1001000011: data <= 13'h0012; 
        10'b1001000100: data <= 13'h001f; 
        10'b1001000101: data <= 13'h0011; 
        10'b1001000110: data <= 13'h1ffd; 
        10'b1001000111: data <= 13'h1ff9; 
        10'b1001001000: data <= 13'h1ff8; 
        10'b1001001001: data <= 13'h1ffe; 
        10'b1001001010: data <= 13'h1ffd; 
        10'b1001001011: data <= 13'h1ffd; 
        10'b1001001100: data <= 13'h1ffb; 
        10'b1001001101: data <= 13'h0000; 
        10'b1001001110: data <= 13'h1ffe; 
        10'b1001001111: data <= 13'h000e; 
        10'b1001010000: data <= 13'h0021; 
        10'b1001010001: data <= 13'h0021; 
        10'b1001010010: data <= 13'h001d; 
        10'b1001010011: data <= 13'h0010; 
        10'b1001010100: data <= 13'h0011; 
        10'b1001010101: data <= 13'h0006; 
        10'b1001010110: data <= 13'h1ffe; 
        10'b1001010111: data <= 13'h1ff8; 
        10'b1001011000: data <= 13'h0002; 
        10'b1001011001: data <= 13'h1fff; 
        10'b1001011010: data <= 13'h1ffe; 
        10'b1001011011: data <= 13'h1ffc; 
        10'b1001011100: data <= 13'h0008; 
        10'b1001011101: data <= 13'h0003; 
        10'b1001011110: data <= 13'h0010; 
        10'b1001011111: data <= 13'h0019; 
        10'b1001100000: data <= 13'h000f; 
        10'b1001100001: data <= 13'h0006; 
        10'b1001100010: data <= 13'h1ffa; 
        10'b1001100011: data <= 13'h1ff1; 
        10'b1001100100: data <= 13'h1ffb; 
        10'b1001100101: data <= 13'h1ffa; 
        10'b1001100110: data <= 13'h1ff8; 
        10'b1001100111: data <= 13'h1ff8; 
        10'b1001101000: data <= 13'h1ffd; 
        10'b1001101001: data <= 13'h1ffe; 
        10'b1001101010: data <= 13'h1ffe; 
        10'b1001101011: data <= 13'h0009; 
        10'b1001101100: data <= 13'h0011; 
        10'b1001101101: data <= 13'h0017; 
        10'b1001101110: data <= 13'h0014; 
        10'b1001101111: data <= 13'h000b; 
        10'b1001110000: data <= 13'h0001; 
        10'b1001110001: data <= 13'h0008; 
        10'b1001110010: data <= 13'h000a; 
        10'b1001110011: data <= 13'h000c; 
        10'b1001110100: data <= 13'h0003; 
        10'b1001110101: data <= 13'h1ffc; 
        10'b1001110110: data <= 13'h1ffb; 
        10'b1001110111: data <= 13'h1ff9; 
        10'b1001111000: data <= 13'h0005; 
        10'b1001111001: data <= 13'h0004; 
        10'b1001111010: data <= 13'h0004; 
        10'b1001111011: data <= 13'h0012; 
        10'b1001111100: data <= 13'h0009; 
        10'b1001111101: data <= 13'h1ffd; 
        10'b1001111110: data <= 13'h1ffc; 
        10'b1001111111: data <= 13'h1ffb; 
        10'b1010000000: data <= 13'h1ff5; 
        10'b1010000001: data <= 13'h1ff8; 
        10'b1010000010: data <= 13'h1ffe; 
        10'b1010000011: data <= 13'h0000; 
        10'b1010000100: data <= 13'h1ffe; 
        10'b1010000101: data <= 13'h1ffa; 
        10'b1010000110: data <= 13'h1ffb; 
        10'b1010000111: data <= 13'h0006; 
        10'b1010001000: data <= 13'h0012; 
        10'b1010001001: data <= 13'h001b; 
        10'b1010001010: data <= 13'h0014; 
        10'b1010001011: data <= 13'h0015; 
        10'b1010001100: data <= 13'h0005; 
        10'b1010001101: data <= 13'h000e; 
        10'b1010001110: data <= 13'h0009; 
        10'b1010001111: data <= 13'h0000; 
        10'b1010010000: data <= 13'h1ff9; 
        10'b1010010001: data <= 13'h0001; 
        10'b1010010010: data <= 13'h0003; 
        10'b1010010011: data <= 13'h0007; 
        10'b1010010100: data <= 13'h0005; 
        10'b1010010101: data <= 13'h000b; 
        10'b1010010110: data <= 13'h0011; 
        10'b1010010111: data <= 13'h1ffd; 
        10'b1010011000: data <= 13'h1ff5; 
        10'b1010011001: data <= 13'h1ff5; 
        10'b1010011010: data <= 13'h1ffa; 
        10'b1010011011: data <= 13'h1ff9; 
        10'b1010011100: data <= 13'h1fff; 
        10'b1010011101: data <= 13'h1ffe; 
        10'b1010011110: data <= 13'h1ff9; 
        10'b1010011111: data <= 13'h1ffa; 
        10'b1010100000: data <= 13'h1ffb; 
        10'b1010100001: data <= 13'h0001; 
        10'b1010100010: data <= 13'h0001; 
        10'b1010100011: data <= 13'h0000; 
        10'b1010100100: data <= 13'h000c; 
        10'b1010100101: data <= 13'h0013; 
        10'b1010100110: data <= 13'h0016; 
        10'b1010100111: data <= 13'h001a; 
        10'b1010101000: data <= 13'h001a; 
        10'b1010101001: data <= 13'h0016; 
        10'b1010101010: data <= 13'h0020; 
        10'b1010101011: data <= 13'h0021; 
        10'b1010101100: data <= 13'h0022; 
        10'b1010101101: data <= 13'h001b; 
        10'b1010101110: data <= 13'h0018; 
        10'b1010101111: data <= 13'h0012; 
        10'b1010110000: data <= 13'h0011; 
        10'b1010110001: data <= 13'h1fff; 
        10'b1010110010: data <= 13'h1ff2; 
        10'b1010110011: data <= 13'h1fed; 
        10'b1010110100: data <= 13'h1fef; 
        10'b1010110101: data <= 13'h1ff6; 
        10'b1010110110: data <= 13'h1ff6; 
        10'b1010110111: data <= 13'h1ffd; 
        10'b1010111000: data <= 13'h1ffb; 
        10'b1010111001: data <= 13'h0000; 
        10'b1010111010: data <= 13'h1ffb; 
        10'b1010111011: data <= 13'h0001; 
        10'b1010111100: data <= 13'h1fff; 
        10'b1010111101: data <= 13'h1ff8; 
        10'b1010111110: data <= 13'h0001; 
        10'b1010111111: data <= 13'h0001; 
        10'b1011000000: data <= 13'h1ffe; 
        10'b1011000001: data <= 13'h0007; 
        10'b1011000010: data <= 13'h000b; 
        10'b1011000011: data <= 13'h0006; 
        10'b1011000100: data <= 13'h000f; 
        10'b1011000101: data <= 13'h000f; 
        10'b1011000110: data <= 13'h001c; 
        10'b1011000111: data <= 13'h0020; 
        10'b1011001000: data <= 13'h0022; 
        10'b1011001001: data <= 13'h001b; 
        10'b1011001010: data <= 13'h0013; 
        10'b1011001011: data <= 13'h0008; 
        10'b1011001100: data <= 13'h1ffd; 
        10'b1011001101: data <= 13'h1ff4; 
        10'b1011001110: data <= 13'h1ff4; 
        10'b1011001111: data <= 13'h1ff6; 
        10'b1011010000: data <= 13'h1ff6; 
        10'b1011010001: data <= 13'h1ffb; 
        10'b1011010010: data <= 13'h1ffb; 
        10'b1011010011: data <= 13'h1fff; 
        10'b1011010100: data <= 13'h1ffa; 
        10'b1011010101: data <= 13'h0001; 
        10'b1011010110: data <= 13'h1ff8; 
        10'b1011010111: data <= 13'h1fff; 
        10'b1011011000: data <= 13'h1ffa; 
        10'b1011011001: data <= 13'h1ff8; 
        10'b1011011010: data <= 13'h1ff8; 
        10'b1011011011: data <= 13'h1ffe; 
        10'b1011011100: data <= 13'h1ffe; 
        10'b1011011101: data <= 13'h1ffb; 
        10'b1011011110: data <= 13'h1ffa; 
        10'b1011011111: data <= 13'h1ffe; 
        10'b1011100000: data <= 13'h1ffe; 
        10'b1011100001: data <= 13'h1ffd; 
        10'b1011100010: data <= 13'h1ffc; 
        10'b1011100011: data <= 13'h1ffd; 
        10'b1011100100: data <= 13'h1ffb; 
        10'b1011100101: data <= 13'h1ffe; 
        10'b1011100110: data <= 13'h1ffb; 
        10'b1011100111: data <= 13'h1ff7; 
        10'b1011101000: data <= 13'h1ffb; 
        10'b1011101001: data <= 13'h1ffd; 
        10'b1011101010: data <= 13'h1ffc; 
        10'b1011101011: data <= 13'h1ffe; 
        10'b1011101100: data <= 13'h1ff8; 
        10'b1011101101: data <= 13'h1ff8; 
        10'b1011101110: data <= 13'h1fff; 
        10'b1011101111: data <= 13'h1ffc; 
        10'b1011110000: data <= 13'h0000; 
        10'b1011110001: data <= 13'h1ffa; 
        10'b1011110010: data <= 13'h1fff; 
        10'b1011110011: data <= 13'h0001; 
        10'b1011110100: data <= 13'h1ffc; 
        10'b1011110101: data <= 13'h1ffa; 
        10'b1011110110: data <= 13'h1ffd; 
        10'b1011110111: data <= 13'h1ff8; 
        10'b1011111000: data <= 13'h0000; 
        10'b1011111001: data <= 13'h1ffe; 
        10'b1011111010: data <= 13'h0000; 
        10'b1011111011: data <= 13'h1ffe; 
        10'b1011111100: data <= 13'h1fff; 
        10'b1011111101: data <= 13'h1ff8; 
        10'b1011111110: data <= 13'h1ffa; 
        10'b1011111111: data <= 13'h1ffe; 
        10'b1100000000: data <= 13'h1ffa; 
        10'b1100000001: data <= 13'h1fff; 
        10'b1100000010: data <= 13'h1ffb; 
        10'b1100000011: data <= 13'h1ffd; 
        10'b1100000100: data <= 13'h1ffb; 
        10'b1100000101: data <= 13'h0000; 
        10'b1100000110: data <= 13'h1ff9; 
        10'b1100000111: data <= 13'h1ffa; 
        10'b1100001000: data <= 13'h1fff; 
        10'b1100001001: data <= 13'h1ffd; 
        10'b1100001010: data <= 13'h1ffa; 
        10'b1100001011: data <= 13'h1ffe; 
        10'b1100001100: data <= 13'h1ff9; 
        10'b1100001101: data <= 13'h1ff8; 
        10'b1100001110: data <= 13'h0000; 
        10'b1100001111: data <= 13'h1ffc; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 8) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 14'h3ffb; 
        10'b0000000001: data <= 14'h3ff4; 
        10'b0000000010: data <= 14'h3fff; 
        10'b0000000011: data <= 14'h0001; 
        10'b0000000100: data <= 14'h0001; 
        10'b0000000101: data <= 14'h3fff; 
        10'b0000000110: data <= 14'h3ffb; 
        10'b0000000111: data <= 14'h0001; 
        10'b0000001000: data <= 14'h3ff6; 
        10'b0000001001: data <= 14'h0001; 
        10'b0000001010: data <= 14'h0001; 
        10'b0000001011: data <= 14'h3ff7; 
        10'b0000001100: data <= 14'h3ff7; 
        10'b0000001101: data <= 14'h3ff7; 
        10'b0000001110: data <= 14'h3ff8; 
        10'b0000001111: data <= 14'h3ff9; 
        10'b0000010000: data <= 14'h0000; 
        10'b0000010001: data <= 14'h0001; 
        10'b0000010010: data <= 14'h3ff4; 
        10'b0000010011: data <= 14'h0001; 
        10'b0000010100: data <= 14'h3ffc; 
        10'b0000010101: data <= 14'h3ffd; 
        10'b0000010110: data <= 14'h3ff0; 
        10'b0000010111: data <= 14'h3fff; 
        10'b0000011000: data <= 14'h3fff; 
        10'b0000011001: data <= 14'h3ff1; 
        10'b0000011010: data <= 14'h3ff8; 
        10'b0000011011: data <= 14'h0000; 
        10'b0000011100: data <= 14'h3ff3; 
        10'b0000011101: data <= 14'h3ff8; 
        10'b0000011110: data <= 14'h3ff3; 
        10'b0000011111: data <= 14'h3ffc; 
        10'b0000100000: data <= 14'h3ff2; 
        10'b0000100001: data <= 14'h3ff9; 
        10'b0000100010: data <= 14'h0002; 
        10'b0000100011: data <= 14'h0001; 
        10'b0000100100: data <= 14'h3ff1; 
        10'b0000100101: data <= 14'h3ff0; 
        10'b0000100110: data <= 14'h3ff1; 
        10'b0000100111: data <= 14'h3ffb; 
        10'b0000101000: data <= 14'h3ffd; 
        10'b0000101001: data <= 14'h3ff9; 
        10'b0000101010: data <= 14'h3ff7; 
        10'b0000101011: data <= 14'h3ff4; 
        10'b0000101100: data <= 14'h0002; 
        10'b0000101101: data <= 14'h3ff4; 
        10'b0000101110: data <= 14'h3ffd; 
        10'b0000101111: data <= 14'h3ff7; 
        10'b0000110000: data <= 14'h3ff7; 
        10'b0000110001: data <= 14'h3ff1; 
        10'b0000110010: data <= 14'h3ffa; 
        10'b0000110011: data <= 14'h3fff; 
        10'b0000110100: data <= 14'h3ff2; 
        10'b0000110101: data <= 14'h3fff; 
        10'b0000110110: data <= 14'h3ffb; 
        10'b0000110111: data <= 14'h3ff3; 
        10'b0000111000: data <= 14'h3ff5; 
        10'b0000111001: data <= 14'h3ffa; 
        10'b0000111010: data <= 14'h3ff9; 
        10'b0000111011: data <= 14'h3ff4; 
        10'b0000111100: data <= 14'h3ffc; 
        10'b0000111101: data <= 14'h3ffd; 
        10'b0000111110: data <= 14'h3ff5; 
        10'b0000111111: data <= 14'h3ffd; 
        10'b0001000000: data <= 14'h3fff; 
        10'b0001000001: data <= 14'h3ff9; 
        10'b0001000010: data <= 14'h3ff2; 
        10'b0001000011: data <= 14'h3ff3; 
        10'b0001000100: data <= 14'h3ff1; 
        10'b0001000101: data <= 14'h3ff3; 
        10'b0001000110: data <= 14'h3ff8; 
        10'b0001000111: data <= 14'h3ff6; 
        10'b0001001000: data <= 14'h3ff5; 
        10'b0001001001: data <= 14'h3ff5; 
        10'b0001001010: data <= 14'h3ffd; 
        10'b0001001011: data <= 14'h0000; 
        10'b0001001100: data <= 14'h3ff8; 
        10'b0001001101: data <= 14'h3ff3; 
        10'b0001001110: data <= 14'h0001; 
        10'b0001001111: data <= 14'h3fff; 
        10'b0001010000: data <= 14'h0000; 
        10'b0001010001: data <= 14'h3ff6; 
        10'b0001010010: data <= 14'h3ff0; 
        10'b0001010011: data <= 14'h3ff9; 
        10'b0001010100: data <= 14'h0002; 
        10'b0001010101: data <= 14'h3ffd; 
        10'b0001010110: data <= 14'h3ff9; 
        10'b0001010111: data <= 14'h3ffe; 
        10'b0001011000: data <= 14'h3ffd; 
        10'b0001011001: data <= 14'h0000; 
        10'b0001011010: data <= 14'h3ffb; 
        10'b0001011011: data <= 14'h3fff; 
        10'b0001011100: data <= 14'h3ffe; 
        10'b0001011101: data <= 14'h3ffa; 
        10'b0001011110: data <= 14'h0006; 
        10'b0001011111: data <= 14'h0013; 
        10'b0001100000: data <= 14'h0027; 
        10'b0001100001: data <= 14'h0020; 
        10'b0001100010: data <= 14'h0021; 
        10'b0001100011: data <= 14'h0025; 
        10'b0001100100: data <= 14'h0019; 
        10'b0001100101: data <= 14'h001d; 
        10'b0001100110: data <= 14'h0016; 
        10'b0001100111: data <= 14'h0002; 
        10'b0001101000: data <= 14'h3ffe; 
        10'b0001101001: data <= 14'h3fe5; 
        10'b0001101010: data <= 14'h3ff0; 
        10'b0001101011: data <= 14'h3fff; 
        10'b0001101100: data <= 14'h0001; 
        10'b0001101101: data <= 14'h3ff4; 
        10'b0001101110: data <= 14'h3ffb; 
        10'b0001101111: data <= 14'h3ff5; 
        10'b0001110000: data <= 14'h3ffa; 
        10'b0001110001: data <= 14'h3fff; 
        10'b0001110010: data <= 14'h3ffc; 
        10'b0001110011: data <= 14'h0000; 
        10'b0001110100: data <= 14'h0006; 
        10'b0001110101: data <= 14'h0000; 
        10'b0001110110: data <= 14'h0017; 
        10'b0001110111: data <= 14'h0013; 
        10'b0001111000: data <= 14'h0035; 
        10'b0001111001: data <= 14'h002d; 
        10'b0001111010: data <= 14'h0038; 
        10'b0001111011: data <= 14'h0044; 
        10'b0001111100: data <= 14'h004f; 
        10'b0001111101: data <= 14'h0054; 
        10'b0001111110: data <= 14'h004c; 
        10'b0001111111: data <= 14'h0038; 
        10'b0010000000: data <= 14'h001f; 
        10'b0010000001: data <= 14'h0019; 
        10'b0010000010: data <= 14'h0029; 
        10'b0010000011: data <= 14'h0005; 
        10'b0010000100: data <= 14'h3fe4; 
        10'b0010000101: data <= 14'h3fd4; 
        10'b0010000110: data <= 14'h3fdb; 
        10'b0010000111: data <= 14'h3fdb; 
        10'b0010001000: data <= 14'h3ffc; 
        10'b0010001001: data <= 14'h3ff9; 
        10'b0010001010: data <= 14'h3ff6; 
        10'b0010001011: data <= 14'h3ffe; 
        10'b0010001100: data <= 14'h3ff2; 
        10'b0010001101: data <= 14'h3ff0; 
        10'b0010001110: data <= 14'h3ff4; 
        10'b0010001111: data <= 14'h3ff4; 
        10'b0010010000: data <= 14'h0003; 
        10'b0010010001: data <= 14'h0018; 
        10'b0010010010: data <= 14'h002c; 
        10'b0010010011: data <= 14'h0023; 
        10'b0010010100: data <= 14'h0028; 
        10'b0010010101: data <= 14'h0023; 
        10'b0010010110: data <= 14'h0020; 
        10'b0010010111: data <= 14'h002a; 
        10'b0010011000: data <= 14'h002a; 
        10'b0010011001: data <= 14'h0033; 
        10'b0010011010: data <= 14'h0009; 
        10'b0010011011: data <= 14'h0022; 
        10'b0010011100: data <= 14'h0027; 
        10'b0010011101: data <= 14'h3ffd; 
        10'b0010011110: data <= 14'h3ffe; 
        10'b0010011111: data <= 14'h3fee; 
        10'b0010100000: data <= 14'h3fe7; 
        10'b0010100001: data <= 14'h3fcc; 
        10'b0010100010: data <= 14'h3fbd; 
        10'b0010100011: data <= 14'h3fc8; 
        10'b0010100100: data <= 14'h3ff0; 
        10'b0010100101: data <= 14'h0000; 
        10'b0010100110: data <= 14'h3ff5; 
        10'b0010100111: data <= 14'h3ff9; 
        10'b0010101000: data <= 14'h3ff4; 
        10'b0010101001: data <= 14'h3ff6; 
        10'b0010101010: data <= 14'h3ff5; 
        10'b0010101011: data <= 14'h0005; 
        10'b0010101100: data <= 14'h001e; 
        10'b0010101101: data <= 14'h0037; 
        10'b0010101110: data <= 14'h002a; 
        10'b0010101111: data <= 14'h0020; 
        10'b0010110000: data <= 14'h0031; 
        10'b0010110001: data <= 14'h0028; 
        10'b0010110010: data <= 14'h0023; 
        10'b0010110011: data <= 14'h0022; 
        10'b0010110100: data <= 14'h002d; 
        10'b0010110101: data <= 14'h0041; 
        10'b0010110110: data <= 14'h002d; 
        10'b0010110111: data <= 14'h0010; 
        10'b0010111000: data <= 14'h002b; 
        10'b0010111001: data <= 14'h0027; 
        10'b0010111010: data <= 14'h0026; 
        10'b0010111011: data <= 14'h3fef; 
        10'b0010111100: data <= 14'h0010; 
        10'b0010111101: data <= 14'h3ff0; 
        10'b0010111110: data <= 14'h3fc7; 
        10'b0010111111: data <= 14'h3fc7; 
        10'b0011000000: data <= 14'h3fdd; 
        10'b0011000001: data <= 14'h3ff9; 
        10'b0011000010: data <= 14'h3ffe; 
        10'b0011000011: data <= 14'h3ffb; 
        10'b0011000100: data <= 14'h0001; 
        10'b0011000101: data <= 14'h3ffe; 
        10'b0011000110: data <= 14'h0003; 
        10'b0011000111: data <= 14'h0019; 
        10'b0011001000: data <= 14'h0041; 
        10'b0011001001: data <= 14'h0041; 
        10'b0011001010: data <= 14'h002e; 
        10'b0011001011: data <= 14'h000d; 
        10'b0011001100: data <= 14'h000e; 
        10'b0011001101: data <= 14'h001d; 
        10'b0011001110: data <= 14'h0009; 
        10'b0011001111: data <= 14'h000d; 
        10'b0011010000: data <= 14'h0026; 
        10'b0011010001: data <= 14'h0024; 
        10'b0011010010: data <= 14'h003c; 
        10'b0011010011: data <= 14'h0023; 
        10'b0011010100: data <= 14'h000b; 
        10'b0011010101: data <= 14'h001e; 
        10'b0011010110: data <= 14'h0019; 
        10'b0011010111: data <= 14'h001b; 
        10'b0011011000: data <= 14'h001b; 
        10'b0011011001: data <= 14'h0004; 
        10'b0011011010: data <= 14'h3fe4; 
        10'b0011011011: data <= 14'h3fc0; 
        10'b0011011100: data <= 14'h3fd2; 
        10'b0011011101: data <= 14'h3ff4; 
        10'b0011011110: data <= 14'h3ff0; 
        10'b0011011111: data <= 14'h3ff8; 
        10'b0011100000: data <= 14'h3ffa; 
        10'b0011100001: data <= 14'h3ff7; 
        10'b0011100010: data <= 14'h0003; 
        10'b0011100011: data <= 14'h0017; 
        10'b0011100100: data <= 14'h0036; 
        10'b0011100101: data <= 14'h0033; 
        10'b0011100110: data <= 14'h0026; 
        10'b0011100111: data <= 14'h0010; 
        10'b0011101000: data <= 14'h001a; 
        10'b0011101001: data <= 14'h000c; 
        10'b0011101010: data <= 14'h0021; 
        10'b0011101011: data <= 14'h000a; 
        10'b0011101100: data <= 14'h0009; 
        10'b0011101101: data <= 14'h0010; 
        10'b0011101110: data <= 14'h0041; 
        10'b0011101111: data <= 14'h0036; 
        10'b0011110000: data <= 14'h000c; 
        10'b0011110001: data <= 14'h001e; 
        10'b0011110010: data <= 14'h002b; 
        10'b0011110011: data <= 14'h001c; 
        10'b0011110100: data <= 14'h0029; 
        10'b0011110101: data <= 14'h0015; 
        10'b0011110110: data <= 14'h3ff5; 
        10'b0011110111: data <= 14'h3fc5; 
        10'b0011111000: data <= 14'h3fd4; 
        10'b0011111001: data <= 14'h3ff0; 
        10'b0011111010: data <= 14'h3ff2; 
        10'b0011111011: data <= 14'h3ff6; 
        10'b0011111100: data <= 14'h3ff8; 
        10'b0011111101: data <= 14'h3ff1; 
        10'b0011111110: data <= 14'h3ffb; 
        10'b0011111111: data <= 14'h000a; 
        10'b0100000000: data <= 14'h001c; 
        10'b0100000001: data <= 14'h0025; 
        10'b0100000010: data <= 14'h001e; 
        10'b0100000011: data <= 14'h0007; 
        10'b0100000100: data <= 14'h3ffc; 
        10'b0100000101: data <= 14'h3fe4; 
        10'b0100000110: data <= 14'h3fca; 
        10'b0100000111: data <= 14'h3f9d; 
        10'b0100001000: data <= 14'h3faf; 
        10'b0100001001: data <= 14'h3ff5; 
        10'b0100001010: data <= 14'h004d; 
        10'b0100001011: data <= 14'h0077; 
        10'b0100001100: data <= 14'h0045; 
        10'b0100001101: data <= 14'h0028; 
        10'b0100001110: data <= 14'h002c; 
        10'b0100001111: data <= 14'h0028; 
        10'b0100010000: data <= 14'h003c; 
        10'b0100010001: data <= 14'h0027; 
        10'b0100010010: data <= 14'h3ff4; 
        10'b0100010011: data <= 14'h3fc5; 
        10'b0100010100: data <= 14'h3fe2; 
        10'b0100010101: data <= 14'h3fef; 
        10'b0100010110: data <= 14'h3ff3; 
        10'b0100010111: data <= 14'h3ff5; 
        10'b0100011000: data <= 14'h3ffe; 
        10'b0100011001: data <= 14'h3ffd; 
        10'b0100011010: data <= 14'h0001; 
        10'b0100011011: data <= 14'h000f; 
        10'b0100011100: data <= 14'h000d; 
        10'b0100011101: data <= 14'h0006; 
        10'b0100011110: data <= 14'h3fef; 
        10'b0100011111: data <= 14'h3fd4; 
        10'b0100100000: data <= 14'h3fb0; 
        10'b0100100001: data <= 14'h3f8d; 
        10'b0100100010: data <= 14'h3f74; 
        10'b0100100011: data <= 14'h3f70; 
        10'b0100100100: data <= 14'h3f96; 
        10'b0100100101: data <= 14'h3fe5; 
        10'b0100100110: data <= 14'h003f; 
        10'b0100100111: data <= 14'h0049; 
        10'b0100101000: data <= 14'h003e; 
        10'b0100101001: data <= 14'h003a; 
        10'b0100101010: data <= 14'h0024; 
        10'b0100101011: data <= 14'h003e; 
        10'b0100101100: data <= 14'h003a; 
        10'b0100101101: data <= 14'h0017; 
        10'b0100101110: data <= 14'h3feb; 
        10'b0100101111: data <= 14'h3fda; 
        10'b0100110000: data <= 14'h3ff2; 
        10'b0100110001: data <= 14'h3ff0; 
        10'b0100110010: data <= 14'h3ff9; 
        10'b0100110011: data <= 14'h3ffe; 
        10'b0100110100: data <= 14'h0002; 
        10'b0100110101: data <= 14'h3ffe; 
        10'b0100110110: data <= 14'h3ff3; 
        10'b0100110111: data <= 14'h000f; 
        10'b0100111000: data <= 14'h3ff7; 
        10'b0100111001: data <= 14'h3fd3; 
        10'b0100111010: data <= 14'h3fbd; 
        10'b0100111011: data <= 14'h3f9d; 
        10'b0100111100: data <= 14'h3f84; 
        10'b0100111101: data <= 14'h3f95; 
        10'b0100111110: data <= 14'h3faf; 
        10'b0100111111: data <= 14'h3fda; 
        10'b0101000000: data <= 14'h3feb; 
        10'b0101000001: data <= 14'h001b; 
        10'b0101000010: data <= 14'h002a; 
        10'b0101000011: data <= 14'h002a; 
        10'b0101000100: data <= 14'h0013; 
        10'b0101000101: data <= 14'h002c; 
        10'b0101000110: data <= 14'h0036; 
        10'b0101000111: data <= 14'h0035; 
        10'b0101001000: data <= 14'h002e; 
        10'b0101001001: data <= 14'h0000; 
        10'b0101001010: data <= 14'h3fec; 
        10'b0101001011: data <= 14'h3fef; 
        10'b0101001100: data <= 14'h3ff1; 
        10'b0101001101: data <= 14'h3ff7; 
        10'b0101001110: data <= 14'h3ff4; 
        10'b0101001111: data <= 14'h3ff2; 
        10'b0101010000: data <= 14'h0001; 
        10'b0101010001: data <= 14'h3ff6; 
        10'b0101010010: data <= 14'h3ffd; 
        10'b0101010011: data <= 14'h3fff; 
        10'b0101010100: data <= 14'h3ff0; 
        10'b0101010101: data <= 14'h3fd3; 
        10'b0101010110: data <= 14'h3fb1; 
        10'b0101010111: data <= 14'h3f9d; 
        10'b0101011000: data <= 14'h3fa7; 
        10'b0101011001: data <= 14'h3fd0; 
        10'b0101011010: data <= 14'h0001; 
        10'b0101011011: data <= 14'h0008; 
        10'b0101011100: data <= 14'h000d; 
        10'b0101011101: data <= 14'h001d; 
        10'b0101011110: data <= 14'h0047; 
        10'b0101011111: data <= 14'h0025; 
        10'b0101100000: data <= 14'h0019; 
        10'b0101100001: data <= 14'h0023; 
        10'b0101100010: data <= 14'h001c; 
        10'b0101100011: data <= 14'h3ffe; 
        10'b0101100100: data <= 14'h3fdb; 
        10'b0101100101: data <= 14'h3fce; 
        10'b0101100110: data <= 14'h3fcb; 
        10'b0101100111: data <= 14'h3fdf; 
        10'b0101101000: data <= 14'h3ffa; 
        10'b0101101001: data <= 14'h3ff6; 
        10'b0101101010: data <= 14'h3ffb; 
        10'b0101101011: data <= 14'h3ffc; 
        10'b0101101100: data <= 14'h3ff9; 
        10'b0101101101: data <= 14'h3ff5; 
        10'b0101101110: data <= 14'h3ff9; 
        10'b0101101111: data <= 14'h3ffc; 
        10'b0101110000: data <= 14'h3feb; 
        10'b0101110001: data <= 14'h3fe1; 
        10'b0101110010: data <= 14'h3fc0; 
        10'b0101110011: data <= 14'h3fb6; 
        10'b0101110100: data <= 14'h3fce; 
        10'b0101110101: data <= 14'h3ff6; 
        10'b0101110110: data <= 14'h3ff0; 
        10'b0101110111: data <= 14'h3fd5; 
        10'b0101111000: data <= 14'h0003; 
        10'b0101111001: data <= 14'h003d; 
        10'b0101111010: data <= 14'h003d; 
        10'b0101111011: data <= 14'h000b; 
        10'b0101111100: data <= 14'h001c; 
        10'b0101111101: data <= 14'h001e; 
        10'b0101111110: data <= 14'h0010; 
        10'b0101111111: data <= 14'h3feb; 
        10'b0110000000: data <= 14'h3fc8; 
        10'b0110000001: data <= 14'h3fc8; 
        10'b0110000010: data <= 14'h3fd3; 
        10'b0110000011: data <= 14'h3fe1; 
        10'b0110000100: data <= 14'h3fee; 
        10'b0110000101: data <= 14'h0000; 
        10'b0110000110: data <= 14'h3ffd; 
        10'b0110000111: data <= 14'h3ff6; 
        10'b0110001000: data <= 14'h0001; 
        10'b0110001001: data <= 14'h3ff4; 
        10'b0110001010: data <= 14'h3ff8; 
        10'b0110001011: data <= 14'h3ffb; 
        10'b0110001100: data <= 14'h3ffc; 
        10'b0110001101: data <= 14'h3fe6; 
        10'b0110001110: data <= 14'h3fc6; 
        10'b0110001111: data <= 14'h3fcc; 
        10'b0110010000: data <= 14'h3fdc; 
        10'b0110010001: data <= 14'h3ffb; 
        10'b0110010010: data <= 14'h3fdb; 
        10'b0110010011: data <= 14'h3fd8; 
        10'b0110010100: data <= 14'h000b; 
        10'b0110010101: data <= 14'h001d; 
        10'b0110010110: data <= 14'h001f; 
        10'b0110010111: data <= 14'h3ffb; 
        10'b0110011000: data <= 14'h3ff3; 
        10'b0110011001: data <= 14'h3ff6; 
        10'b0110011010: data <= 14'h0004; 
        10'b0110011011: data <= 14'h3fe8; 
        10'b0110011100: data <= 14'h3fdf; 
        10'b0110011101: data <= 14'h3ff0; 
        10'b0110011110: data <= 14'h3fe9; 
        10'b0110011111: data <= 14'h3ff1; 
        10'b0110100000: data <= 14'h3fec; 
        10'b0110100001: data <= 14'h3fee; 
        10'b0110100010: data <= 14'h0000; 
        10'b0110100011: data <= 14'h0001; 
        10'b0110100100: data <= 14'h0001; 
        10'b0110100101: data <= 14'h3ff4; 
        10'b0110100110: data <= 14'h0002; 
        10'b0110100111: data <= 14'h0004; 
        10'b0110101000: data <= 14'h3ffb; 
        10'b0110101001: data <= 14'h3fe3; 
        10'b0110101010: data <= 14'h3fca; 
        10'b0110101011: data <= 14'h3fc6; 
        10'b0110101100: data <= 14'h3fd5; 
        10'b0110101101: data <= 14'h3fe7; 
        10'b0110101110: data <= 14'h3fe4; 
        10'b0110101111: data <= 14'h3ff7; 
        10'b0110110000: data <= 14'h000c; 
        10'b0110110001: data <= 14'h0030; 
        10'b0110110010: data <= 14'h001b; 
        10'b0110110011: data <= 14'h3ffd; 
        10'b0110110100: data <= 14'h3fd8; 
        10'b0110110101: data <= 14'h3ff4; 
        10'b0110110110: data <= 14'h3ffc; 
        10'b0110110111: data <= 14'h000b; 
        10'b0110111000: data <= 14'h0019; 
        10'b0110111001: data <= 14'h0018; 
        10'b0110111010: data <= 14'h0008; 
        10'b0110111011: data <= 14'h0003; 
        10'b0110111100: data <= 14'h3ff1; 
        10'b0110111101: data <= 14'h3ffd; 
        10'b0110111110: data <= 14'h3ffb; 
        10'b0110111111: data <= 14'h3ff4; 
        10'b0111000000: data <= 14'h3ffb; 
        10'b0111000001: data <= 14'h3ffd; 
        10'b0111000010: data <= 14'h000b; 
        10'b0111000011: data <= 14'h0002; 
        10'b0111000100: data <= 14'h0008; 
        10'b0111000101: data <= 14'h3ff3; 
        10'b0111000110: data <= 14'h3fea; 
        10'b0111000111: data <= 14'h3fda; 
        10'b0111001000: data <= 14'h3fad; 
        10'b0111001001: data <= 14'h3fa9; 
        10'b0111001010: data <= 14'h3fb3; 
        10'b0111001011: data <= 14'h3fec; 
        10'b0111001100: data <= 14'h0017; 
        10'b0111001101: data <= 14'h003c; 
        10'b0111001110: data <= 14'h3ffa; 
        10'b0111001111: data <= 14'h3fd4; 
        10'b0111010000: data <= 14'h3fd2; 
        10'b0111010001: data <= 14'h3ff1; 
        10'b0111010010: data <= 14'h0013; 
        10'b0111010011: data <= 14'h0033; 
        10'b0111010100: data <= 14'h0024; 
        10'b0111010101: data <= 14'h002d; 
        10'b0111010110: data <= 14'h002c; 
        10'b0111010111: data <= 14'h0013; 
        10'b0111011000: data <= 14'h3ffa; 
        10'b0111011001: data <= 14'h3ffc; 
        10'b0111011010: data <= 14'h3fff; 
        10'b0111011011: data <= 14'h3fff; 
        10'b0111011100: data <= 14'h3ffe; 
        10'b0111011101: data <= 14'h0002; 
        10'b0111011110: data <= 14'h0000; 
        10'b0111011111: data <= 14'h001c; 
        10'b0111100000: data <= 14'h000f; 
        10'b0111100001: data <= 14'h0005; 
        10'b0111100010: data <= 14'h3ff1; 
        10'b0111100011: data <= 14'h3fce; 
        10'b0111100100: data <= 14'h3fa7; 
        10'b0111100101: data <= 14'h3f72; 
        10'b0111100110: data <= 14'h3f50; 
        10'b0111100111: data <= 14'h3f5f; 
        10'b0111101000: data <= 14'h3f86; 
        10'b0111101001: data <= 14'h3fba; 
        10'b0111101010: data <= 14'h3fbf; 
        10'b0111101011: data <= 14'h3fc6; 
        10'b0111101100: data <= 14'h3ffe; 
        10'b0111101101: data <= 14'h0012; 
        10'b0111101110: data <= 14'h0021; 
        10'b0111101111: data <= 14'h0034; 
        10'b0111110000: data <= 14'h000b; 
        10'b0111110001: data <= 14'h003e; 
        10'b0111110010: data <= 14'h003e; 
        10'b0111110011: data <= 14'h0013; 
        10'b0111110100: data <= 14'h3ff7; 
        10'b0111110101: data <= 14'h3ff3; 
        10'b0111110110: data <= 14'h3ff4; 
        10'b0111110111: data <= 14'h3ff5; 
        10'b0111111000: data <= 14'h3ff9; 
        10'b0111111001: data <= 14'h3ffa; 
        10'b0111111010: data <= 14'h0005; 
        10'b0111111011: data <= 14'h0029; 
        10'b0111111100: data <= 14'h001e; 
        10'b0111111101: data <= 14'h0012; 
        10'b0111111110: data <= 14'h0009; 
        10'b0111111111: data <= 14'h3ff5; 
        10'b1000000000: data <= 14'h3fe0; 
        10'b1000000001: data <= 14'h3f98; 
        10'b1000000010: data <= 14'h3f67; 
        10'b1000000011: data <= 14'h3f6f; 
        10'b1000000100: data <= 14'h3f51; 
        10'b1000000101: data <= 14'h3f71; 
        10'b1000000110: data <= 14'h3fa6; 
        10'b1000000111: data <= 14'h3feb; 
        10'b1000001000: data <= 14'h0024; 
        10'b1000001001: data <= 14'h0031; 
        10'b1000001010: data <= 14'h0035; 
        10'b1000001011: data <= 14'h0034; 
        10'b1000001100: data <= 14'h0025; 
        10'b1000001101: data <= 14'h0049; 
        10'b1000001110: data <= 14'h0044; 
        10'b1000001111: data <= 14'h001a; 
        10'b1000010000: data <= 14'h3fe8; 
        10'b1000010001: data <= 14'h3ff0; 
        10'b1000010010: data <= 14'h3ff4; 
        10'b1000010011: data <= 14'h3ffe; 
        10'b1000010100: data <= 14'h3ffe; 
        10'b1000010101: data <= 14'h3ff4; 
        10'b1000010110: data <= 14'h3ff8; 
        10'b1000010111: data <= 14'h0034; 
        10'b1000011000: data <= 14'h0035; 
        10'b1000011001: data <= 14'h003e; 
        10'b1000011010: data <= 14'h0035; 
        10'b1000011011: data <= 14'h0014; 
        10'b1000011100: data <= 14'h0006; 
        10'b1000011101: data <= 14'h3fea; 
        10'b1000011110: data <= 14'h3ff0; 
        10'b1000011111: data <= 14'h3fcf; 
        10'b1000100000: data <= 14'h3fb8; 
        10'b1000100001: data <= 14'h3fb3; 
        10'b1000100010: data <= 14'h3fcc; 
        10'b1000100011: data <= 14'h0012; 
        10'b1000100100: data <= 14'h0031; 
        10'b1000100101: data <= 14'h003e; 
        10'b1000100110: data <= 14'h0045; 
        10'b1000100111: data <= 14'h003e; 
        10'b1000101000: data <= 14'h0037; 
        10'b1000101001: data <= 14'h0040; 
        10'b1000101010: data <= 14'h0018; 
        10'b1000101011: data <= 14'h0003; 
        10'b1000101100: data <= 14'h3fec; 
        10'b1000101101: data <= 14'h3ffc; 
        10'b1000101110: data <= 14'h3ffe; 
        10'b1000101111: data <= 14'h3ffc; 
        10'b1000110000: data <= 14'h3ffd; 
        10'b1000110001: data <= 14'h3ff0; 
        10'b1000110010: data <= 14'h0009; 
        10'b1000110011: data <= 14'h0038; 
        10'b1000110100: data <= 14'h0044; 
        10'b1000110101: data <= 14'h004a; 
        10'b1000110110: data <= 14'h004e; 
        10'b1000110111: data <= 14'h0027; 
        10'b1000111000: data <= 14'h002e; 
        10'b1000111001: data <= 14'h0035; 
        10'b1000111010: data <= 14'h0013; 
        10'b1000111011: data <= 14'h3ffb; 
        10'b1000111100: data <= 14'h3fee; 
        10'b1000111101: data <= 14'h3fe5; 
        10'b1000111110: data <= 14'h0008; 
        10'b1000111111: data <= 14'h000f; 
        10'b1001000000: data <= 14'h001c; 
        10'b1001000001: data <= 14'h0032; 
        10'b1001000010: data <= 14'h0034; 
        10'b1001000011: data <= 14'h0023; 
        10'b1001000100: data <= 14'h003d; 
        10'b1001000101: data <= 14'h0023; 
        10'b1001000110: data <= 14'h3ff9; 
        10'b1001000111: data <= 14'h3ff2; 
        10'b1001001000: data <= 14'h3ff0; 
        10'b1001001001: data <= 14'h3ffb; 
        10'b1001001010: data <= 14'h3ffb; 
        10'b1001001011: data <= 14'h3ffa; 
        10'b1001001100: data <= 14'h3ff5; 
        10'b1001001101: data <= 14'h3fff; 
        10'b1001001110: data <= 14'h3ffc; 
        10'b1001001111: data <= 14'h001c; 
        10'b1001010000: data <= 14'h0042; 
        10'b1001010001: data <= 14'h0042; 
        10'b1001010010: data <= 14'h0039; 
        10'b1001010011: data <= 14'h0020; 
        10'b1001010100: data <= 14'h0023; 
        10'b1001010101: data <= 14'h000b; 
        10'b1001010110: data <= 14'h3ffb; 
        10'b1001010111: data <= 14'h3ff0; 
        10'b1001011000: data <= 14'h0005; 
        10'b1001011001: data <= 14'h3ffd; 
        10'b1001011010: data <= 14'h3ffc; 
        10'b1001011011: data <= 14'h3ff8; 
        10'b1001011100: data <= 14'h0010; 
        10'b1001011101: data <= 14'h0006; 
        10'b1001011110: data <= 14'h0020; 
        10'b1001011111: data <= 14'h0033; 
        10'b1001100000: data <= 14'h001e; 
        10'b1001100001: data <= 14'h000b; 
        10'b1001100010: data <= 14'h3ff5; 
        10'b1001100011: data <= 14'h3fe2; 
        10'b1001100100: data <= 14'h3ff6; 
        10'b1001100101: data <= 14'h3ff4; 
        10'b1001100110: data <= 14'h3ff0; 
        10'b1001100111: data <= 14'h3ff1; 
        10'b1001101000: data <= 14'h3ff9; 
        10'b1001101001: data <= 14'h3ffb; 
        10'b1001101010: data <= 14'h3ffd; 
        10'b1001101011: data <= 14'h0011; 
        10'b1001101100: data <= 14'h0021; 
        10'b1001101101: data <= 14'h002d; 
        10'b1001101110: data <= 14'h0028; 
        10'b1001101111: data <= 14'h0017; 
        10'b1001110000: data <= 14'h0002; 
        10'b1001110001: data <= 14'h0011; 
        10'b1001110010: data <= 14'h0014; 
        10'b1001110011: data <= 14'h0018; 
        10'b1001110100: data <= 14'h0007; 
        10'b1001110101: data <= 14'h3ff7; 
        10'b1001110110: data <= 14'h3ff7; 
        10'b1001110111: data <= 14'h3ff3; 
        10'b1001111000: data <= 14'h000a; 
        10'b1001111001: data <= 14'h0008; 
        10'b1001111010: data <= 14'h0008; 
        10'b1001111011: data <= 14'h0023; 
        10'b1001111100: data <= 14'h0011; 
        10'b1001111101: data <= 14'h3ffa; 
        10'b1001111110: data <= 14'h3ff8; 
        10'b1001111111: data <= 14'h3ff6; 
        10'b1010000000: data <= 14'h3fe9; 
        10'b1010000001: data <= 14'h3fef; 
        10'b1010000010: data <= 14'h3ffd; 
        10'b1010000011: data <= 14'h0000; 
        10'b1010000100: data <= 14'h3ffb; 
        10'b1010000101: data <= 14'h3ff3; 
        10'b1010000110: data <= 14'h3ff5; 
        10'b1010000111: data <= 14'h000b; 
        10'b1010001000: data <= 14'h0024; 
        10'b1010001001: data <= 14'h0037; 
        10'b1010001010: data <= 14'h0029; 
        10'b1010001011: data <= 14'h002b; 
        10'b1010001100: data <= 14'h000a; 
        10'b1010001101: data <= 14'h001c; 
        10'b1010001110: data <= 14'h0011; 
        10'b1010001111: data <= 14'h0000; 
        10'b1010010000: data <= 14'h3ff2; 
        10'b1010010001: data <= 14'h0002; 
        10'b1010010010: data <= 14'h0006; 
        10'b1010010011: data <= 14'h000e; 
        10'b1010010100: data <= 14'h000a; 
        10'b1010010101: data <= 14'h0015; 
        10'b1010010110: data <= 14'h0022; 
        10'b1010010111: data <= 14'h3ffa; 
        10'b1010011000: data <= 14'h3fe9; 
        10'b1010011001: data <= 14'h3fea; 
        10'b1010011010: data <= 14'h3ff4; 
        10'b1010011011: data <= 14'h3ff1; 
        10'b1010011100: data <= 14'h3fff; 
        10'b1010011101: data <= 14'h3ffc; 
        10'b1010011110: data <= 14'h3ff2; 
        10'b1010011111: data <= 14'h3ff3; 
        10'b1010100000: data <= 14'h3ff6; 
        10'b1010100001: data <= 14'h0002; 
        10'b1010100010: data <= 14'h0002; 
        10'b1010100011: data <= 14'h0000; 
        10'b1010100100: data <= 14'h0017; 
        10'b1010100101: data <= 14'h0025; 
        10'b1010100110: data <= 14'h002c; 
        10'b1010100111: data <= 14'h0034; 
        10'b1010101000: data <= 14'h0035; 
        10'b1010101001: data <= 14'h002b; 
        10'b1010101010: data <= 14'h003f; 
        10'b1010101011: data <= 14'h0043; 
        10'b1010101100: data <= 14'h0044; 
        10'b1010101101: data <= 14'h0036; 
        10'b1010101110: data <= 14'h002f; 
        10'b1010101111: data <= 14'h0023; 
        10'b1010110000: data <= 14'h0022; 
        10'b1010110001: data <= 14'h3ffd; 
        10'b1010110010: data <= 14'h3fe5; 
        10'b1010110011: data <= 14'h3fda; 
        10'b1010110100: data <= 14'h3fde; 
        10'b1010110101: data <= 14'h3feb; 
        10'b1010110110: data <= 14'h3fed; 
        10'b1010110111: data <= 14'h3ffa; 
        10'b1010111000: data <= 14'h3ff6; 
        10'b1010111001: data <= 14'h0000; 
        10'b1010111010: data <= 14'h3ff6; 
        10'b1010111011: data <= 14'h0002; 
        10'b1010111100: data <= 14'h3ffe; 
        10'b1010111101: data <= 14'h3ff0; 
        10'b1010111110: data <= 14'h0001; 
        10'b1010111111: data <= 14'h0003; 
        10'b1011000000: data <= 14'h3ffc; 
        10'b1011000001: data <= 14'h000f; 
        10'b1011000010: data <= 14'h0016; 
        10'b1011000011: data <= 14'h000c; 
        10'b1011000100: data <= 14'h001e; 
        10'b1011000101: data <= 14'h001e; 
        10'b1011000110: data <= 14'h0038; 
        10'b1011000111: data <= 14'h0040; 
        10'b1011001000: data <= 14'h0045; 
        10'b1011001001: data <= 14'h0036; 
        10'b1011001010: data <= 14'h0026; 
        10'b1011001011: data <= 14'h000f; 
        10'b1011001100: data <= 14'h3ffa; 
        10'b1011001101: data <= 14'h3fe8; 
        10'b1011001110: data <= 14'h3fe8; 
        10'b1011001111: data <= 14'h3fec; 
        10'b1011010000: data <= 14'h3fec; 
        10'b1011010001: data <= 14'h3ff6; 
        10'b1011010010: data <= 14'h3ff6; 
        10'b1011010011: data <= 14'h3fff; 
        10'b1011010100: data <= 14'h3ff4; 
        10'b1011010101: data <= 14'h0002; 
        10'b1011010110: data <= 14'h3ff0; 
        10'b1011010111: data <= 14'h3ffe; 
        10'b1011011000: data <= 14'h3ff5; 
        10'b1011011001: data <= 14'h3ff0; 
        10'b1011011010: data <= 14'h3ff0; 
        10'b1011011011: data <= 14'h3ffc; 
        10'b1011011100: data <= 14'h3ffc; 
        10'b1011011101: data <= 14'h3ff5; 
        10'b1011011110: data <= 14'h3ff3; 
        10'b1011011111: data <= 14'h3ffc; 
        10'b1011100000: data <= 14'h3ffc; 
        10'b1011100001: data <= 14'h3ffb; 
        10'b1011100010: data <= 14'h3ff9; 
        10'b1011100011: data <= 14'h3ffa; 
        10'b1011100100: data <= 14'h3ff7; 
        10'b1011100101: data <= 14'h3ffb; 
        10'b1011100110: data <= 14'h3ff7; 
        10'b1011100111: data <= 14'h3fee; 
        10'b1011101000: data <= 14'h3ff5; 
        10'b1011101001: data <= 14'h3ffb; 
        10'b1011101010: data <= 14'h3ff9; 
        10'b1011101011: data <= 14'h3ffb; 
        10'b1011101100: data <= 14'h3ff1; 
        10'b1011101101: data <= 14'h3ff1; 
        10'b1011101110: data <= 14'h3ffe; 
        10'b1011101111: data <= 14'h3ff7; 
        10'b1011110000: data <= 14'h0000; 
        10'b1011110001: data <= 14'h3ff4; 
        10'b1011110010: data <= 14'h3fff; 
        10'b1011110011: data <= 14'h0002; 
        10'b1011110100: data <= 14'h3ff8; 
        10'b1011110101: data <= 14'h3ff4; 
        10'b1011110110: data <= 14'h3ffb; 
        10'b1011110111: data <= 14'h3ff1; 
        10'b1011111000: data <= 14'h0001; 
        10'b1011111001: data <= 14'h3ffc; 
        10'b1011111010: data <= 14'h3fff; 
        10'b1011111011: data <= 14'h3ffb; 
        10'b1011111100: data <= 14'h3ffd; 
        10'b1011111101: data <= 14'h3ff0; 
        10'b1011111110: data <= 14'h3ff3; 
        10'b1011111111: data <= 14'h3ffd; 
        10'b1100000000: data <= 14'h3ff3; 
        10'b1100000001: data <= 14'h3ffe; 
        10'b1100000010: data <= 14'h3ff6; 
        10'b1100000011: data <= 14'h3ffa; 
        10'b1100000100: data <= 14'h3ff7; 
        10'b1100000101: data <= 14'h0000; 
        10'b1100000110: data <= 14'h3ff1; 
        10'b1100000111: data <= 14'h3ff4; 
        10'b1100001000: data <= 14'h3fff; 
        10'b1100001001: data <= 14'h3ffb; 
        10'b1100001010: data <= 14'h3ff4; 
        10'b1100001011: data <= 14'h3ffc; 
        10'b1100001100: data <= 14'h3ff2; 
        10'b1100001101: data <= 14'h3ff0; 
        10'b1100001110: data <= 14'h3fff; 
        10'b1100001111: data <= 14'h3ff9; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 9) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 15'h7ff6; 
        10'b0000000001: data <= 15'h7fe7; 
        10'b0000000010: data <= 15'h7fff; 
        10'b0000000011: data <= 15'h0001; 
        10'b0000000100: data <= 15'h0003; 
        10'b0000000101: data <= 15'h7ffe; 
        10'b0000000110: data <= 15'h7ff7; 
        10'b0000000111: data <= 15'h0003; 
        10'b0000001000: data <= 15'h7fec; 
        10'b0000001001: data <= 15'h0002; 
        10'b0000001010: data <= 15'h0002; 
        10'b0000001011: data <= 15'h7fef; 
        10'b0000001100: data <= 15'h7fee; 
        10'b0000001101: data <= 15'h7fee; 
        10'b0000001110: data <= 15'h7fef; 
        10'b0000001111: data <= 15'h7ff2; 
        10'b0000010000: data <= 15'h0000; 
        10'b0000010001: data <= 15'h0001; 
        10'b0000010010: data <= 15'h7fe7; 
        10'b0000010011: data <= 15'h0003; 
        10'b0000010100: data <= 15'h7ff8; 
        10'b0000010101: data <= 15'h7ff9; 
        10'b0000010110: data <= 15'h7fdf; 
        10'b0000010111: data <= 15'h7ffe; 
        10'b0000011000: data <= 15'h7fff; 
        10'b0000011001: data <= 15'h7fe1; 
        10'b0000011010: data <= 15'h7ff1; 
        10'b0000011011: data <= 15'h0001; 
        10'b0000011100: data <= 15'h7fe6; 
        10'b0000011101: data <= 15'h7ff0; 
        10'b0000011110: data <= 15'h7fe7; 
        10'b0000011111: data <= 15'h7ff7; 
        10'b0000100000: data <= 15'h7fe3; 
        10'b0000100001: data <= 15'h7ff2; 
        10'b0000100010: data <= 15'h0003; 
        10'b0000100011: data <= 15'h0002; 
        10'b0000100100: data <= 15'h7fe1; 
        10'b0000100101: data <= 15'h7fe0; 
        10'b0000100110: data <= 15'h7fe3; 
        10'b0000100111: data <= 15'h7ff6; 
        10'b0000101000: data <= 15'h7ff9; 
        10'b0000101001: data <= 15'h7ff1; 
        10'b0000101010: data <= 15'h7fef; 
        10'b0000101011: data <= 15'h7fe9; 
        10'b0000101100: data <= 15'h0003; 
        10'b0000101101: data <= 15'h7fe7; 
        10'b0000101110: data <= 15'h7ffa; 
        10'b0000101111: data <= 15'h7fed; 
        10'b0000110000: data <= 15'h7fed; 
        10'b0000110001: data <= 15'h7fe2; 
        10'b0000110010: data <= 15'h7ff3; 
        10'b0000110011: data <= 15'h7ffd; 
        10'b0000110100: data <= 15'h7fe5; 
        10'b0000110101: data <= 15'h7ffe; 
        10'b0000110110: data <= 15'h7ff5; 
        10'b0000110111: data <= 15'h7fe5; 
        10'b0000111000: data <= 15'h7fe9; 
        10'b0000111001: data <= 15'h7ff3; 
        10'b0000111010: data <= 15'h7ff2; 
        10'b0000111011: data <= 15'h7fe7; 
        10'b0000111100: data <= 15'h7ff8; 
        10'b0000111101: data <= 15'h7ffb; 
        10'b0000111110: data <= 15'h7feb; 
        10'b0000111111: data <= 15'h7ffa; 
        10'b0001000000: data <= 15'h7ffd; 
        10'b0001000001: data <= 15'h7ff1; 
        10'b0001000010: data <= 15'h7fe4; 
        10'b0001000011: data <= 15'h7fe5; 
        10'b0001000100: data <= 15'h7fe2; 
        10'b0001000101: data <= 15'h7fe6; 
        10'b0001000110: data <= 15'h7fef; 
        10'b0001000111: data <= 15'h7fed; 
        10'b0001001000: data <= 15'h7feb; 
        10'b0001001001: data <= 15'h7fea; 
        10'b0001001010: data <= 15'h7ffa; 
        10'b0001001011: data <= 15'h7fff; 
        10'b0001001100: data <= 15'h7ff1; 
        10'b0001001101: data <= 15'h7fe7; 
        10'b0001001110: data <= 15'h0003; 
        10'b0001001111: data <= 15'h7ffe; 
        10'b0001010000: data <= 15'h0000; 
        10'b0001010001: data <= 15'h7fec; 
        10'b0001010010: data <= 15'h7fe1; 
        10'b0001010011: data <= 15'h7ff1; 
        10'b0001010100: data <= 15'h0003; 
        10'b0001010101: data <= 15'h7ffa; 
        10'b0001010110: data <= 15'h7ff2; 
        10'b0001010111: data <= 15'h7ffc; 
        10'b0001011000: data <= 15'h7ffa; 
        10'b0001011001: data <= 15'h0000; 
        10'b0001011010: data <= 15'h7ff7; 
        10'b0001011011: data <= 15'h7ffe; 
        10'b0001011100: data <= 15'h7ffc; 
        10'b0001011101: data <= 15'h7ff4; 
        10'b0001011110: data <= 15'h000b; 
        10'b0001011111: data <= 15'h0025; 
        10'b0001100000: data <= 15'h004e; 
        10'b0001100001: data <= 15'h0041; 
        10'b0001100010: data <= 15'h0042; 
        10'b0001100011: data <= 15'h0049; 
        10'b0001100100: data <= 15'h0033; 
        10'b0001100101: data <= 15'h0039; 
        10'b0001100110: data <= 15'h002d; 
        10'b0001100111: data <= 15'h0003; 
        10'b0001101000: data <= 15'h7ffc; 
        10'b0001101001: data <= 15'h7fc9; 
        10'b0001101010: data <= 15'h7fe0; 
        10'b0001101011: data <= 15'h7ffd; 
        10'b0001101100: data <= 15'h0002; 
        10'b0001101101: data <= 15'h7fe8; 
        10'b0001101110: data <= 15'h7ff5; 
        10'b0001101111: data <= 15'h7feb; 
        10'b0001110000: data <= 15'h7ff5; 
        10'b0001110001: data <= 15'h7ffe; 
        10'b0001110010: data <= 15'h7ff7; 
        10'b0001110011: data <= 15'h0001; 
        10'b0001110100: data <= 15'h000c; 
        10'b0001110101: data <= 15'h0000; 
        10'b0001110110: data <= 15'h002e; 
        10'b0001110111: data <= 15'h0027; 
        10'b0001111000: data <= 15'h006a; 
        10'b0001111001: data <= 15'h005b; 
        10'b0001111010: data <= 15'h0071; 
        10'b0001111011: data <= 15'h0088; 
        10'b0001111100: data <= 15'h009d; 
        10'b0001111101: data <= 15'h00a9; 
        10'b0001111110: data <= 15'h0098; 
        10'b0001111111: data <= 15'h006f; 
        10'b0010000000: data <= 15'h003f; 
        10'b0010000001: data <= 15'h0032; 
        10'b0010000010: data <= 15'h0052; 
        10'b0010000011: data <= 15'h000a; 
        10'b0010000100: data <= 15'h7fc8; 
        10'b0010000101: data <= 15'h7fa9; 
        10'b0010000110: data <= 15'h7fb5; 
        10'b0010000111: data <= 15'h7fb7; 
        10'b0010001000: data <= 15'h7ff7; 
        10'b0010001001: data <= 15'h7ff3; 
        10'b0010001010: data <= 15'h7fed; 
        10'b0010001011: data <= 15'h7ffb; 
        10'b0010001100: data <= 15'h7fe4; 
        10'b0010001101: data <= 15'h7fe0; 
        10'b0010001110: data <= 15'h7fe8; 
        10'b0010001111: data <= 15'h7fe8; 
        10'b0010010000: data <= 15'h0006; 
        10'b0010010001: data <= 15'h0030; 
        10'b0010010010: data <= 15'h0057; 
        10'b0010010011: data <= 15'h0046; 
        10'b0010010100: data <= 15'h0050; 
        10'b0010010101: data <= 15'h0046; 
        10'b0010010110: data <= 15'h0040; 
        10'b0010010111: data <= 15'h0053; 
        10'b0010011000: data <= 15'h0054; 
        10'b0010011001: data <= 15'h0065; 
        10'b0010011010: data <= 15'h0011; 
        10'b0010011011: data <= 15'h0043; 
        10'b0010011100: data <= 15'h004e; 
        10'b0010011101: data <= 15'h7ffa; 
        10'b0010011110: data <= 15'h7ffc; 
        10'b0010011111: data <= 15'h7fdd; 
        10'b0010100000: data <= 15'h7fcf; 
        10'b0010100001: data <= 15'h7f98; 
        10'b0010100010: data <= 15'h7f7b; 
        10'b0010100011: data <= 15'h7f8f; 
        10'b0010100100: data <= 15'h7fdf; 
        10'b0010100101: data <= 15'h0000; 
        10'b0010100110: data <= 15'h7fea; 
        10'b0010100111: data <= 15'h7ff2; 
        10'b0010101000: data <= 15'h7fe7; 
        10'b0010101001: data <= 15'h7fed; 
        10'b0010101010: data <= 15'h7fea; 
        10'b0010101011: data <= 15'h000a; 
        10'b0010101100: data <= 15'h003b; 
        10'b0010101101: data <= 15'h006e; 
        10'b0010101110: data <= 15'h0054; 
        10'b0010101111: data <= 15'h0040; 
        10'b0010110000: data <= 15'h0062; 
        10'b0010110001: data <= 15'h0050; 
        10'b0010110010: data <= 15'h0047; 
        10'b0010110011: data <= 15'h0044; 
        10'b0010110100: data <= 15'h005b; 
        10'b0010110101: data <= 15'h0082; 
        10'b0010110110: data <= 15'h005a; 
        10'b0010110111: data <= 15'h0021; 
        10'b0010111000: data <= 15'h0056; 
        10'b0010111001: data <= 15'h004f; 
        10'b0010111010: data <= 15'h004b; 
        10'b0010111011: data <= 15'h7fde; 
        10'b0010111100: data <= 15'h0020; 
        10'b0010111101: data <= 15'h7fe0; 
        10'b0010111110: data <= 15'h7f8e; 
        10'b0010111111: data <= 15'h7f8e; 
        10'b0011000000: data <= 15'h7fba; 
        10'b0011000001: data <= 15'h7ff2; 
        10'b0011000010: data <= 15'h7ffd; 
        10'b0011000011: data <= 15'h7ff5; 
        10'b0011000100: data <= 15'h0001; 
        10'b0011000101: data <= 15'h7ffc; 
        10'b0011000110: data <= 15'h0007; 
        10'b0011000111: data <= 15'h0031; 
        10'b0011001000: data <= 15'h0082; 
        10'b0011001001: data <= 15'h0081; 
        10'b0011001010: data <= 15'h005b; 
        10'b0011001011: data <= 15'h001a; 
        10'b0011001100: data <= 15'h001b; 
        10'b0011001101: data <= 15'h003a; 
        10'b0011001110: data <= 15'h0012; 
        10'b0011001111: data <= 15'h001a; 
        10'b0011010000: data <= 15'h004c; 
        10'b0011010001: data <= 15'h0048; 
        10'b0011010010: data <= 15'h0078; 
        10'b0011010011: data <= 15'h0046; 
        10'b0011010100: data <= 15'h0016; 
        10'b0011010101: data <= 15'h003c; 
        10'b0011010110: data <= 15'h0032; 
        10'b0011010111: data <= 15'h0036; 
        10'b0011011000: data <= 15'h0037; 
        10'b0011011001: data <= 15'h0008; 
        10'b0011011010: data <= 15'h7fc9; 
        10'b0011011011: data <= 15'h7f80; 
        10'b0011011100: data <= 15'h7fa4; 
        10'b0011011101: data <= 15'h7fe8; 
        10'b0011011110: data <= 15'h7fe1; 
        10'b0011011111: data <= 15'h7fef; 
        10'b0011100000: data <= 15'h7ff4; 
        10'b0011100001: data <= 15'h7fed; 
        10'b0011100010: data <= 15'h0005; 
        10'b0011100011: data <= 15'h002e; 
        10'b0011100100: data <= 15'h006b; 
        10'b0011100101: data <= 15'h0066; 
        10'b0011100110: data <= 15'h004c; 
        10'b0011100111: data <= 15'h001f; 
        10'b0011101000: data <= 15'h0034; 
        10'b0011101001: data <= 15'h0019; 
        10'b0011101010: data <= 15'h0041; 
        10'b0011101011: data <= 15'h0015; 
        10'b0011101100: data <= 15'h0012; 
        10'b0011101101: data <= 15'h0020; 
        10'b0011101110: data <= 15'h0082; 
        10'b0011101111: data <= 15'h006c; 
        10'b0011110000: data <= 15'h0019; 
        10'b0011110001: data <= 15'h003c; 
        10'b0011110010: data <= 15'h0056; 
        10'b0011110011: data <= 15'h0038; 
        10'b0011110100: data <= 15'h0052; 
        10'b0011110101: data <= 15'h002a; 
        10'b0011110110: data <= 15'h7fea; 
        10'b0011110111: data <= 15'h7f89; 
        10'b0011111000: data <= 15'h7fa7; 
        10'b0011111001: data <= 15'h7fe0; 
        10'b0011111010: data <= 15'h7fe4; 
        10'b0011111011: data <= 15'h7fec; 
        10'b0011111100: data <= 15'h7ff0; 
        10'b0011111101: data <= 15'h7fe1; 
        10'b0011111110: data <= 15'h7ff6; 
        10'b0011111111: data <= 15'h0014; 
        10'b0100000000: data <= 15'h0037; 
        10'b0100000001: data <= 15'h0049; 
        10'b0100000010: data <= 15'h003d; 
        10'b0100000011: data <= 15'h000f; 
        10'b0100000100: data <= 15'h7ff8; 
        10'b0100000101: data <= 15'h7fc7; 
        10'b0100000110: data <= 15'h7f94; 
        10'b0100000111: data <= 15'h7f3a; 
        10'b0100001000: data <= 15'h7f5f; 
        10'b0100001001: data <= 15'h7feb; 
        10'b0100001010: data <= 15'h009b; 
        10'b0100001011: data <= 15'h00ee; 
        10'b0100001100: data <= 15'h0089; 
        10'b0100001101: data <= 15'h0050; 
        10'b0100001110: data <= 15'h0057; 
        10'b0100001111: data <= 15'h0051; 
        10'b0100010000: data <= 15'h0079; 
        10'b0100010001: data <= 15'h004d; 
        10'b0100010010: data <= 15'h7fe9; 
        10'b0100010011: data <= 15'h7f8a; 
        10'b0100010100: data <= 15'h7fc5; 
        10'b0100010101: data <= 15'h7fdf; 
        10'b0100010110: data <= 15'h7fe7; 
        10'b0100010111: data <= 15'h7feb; 
        10'b0100011000: data <= 15'h7ffd; 
        10'b0100011001: data <= 15'h7ffb; 
        10'b0100011010: data <= 15'h0002; 
        10'b0100011011: data <= 15'h001e; 
        10'b0100011100: data <= 15'h001b; 
        10'b0100011101: data <= 15'h000b; 
        10'b0100011110: data <= 15'h7fdd; 
        10'b0100011111: data <= 15'h7fa8; 
        10'b0100100000: data <= 15'h7f60; 
        10'b0100100001: data <= 15'h7f1b; 
        10'b0100100010: data <= 15'h7ee7; 
        10'b0100100011: data <= 15'h7ee0; 
        10'b0100100100: data <= 15'h7f2c; 
        10'b0100100101: data <= 15'h7fca; 
        10'b0100100110: data <= 15'h007f; 
        10'b0100100111: data <= 15'h0093; 
        10'b0100101000: data <= 15'h007d; 
        10'b0100101001: data <= 15'h0074; 
        10'b0100101010: data <= 15'h0048; 
        10'b0100101011: data <= 15'h007d; 
        10'b0100101100: data <= 15'h0074; 
        10'b0100101101: data <= 15'h002e; 
        10'b0100101110: data <= 15'h7fd6; 
        10'b0100101111: data <= 15'h7fb3; 
        10'b0100110000: data <= 15'h7fe3; 
        10'b0100110001: data <= 15'h7fe0; 
        10'b0100110010: data <= 15'h7ff2; 
        10'b0100110011: data <= 15'h7ffd; 
        10'b0100110100: data <= 15'h0004; 
        10'b0100110101: data <= 15'h7ffd; 
        10'b0100110110: data <= 15'h7fe5; 
        10'b0100110111: data <= 15'h001d; 
        10'b0100111000: data <= 15'h7fef; 
        10'b0100111001: data <= 15'h7fa6; 
        10'b0100111010: data <= 15'h7f79; 
        10'b0100111011: data <= 15'h7f3a; 
        10'b0100111100: data <= 15'h7f08; 
        10'b0100111101: data <= 15'h7f2a; 
        10'b0100111110: data <= 15'h7f5d; 
        10'b0100111111: data <= 15'h7fb3; 
        10'b0101000000: data <= 15'h7fd6; 
        10'b0101000001: data <= 15'h0036; 
        10'b0101000010: data <= 15'h0054; 
        10'b0101000011: data <= 15'h0055; 
        10'b0101000100: data <= 15'h0027; 
        10'b0101000101: data <= 15'h0058; 
        10'b0101000110: data <= 15'h006d; 
        10'b0101000111: data <= 15'h006a; 
        10'b0101001000: data <= 15'h005d; 
        10'b0101001001: data <= 15'h0000; 
        10'b0101001010: data <= 15'h7fd7; 
        10'b0101001011: data <= 15'h7fde; 
        10'b0101001100: data <= 15'h7fe2; 
        10'b0101001101: data <= 15'h7fee; 
        10'b0101001110: data <= 15'h7fe7; 
        10'b0101001111: data <= 15'h7fe4; 
        10'b0101010000: data <= 15'h0001; 
        10'b0101010001: data <= 15'h7feb; 
        10'b0101010010: data <= 15'h7ffb; 
        10'b0101010011: data <= 15'h7ffe; 
        10'b0101010100: data <= 15'h7fdf; 
        10'b0101010101: data <= 15'h7fa6; 
        10'b0101010110: data <= 15'h7f62; 
        10'b0101010111: data <= 15'h7f3a; 
        10'b0101011000: data <= 15'h7f4d; 
        10'b0101011001: data <= 15'h7fa1; 
        10'b0101011010: data <= 15'h0002; 
        10'b0101011011: data <= 15'h0010; 
        10'b0101011100: data <= 15'h0019; 
        10'b0101011101: data <= 15'h0039; 
        10'b0101011110: data <= 15'h008d; 
        10'b0101011111: data <= 15'h0049; 
        10'b0101100000: data <= 15'h0032; 
        10'b0101100001: data <= 15'h0047; 
        10'b0101100010: data <= 15'h0039; 
        10'b0101100011: data <= 15'h7ffb; 
        10'b0101100100: data <= 15'h7fb7; 
        10'b0101100101: data <= 15'h7f9b; 
        10'b0101100110: data <= 15'h7f97; 
        10'b0101100111: data <= 15'h7fbd; 
        10'b0101101000: data <= 15'h7ff4; 
        10'b0101101001: data <= 15'h7fec; 
        10'b0101101010: data <= 15'h7ff5; 
        10'b0101101011: data <= 15'h7ff8; 
        10'b0101101100: data <= 15'h7ff2; 
        10'b0101101101: data <= 15'h7fea; 
        10'b0101101110: data <= 15'h7ff3; 
        10'b0101101111: data <= 15'h7ff7; 
        10'b0101110000: data <= 15'h7fd6; 
        10'b0101110001: data <= 15'h7fc2; 
        10'b0101110010: data <= 15'h7f80; 
        10'b0101110011: data <= 15'h7f6c; 
        10'b0101110100: data <= 15'h7f9b; 
        10'b0101110101: data <= 15'h7fec; 
        10'b0101110110: data <= 15'h7fdf; 
        10'b0101110111: data <= 15'h7fab; 
        10'b0101111000: data <= 15'h0007; 
        10'b0101111001: data <= 15'h007a; 
        10'b0101111010: data <= 15'h007b; 
        10'b0101111011: data <= 15'h0016; 
        10'b0101111100: data <= 15'h0038; 
        10'b0101111101: data <= 15'h003b; 
        10'b0101111110: data <= 15'h0020; 
        10'b0101111111: data <= 15'h7fd6; 
        10'b0110000000: data <= 15'h7f90; 
        10'b0110000001: data <= 15'h7f8f; 
        10'b0110000010: data <= 15'h7fa7; 
        10'b0110000011: data <= 15'h7fc1; 
        10'b0110000100: data <= 15'h7fdc; 
        10'b0110000101: data <= 15'h7fff; 
        10'b0110000110: data <= 15'h7ff9; 
        10'b0110000111: data <= 15'h7fed; 
        10'b0110001000: data <= 15'h0003; 
        10'b0110001001: data <= 15'h7fe8; 
        10'b0110001010: data <= 15'h7ff0; 
        10'b0110001011: data <= 15'h7ff6; 
        10'b0110001100: data <= 15'h7ff8; 
        10'b0110001101: data <= 15'h7fcc; 
        10'b0110001110: data <= 15'h7f8c; 
        10'b0110001111: data <= 15'h7f97; 
        10'b0110010000: data <= 15'h7fb9; 
        10'b0110010001: data <= 15'h7ff6; 
        10'b0110010010: data <= 15'h7fb5; 
        10'b0110010011: data <= 15'h7fb0; 
        10'b0110010100: data <= 15'h0017; 
        10'b0110010101: data <= 15'h003b; 
        10'b0110010110: data <= 15'h003f; 
        10'b0110010111: data <= 15'h7ff7; 
        10'b0110011000: data <= 15'h7fe6; 
        10'b0110011001: data <= 15'h7fed; 
        10'b0110011010: data <= 15'h0009; 
        10'b0110011011: data <= 15'h7fcf; 
        10'b0110011100: data <= 15'h7fbe; 
        10'b0110011101: data <= 15'h7fe0; 
        10'b0110011110: data <= 15'h7fd3; 
        10'b0110011111: data <= 15'h7fe1; 
        10'b0110100000: data <= 15'h7fd8; 
        10'b0110100001: data <= 15'h7fdc; 
        10'b0110100010: data <= 15'h0001; 
        10'b0110100011: data <= 15'h0002; 
        10'b0110100100: data <= 15'h0003; 
        10'b0110100101: data <= 15'h7fe8; 
        10'b0110100110: data <= 15'h0004; 
        10'b0110100111: data <= 15'h0009; 
        10'b0110101000: data <= 15'h7ff6; 
        10'b0110101001: data <= 15'h7fc6; 
        10'b0110101010: data <= 15'h7f94; 
        10'b0110101011: data <= 15'h7f8d; 
        10'b0110101100: data <= 15'h7faa; 
        10'b0110101101: data <= 15'h7fce; 
        10'b0110101110: data <= 15'h7fc8; 
        10'b0110101111: data <= 15'h7fed; 
        10'b0110110000: data <= 15'h0017; 
        10'b0110110001: data <= 15'h0060; 
        10'b0110110010: data <= 15'h0037; 
        10'b0110110011: data <= 15'h7ffb; 
        10'b0110110100: data <= 15'h7fb0; 
        10'b0110110101: data <= 15'h7fe9; 
        10'b0110110110: data <= 15'h7ff8; 
        10'b0110110111: data <= 15'h0015; 
        10'b0110111000: data <= 15'h0032; 
        10'b0110111001: data <= 15'h0030; 
        10'b0110111010: data <= 15'h0011; 
        10'b0110111011: data <= 15'h0006; 
        10'b0110111100: data <= 15'h7fe2; 
        10'b0110111101: data <= 15'h7ff9; 
        10'b0110111110: data <= 15'h7ff6; 
        10'b0110111111: data <= 15'h7fe8; 
        10'b0111000000: data <= 15'h7ff7; 
        10'b0111000001: data <= 15'h7ffb; 
        10'b0111000010: data <= 15'h0016; 
        10'b0111000011: data <= 15'h0004; 
        10'b0111000100: data <= 15'h0010; 
        10'b0111000101: data <= 15'h7fe5; 
        10'b0111000110: data <= 15'h7fd4; 
        10'b0111000111: data <= 15'h7fb4; 
        10'b0111001000: data <= 15'h7f5a; 
        10'b0111001001: data <= 15'h7f52; 
        10'b0111001010: data <= 15'h7f65; 
        10'b0111001011: data <= 15'h7fd9; 
        10'b0111001100: data <= 15'h002e; 
        10'b0111001101: data <= 15'h0077; 
        10'b0111001110: data <= 15'h7ff3; 
        10'b0111001111: data <= 15'h7fa9; 
        10'b0111010000: data <= 15'h7fa4; 
        10'b0111010001: data <= 15'h7fe2; 
        10'b0111010010: data <= 15'h0027; 
        10'b0111010011: data <= 15'h0066; 
        10'b0111010100: data <= 15'h0048; 
        10'b0111010101: data <= 15'h005a; 
        10'b0111010110: data <= 15'h0058; 
        10'b0111010111: data <= 15'h0027; 
        10'b0111011000: data <= 15'h7ff5; 
        10'b0111011001: data <= 15'h7ff8; 
        10'b0111011010: data <= 15'h7fff; 
        10'b0111011011: data <= 15'h7ffd; 
        10'b0111011100: data <= 15'h7ffc; 
        10'b0111011101: data <= 15'h0004; 
        10'b0111011110: data <= 15'h0000; 
        10'b0111011111: data <= 15'h0038; 
        10'b0111100000: data <= 15'h001f; 
        10'b0111100001: data <= 15'h000a; 
        10'b0111100010: data <= 15'h7fe2; 
        10'b0111100011: data <= 15'h7f9c; 
        10'b0111100100: data <= 15'h7f4d; 
        10'b0111100101: data <= 15'h7ee4; 
        10'b0111100110: data <= 15'h7e9f; 
        10'b0111100111: data <= 15'h7ebe; 
        10'b0111101000: data <= 15'h7f0b; 
        10'b0111101001: data <= 15'h7f75; 
        10'b0111101010: data <= 15'h7f7f; 
        10'b0111101011: data <= 15'h7f8d; 
        10'b0111101100: data <= 15'h7ffb; 
        10'b0111101101: data <= 15'h0024; 
        10'b0111101110: data <= 15'h0041; 
        10'b0111101111: data <= 15'h0067; 
        10'b0111110000: data <= 15'h0015; 
        10'b0111110001: data <= 15'h007d; 
        10'b0111110010: data <= 15'h007d; 
        10'b0111110011: data <= 15'h0026; 
        10'b0111110100: data <= 15'h7fee; 
        10'b0111110101: data <= 15'h7fe5; 
        10'b0111110110: data <= 15'h7fe8; 
        10'b0111110111: data <= 15'h7fea; 
        10'b0111111000: data <= 15'h7ff2; 
        10'b0111111001: data <= 15'h7ff3; 
        10'b0111111010: data <= 15'h000b; 
        10'b0111111011: data <= 15'h0053; 
        10'b0111111100: data <= 15'h003b; 
        10'b0111111101: data <= 15'h0024; 
        10'b0111111110: data <= 15'h0013; 
        10'b0111111111: data <= 15'h7fea; 
        10'b1000000000: data <= 15'h7fc0; 
        10'b1000000001: data <= 15'h7f30; 
        10'b1000000010: data <= 15'h7ece; 
        10'b1000000011: data <= 15'h7edf; 
        10'b1000000100: data <= 15'h7ea3; 
        10'b1000000101: data <= 15'h7ee3; 
        10'b1000000110: data <= 15'h7f4c; 
        10'b1000000111: data <= 15'h7fd7; 
        10'b1000001000: data <= 15'h0049; 
        10'b1000001001: data <= 15'h0062; 
        10'b1000001010: data <= 15'h006a; 
        10'b1000001011: data <= 15'h0069; 
        10'b1000001100: data <= 15'h0049; 
        10'b1000001101: data <= 15'h0092; 
        10'b1000001110: data <= 15'h0088; 
        10'b1000001111: data <= 15'h0034; 
        10'b1000010000: data <= 15'h7fd0; 
        10'b1000010001: data <= 15'h7fe0; 
        10'b1000010010: data <= 15'h7fe8; 
        10'b1000010011: data <= 15'h7ffc; 
        10'b1000010100: data <= 15'h7ffc; 
        10'b1000010101: data <= 15'h7fe8; 
        10'b1000010110: data <= 15'h7ff1; 
        10'b1000010111: data <= 15'h0068; 
        10'b1000011000: data <= 15'h006a; 
        10'b1000011001: data <= 15'h007c; 
        10'b1000011010: data <= 15'h006b; 
        10'b1000011011: data <= 15'h0027; 
        10'b1000011100: data <= 15'h000c; 
        10'b1000011101: data <= 15'h7fd4; 
        10'b1000011110: data <= 15'h7fe1; 
        10'b1000011111: data <= 15'h7f9d; 
        10'b1000100000: data <= 15'h7f70; 
        10'b1000100001: data <= 15'h7f67; 
        10'b1000100010: data <= 15'h7f98; 
        10'b1000100011: data <= 15'h0025; 
        10'b1000100100: data <= 15'h0063; 
        10'b1000100101: data <= 15'h007b; 
        10'b1000100110: data <= 15'h008a; 
        10'b1000100111: data <= 15'h007b; 
        10'b1000101000: data <= 15'h006d; 
        10'b1000101001: data <= 15'h0080; 
        10'b1000101010: data <= 15'h0031; 
        10'b1000101011: data <= 15'h0006; 
        10'b1000101100: data <= 15'h7fd7; 
        10'b1000101101: data <= 15'h7ff9; 
        10'b1000101110: data <= 15'h7ffc; 
        10'b1000101111: data <= 15'h7ff7; 
        10'b1000110000: data <= 15'h7ffb; 
        10'b1000110001: data <= 15'h7fe1; 
        10'b1000110010: data <= 15'h0013; 
        10'b1000110011: data <= 15'h006f; 
        10'b1000110100: data <= 15'h0089; 
        10'b1000110101: data <= 15'h0094; 
        10'b1000110110: data <= 15'h009c; 
        10'b1000110111: data <= 15'h004f; 
        10'b1000111000: data <= 15'h005d; 
        10'b1000111001: data <= 15'h0069; 
        10'b1000111010: data <= 15'h0027; 
        10'b1000111011: data <= 15'h7ff5; 
        10'b1000111100: data <= 15'h7fdd; 
        10'b1000111101: data <= 15'h7fca; 
        10'b1000111110: data <= 15'h0010; 
        10'b1000111111: data <= 15'h001d; 
        10'b1001000000: data <= 15'h0038; 
        10'b1001000001: data <= 15'h0063; 
        10'b1001000010: data <= 15'h0068; 
        10'b1001000011: data <= 15'h0047; 
        10'b1001000100: data <= 15'h007b; 
        10'b1001000101: data <= 15'h0046; 
        10'b1001000110: data <= 15'h7ff3; 
        10'b1001000111: data <= 15'h7fe4; 
        10'b1001001000: data <= 15'h7fe0; 
        10'b1001001001: data <= 15'h7ff6; 
        10'b1001001010: data <= 15'h7ff6; 
        10'b1001001011: data <= 15'h7ff5; 
        10'b1001001100: data <= 15'h7feb; 
        10'b1001001101: data <= 15'h7fff; 
        10'b1001001110: data <= 15'h7ff8; 
        10'b1001001111: data <= 15'h0037; 
        10'b1001010000: data <= 15'h0084; 
        10'b1001010001: data <= 15'h0084; 
        10'b1001010010: data <= 15'h0073; 
        10'b1001010011: data <= 15'h0041; 
        10'b1001010100: data <= 15'h0045; 
        10'b1001010101: data <= 15'h0017; 
        10'b1001010110: data <= 15'h7ff7; 
        10'b1001010111: data <= 15'h7fe1; 
        10'b1001011000: data <= 15'h000a; 
        10'b1001011001: data <= 15'h7ffa; 
        10'b1001011010: data <= 15'h7ff8; 
        10'b1001011011: data <= 15'h7ff1; 
        10'b1001011100: data <= 15'h0020; 
        10'b1001011101: data <= 15'h000c; 
        10'b1001011110: data <= 15'h003f; 
        10'b1001011111: data <= 15'h0066; 
        10'b1001100000: data <= 15'h003b; 
        10'b1001100001: data <= 15'h0017; 
        10'b1001100010: data <= 15'h7fe9; 
        10'b1001100011: data <= 15'h7fc5; 
        10'b1001100100: data <= 15'h7fed; 
        10'b1001100101: data <= 15'h7fe8; 
        10'b1001100110: data <= 15'h7fe0; 
        10'b1001100111: data <= 15'h7fe2; 
        10'b1001101000: data <= 15'h7ff3; 
        10'b1001101001: data <= 15'h7ff7; 
        10'b1001101010: data <= 15'h7ffa; 
        10'b1001101011: data <= 15'h0022; 
        10'b1001101100: data <= 15'h0042; 
        10'b1001101101: data <= 15'h005a; 
        10'b1001101110: data <= 15'h0050; 
        10'b1001101111: data <= 15'h002e; 
        10'b1001110000: data <= 15'h0004; 
        10'b1001110001: data <= 15'h0021; 
        10'b1001110010: data <= 15'h0028; 
        10'b1001110011: data <= 15'h0031; 
        10'b1001110100: data <= 15'h000d; 
        10'b1001110101: data <= 15'h7fee; 
        10'b1001110110: data <= 15'h7fed; 
        10'b1001110111: data <= 15'h7fe5; 
        10'b1001111000: data <= 15'h0015; 
        10'b1001111001: data <= 15'h0010; 
        10'b1001111010: data <= 15'h0010; 
        10'b1001111011: data <= 15'h0046; 
        10'b1001111100: data <= 15'h0022; 
        10'b1001111101: data <= 15'h7ff4; 
        10'b1001111110: data <= 15'h7ff0; 
        10'b1001111111: data <= 15'h7feb; 
        10'b1010000000: data <= 15'h7fd3; 
        10'b1010000001: data <= 15'h7fde; 
        10'b1010000010: data <= 15'h7ffa; 
        10'b1010000011: data <= 15'h7fff; 
        10'b1010000100: data <= 15'h7ff7; 
        10'b1010000101: data <= 15'h7fe7; 
        10'b1010000110: data <= 15'h7feb; 
        10'b1010000111: data <= 15'h0017; 
        10'b1010001000: data <= 15'h0048; 
        10'b1010001001: data <= 15'h006d; 
        10'b1010001010: data <= 15'h0051; 
        10'b1010001011: data <= 15'h0056; 
        10'b1010001100: data <= 15'h0015; 
        10'b1010001101: data <= 15'h0037; 
        10'b1010001110: data <= 15'h0023; 
        10'b1010001111: data <= 15'h7fff; 
        10'b1010010000: data <= 15'h7fe4; 
        10'b1010010001: data <= 15'h0004; 
        10'b1010010010: data <= 15'h000b; 
        10'b1010010011: data <= 15'h001c; 
        10'b1010010100: data <= 15'h0014; 
        10'b1010010101: data <= 15'h002b; 
        10'b1010010110: data <= 15'h0044; 
        10'b1010010111: data <= 15'h7ff5; 
        10'b1010011000: data <= 15'h7fd3; 
        10'b1010011001: data <= 15'h7fd3; 
        10'b1010011010: data <= 15'h7fe8; 
        10'b1010011011: data <= 15'h7fe2; 
        10'b1010011100: data <= 15'h7ffd; 
        10'b1010011101: data <= 15'h7ff8; 
        10'b1010011110: data <= 15'h7fe4; 
        10'b1010011111: data <= 15'h7fe6; 
        10'b1010100000: data <= 15'h7fec; 
        10'b1010100001: data <= 15'h0003; 
        10'b1010100010: data <= 15'h0003; 
        10'b1010100011: data <= 15'h0000; 
        10'b1010100100: data <= 15'h002e; 
        10'b1010100101: data <= 15'h004b; 
        10'b1010100110: data <= 15'h0058; 
        10'b1010100111: data <= 15'h0068; 
        10'b1010101000: data <= 15'h006a; 
        10'b1010101001: data <= 15'h0057; 
        10'b1010101010: data <= 15'h007e; 
        10'b1010101011: data <= 15'h0085; 
        10'b1010101100: data <= 15'h0089; 
        10'b1010101101: data <= 15'h006c; 
        10'b1010101110: data <= 15'h005f; 
        10'b1010101111: data <= 15'h0046; 
        10'b1010110000: data <= 15'h0043; 
        10'b1010110001: data <= 15'h7ffa; 
        10'b1010110010: data <= 15'h7fca; 
        10'b1010110011: data <= 15'h7fb5; 
        10'b1010110100: data <= 15'h7fbc; 
        10'b1010110101: data <= 15'h7fd7; 
        10'b1010110110: data <= 15'h7fd9; 
        10'b1010110111: data <= 15'h7ff5; 
        10'b1010111000: data <= 15'h7fed; 
        10'b1010111001: data <= 15'h0000; 
        10'b1010111010: data <= 15'h7fec; 
        10'b1010111011: data <= 15'h0004; 
        10'b1010111100: data <= 15'h7ffd; 
        10'b1010111101: data <= 15'h7fe0; 
        10'b1010111110: data <= 15'h0002; 
        10'b1010111111: data <= 15'h0005; 
        10'b1011000000: data <= 15'h7ff8; 
        10'b1011000001: data <= 15'h001d; 
        10'b1011000010: data <= 15'h002c; 
        10'b1011000011: data <= 15'h0019; 
        10'b1011000100: data <= 15'h003b; 
        10'b1011000101: data <= 15'h003c; 
        10'b1011000110: data <= 15'h0070; 
        10'b1011000111: data <= 15'h0080; 
        10'b1011001000: data <= 15'h0089; 
        10'b1011001001: data <= 15'h006c; 
        10'b1011001010: data <= 15'h004c; 
        10'b1011001011: data <= 15'h001f; 
        10'b1011001100: data <= 15'h7ff4; 
        10'b1011001101: data <= 15'h7fd0; 
        10'b1011001110: data <= 15'h7fcf; 
        10'b1011001111: data <= 15'h7fd8; 
        10'b1011010000: data <= 15'h7fd8; 
        10'b1011010001: data <= 15'h7fec; 
        10'b1011010010: data <= 15'h7fec; 
        10'b1011010011: data <= 15'h7ffe; 
        10'b1011010100: data <= 15'h7fe8; 
        10'b1011010101: data <= 15'h0003; 
        10'b1011010110: data <= 15'h7fe0; 
        10'b1011010111: data <= 15'h7ffc; 
        10'b1011011000: data <= 15'h7fe9; 
        10'b1011011001: data <= 15'h7fdf; 
        10'b1011011010: data <= 15'h7fe1; 
        10'b1011011011: data <= 15'h7ff8; 
        10'b1011011100: data <= 15'h7ff8; 
        10'b1011011101: data <= 15'h7fea; 
        10'b1011011110: data <= 15'h7fe7; 
        10'b1011011111: data <= 15'h7ff7; 
        10'b1011100000: data <= 15'h7ff8; 
        10'b1011100001: data <= 15'h7ff6; 
        10'b1011100010: data <= 15'h7ff1; 
        10'b1011100011: data <= 15'h7ff4; 
        10'b1011100100: data <= 15'h7fee; 
        10'b1011100101: data <= 15'h7ff6; 
        10'b1011100110: data <= 15'h7fee; 
        10'b1011100111: data <= 15'h7fdd; 
        10'b1011101000: data <= 15'h7fea; 
        10'b1011101001: data <= 15'h7ff6; 
        10'b1011101010: data <= 15'h7ff2; 
        10'b1011101011: data <= 15'h7ff7; 
        10'b1011101100: data <= 15'h7fe1; 
        10'b1011101101: data <= 15'h7fe2; 
        10'b1011101110: data <= 15'h7ffb; 
        10'b1011101111: data <= 15'h7fef; 
        10'b1011110000: data <= 15'h0001; 
        10'b1011110001: data <= 15'h7fe8; 
        10'b1011110010: data <= 15'h7ffd; 
        10'b1011110011: data <= 15'h0004; 
        10'b1011110100: data <= 15'h7ff0; 
        10'b1011110101: data <= 15'h7fe8; 
        10'b1011110110: data <= 15'h7ff5; 
        10'b1011110111: data <= 15'h7fe1; 
        10'b1011111000: data <= 15'h0002; 
        10'b1011111001: data <= 15'h7ff8; 
        10'b1011111010: data <= 15'h7ffe; 
        10'b1011111011: data <= 15'h7ff6; 
        10'b1011111100: data <= 15'h7ffb; 
        10'b1011111101: data <= 15'h7fe1; 
        10'b1011111110: data <= 15'h7fe7; 
        10'b1011111111: data <= 15'h7ff9; 
        10'b1100000000: data <= 15'h7fe6; 
        10'b1100000001: data <= 15'h7ffb; 
        10'b1100000010: data <= 15'h7fed; 
        10'b1100000011: data <= 15'h7ff5; 
        10'b1100000100: data <= 15'h7fee; 
        10'b1100000101: data <= 15'h7fff; 
        10'b1100000110: data <= 15'h7fe3; 
        10'b1100000111: data <= 15'h7fe8; 
        10'b1100001000: data <= 15'h7ffe; 
        10'b1100001001: data <= 15'h7ff5; 
        10'b1100001010: data <= 15'h7fe7; 
        10'b1100001011: data <= 15'h7ff8; 
        10'b1100001100: data <= 15'h7fe3; 
        10'b1100001101: data <= 15'h7fe1; 
        10'b1100001110: data <= 15'h7ffe; 
        10'b1100001111: data <= 15'h7ff1; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 10) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 16'hffec; 
        10'b0000000001: data <= 16'hffce; 
        10'b0000000010: data <= 16'hfffe; 
        10'b0000000011: data <= 16'h0002; 
        10'b0000000100: data <= 16'h0005; 
        10'b0000000101: data <= 16'hfffc; 
        10'b0000000110: data <= 16'hffed; 
        10'b0000000111: data <= 16'h0005; 
        10'b0000001000: data <= 16'hffd8; 
        10'b0000001001: data <= 16'h0003; 
        10'b0000001010: data <= 16'h0003; 
        10'b0000001011: data <= 16'hffde; 
        10'b0000001100: data <= 16'hffdd; 
        10'b0000001101: data <= 16'hffdc; 
        10'b0000001110: data <= 16'hffdf; 
        10'b0000001111: data <= 16'hffe3; 
        10'b0000010000: data <= 16'h0001; 
        10'b0000010001: data <= 16'h0002; 
        10'b0000010010: data <= 16'hffce; 
        10'b0000010011: data <= 16'h0005; 
        10'b0000010100: data <= 16'hfff0; 
        10'b0000010101: data <= 16'hfff2; 
        10'b0000010110: data <= 16'hffbf; 
        10'b0000010111: data <= 16'hfffc; 
        10'b0000011000: data <= 16'hfffe; 
        10'b0000011001: data <= 16'hffc3; 
        10'b0000011010: data <= 16'hffe2; 
        10'b0000011011: data <= 16'h0002; 
        10'b0000011100: data <= 16'hffcd; 
        10'b0000011101: data <= 16'hffe0; 
        10'b0000011110: data <= 16'hffcd; 
        10'b0000011111: data <= 16'hffee; 
        10'b0000100000: data <= 16'hffc6; 
        10'b0000100001: data <= 16'hffe4; 
        10'b0000100010: data <= 16'h0007; 
        10'b0000100011: data <= 16'h0004; 
        10'b0000100100: data <= 16'hffc2; 
        10'b0000100101: data <= 16'hffbf; 
        10'b0000100110: data <= 16'hffc6; 
        10'b0000100111: data <= 16'hffed; 
        10'b0000101000: data <= 16'hfff2; 
        10'b0000101001: data <= 16'hffe2; 
        10'b0000101010: data <= 16'hffdd; 
        10'b0000101011: data <= 16'hffd2; 
        10'b0000101100: data <= 16'h0006; 
        10'b0000101101: data <= 16'hffce; 
        10'b0000101110: data <= 16'hfff5; 
        10'b0000101111: data <= 16'hffda; 
        10'b0000110000: data <= 16'hffdb; 
        10'b0000110001: data <= 16'hffc4; 
        10'b0000110010: data <= 16'hffe7; 
        10'b0000110011: data <= 16'hfffa; 
        10'b0000110100: data <= 16'hffca; 
        10'b0000110101: data <= 16'hfffd; 
        10'b0000110110: data <= 16'hffeb; 
        10'b0000110111: data <= 16'hffca; 
        10'b0000111000: data <= 16'hffd3; 
        10'b0000111001: data <= 16'hffe7; 
        10'b0000111010: data <= 16'hffe5; 
        10'b0000111011: data <= 16'hffce; 
        10'b0000111100: data <= 16'hfff0; 
        10'b0000111101: data <= 16'hfff5; 
        10'b0000111110: data <= 16'hffd6; 
        10'b0000111111: data <= 16'hfff5; 
        10'b0001000000: data <= 16'hfffa; 
        10'b0001000001: data <= 16'hffe2; 
        10'b0001000010: data <= 16'hffc9; 
        10'b0001000011: data <= 16'hffca; 
        10'b0001000100: data <= 16'hffc3; 
        10'b0001000101: data <= 16'hffcc; 
        10'b0001000110: data <= 16'hffdf; 
        10'b0001000111: data <= 16'hffda; 
        10'b0001001000: data <= 16'hffd5; 
        10'b0001001001: data <= 16'hffd3; 
        10'b0001001010: data <= 16'hfff5; 
        10'b0001001011: data <= 16'hffff; 
        10'b0001001100: data <= 16'hffe1; 
        10'b0001001101: data <= 16'hffcd; 
        10'b0001001110: data <= 16'h0006; 
        10'b0001001111: data <= 16'hfffc; 
        10'b0001010000: data <= 16'h0000; 
        10'b0001010001: data <= 16'hffd8; 
        10'b0001010010: data <= 16'hffc1; 
        10'b0001010011: data <= 16'hffe3; 
        10'b0001010100: data <= 16'h0007; 
        10'b0001010101: data <= 16'hfff4; 
        10'b0001010110: data <= 16'hffe4; 
        10'b0001010111: data <= 16'hfff8; 
        10'b0001011000: data <= 16'hfff3; 
        10'b0001011001: data <= 16'h0000; 
        10'b0001011010: data <= 16'hffed; 
        10'b0001011011: data <= 16'hfffc; 
        10'b0001011100: data <= 16'hfff9; 
        10'b0001011101: data <= 16'hffe8; 
        10'b0001011110: data <= 16'h0016; 
        10'b0001011111: data <= 16'h004a; 
        10'b0001100000: data <= 16'h009c; 
        10'b0001100001: data <= 16'h0082; 
        10'b0001100010: data <= 16'h0084; 
        10'b0001100011: data <= 16'h0092; 
        10'b0001100100: data <= 16'h0065; 
        10'b0001100101: data <= 16'h0072; 
        10'b0001100110: data <= 16'h0059; 
        10'b0001100111: data <= 16'h0007; 
        10'b0001101000: data <= 16'hfff7; 
        10'b0001101001: data <= 16'hff93; 
        10'b0001101010: data <= 16'hffc1; 
        10'b0001101011: data <= 16'hfffb; 
        10'b0001101100: data <= 16'h0003; 
        10'b0001101101: data <= 16'hffd0; 
        10'b0001101110: data <= 16'hffea; 
        10'b0001101111: data <= 16'hffd6; 
        10'b0001110000: data <= 16'hffea; 
        10'b0001110001: data <= 16'hfffc; 
        10'b0001110010: data <= 16'hffef; 
        10'b0001110011: data <= 16'h0002; 
        10'b0001110100: data <= 16'h0018; 
        10'b0001110101: data <= 16'h0000; 
        10'b0001110110: data <= 16'h005c; 
        10'b0001110111: data <= 16'h004e; 
        10'b0001111000: data <= 16'h00d4; 
        10'b0001111001: data <= 16'h00b6; 
        10'b0001111010: data <= 16'h00e1; 
        10'b0001111011: data <= 16'h010f; 
        10'b0001111100: data <= 16'h013a; 
        10'b0001111101: data <= 16'h0151; 
        10'b0001111110: data <= 16'h012f; 
        10'b0001111111: data <= 16'h00de; 
        10'b0010000000: data <= 16'h007d; 
        10'b0010000001: data <= 16'h0064; 
        10'b0010000010: data <= 16'h00a4; 
        10'b0010000011: data <= 16'h0014; 
        10'b0010000100: data <= 16'hff90; 
        10'b0010000101: data <= 16'hff51; 
        10'b0010000110: data <= 16'hff6a; 
        10'b0010000111: data <= 16'hff6e; 
        10'b0010001000: data <= 16'hffee; 
        10'b0010001001: data <= 16'hffe5; 
        10'b0010001010: data <= 16'hffda; 
        10'b0010001011: data <= 16'hfff6; 
        10'b0010001100: data <= 16'hffc9; 
        10'b0010001101: data <= 16'hffc1; 
        10'b0010001110: data <= 16'hffd1; 
        10'b0010001111: data <= 16'hffd1; 
        10'b0010010000: data <= 16'h000c; 
        10'b0010010001: data <= 16'h0060; 
        10'b0010010010: data <= 16'h00af; 
        10'b0010010011: data <= 16'h008c; 
        10'b0010010100: data <= 16'h00a0; 
        10'b0010010101: data <= 16'h008d; 
        10'b0010010110: data <= 16'h0080; 
        10'b0010010111: data <= 16'h00a6; 
        10'b0010011000: data <= 16'h00a9; 
        10'b0010011001: data <= 16'h00ca; 
        10'b0010011010: data <= 16'h0023; 
        10'b0010011011: data <= 16'h0087; 
        10'b0010011100: data <= 16'h009c; 
        10'b0010011101: data <= 16'hfff4; 
        10'b0010011110: data <= 16'hfff8; 
        10'b0010011111: data <= 16'hffb9; 
        10'b0010100000: data <= 16'hff9e; 
        10'b0010100001: data <= 16'hff30; 
        10'b0010100010: data <= 16'hfef6; 
        10'b0010100011: data <= 16'hff1f; 
        10'b0010100100: data <= 16'hffbf; 
        10'b0010100101: data <= 16'h0000; 
        10'b0010100110: data <= 16'hffd3; 
        10'b0010100111: data <= 16'hffe4; 
        10'b0010101000: data <= 16'hffcf; 
        10'b0010101001: data <= 16'hffd9; 
        10'b0010101010: data <= 16'hffd5; 
        10'b0010101011: data <= 16'h0014; 
        10'b0010101100: data <= 16'h0076; 
        10'b0010101101: data <= 16'h00dc; 
        10'b0010101110: data <= 16'h00a8; 
        10'b0010101111: data <= 16'h0081; 
        10'b0010110000: data <= 16'h00c3; 
        10'b0010110001: data <= 16'h009f; 
        10'b0010110010: data <= 16'h008e; 
        10'b0010110011: data <= 16'h0087; 
        10'b0010110100: data <= 16'h00b5; 
        10'b0010110101: data <= 16'h0104; 
        10'b0010110110: data <= 16'h00b5; 
        10'b0010110111: data <= 16'h0041; 
        10'b0010111000: data <= 16'h00ac; 
        10'b0010111001: data <= 16'h009e; 
        10'b0010111010: data <= 16'h0096; 
        10'b0010111011: data <= 16'hffbd; 
        10'b0010111100: data <= 16'h0040; 
        10'b0010111101: data <= 16'hffc1; 
        10'b0010111110: data <= 16'hff1b; 
        10'b0010111111: data <= 16'hff1b; 
        10'b0011000000: data <= 16'hff74; 
        10'b0011000001: data <= 16'hffe4; 
        10'b0011000010: data <= 16'hfffa; 
        10'b0011000011: data <= 16'hffea; 
        10'b0011000100: data <= 16'h0003; 
        10'b0011000101: data <= 16'hfff8; 
        10'b0011000110: data <= 16'h000d; 
        10'b0011000111: data <= 16'h0063; 
        10'b0011001000: data <= 16'h0104; 
        10'b0011001001: data <= 16'h0102; 
        10'b0011001010: data <= 16'h00b6; 
        10'b0011001011: data <= 16'h0033; 
        10'b0011001100: data <= 16'h0037; 
        10'b0011001101: data <= 16'h0074; 
        10'b0011001110: data <= 16'h0024; 
        10'b0011001111: data <= 16'h0035; 
        10'b0011010000: data <= 16'h0098; 
        10'b0011010001: data <= 16'h0090; 
        10'b0011010010: data <= 16'h00ef; 
        10'b0011010011: data <= 16'h008c; 
        10'b0011010100: data <= 16'h002b; 
        10'b0011010101: data <= 16'h0078; 
        10'b0011010110: data <= 16'h0063; 
        10'b0011010111: data <= 16'h006c; 
        10'b0011011000: data <= 16'h006e; 
        10'b0011011001: data <= 16'h000f; 
        10'b0011011010: data <= 16'hff92; 
        10'b0011011011: data <= 16'hff00; 
        10'b0011011100: data <= 16'hff48; 
        10'b0011011101: data <= 16'hffd0; 
        10'b0011011110: data <= 16'hffc1; 
        10'b0011011111: data <= 16'hffde; 
        10'b0011100000: data <= 16'hffe8; 
        10'b0011100001: data <= 16'hffda; 
        10'b0011100010: data <= 16'h000b; 
        10'b0011100011: data <= 16'h005c; 
        10'b0011100100: data <= 16'h00d6; 
        10'b0011100101: data <= 16'h00cb; 
        10'b0011100110: data <= 16'h0099; 
        10'b0011100111: data <= 16'h003e; 
        10'b0011101000: data <= 16'h0068; 
        10'b0011101001: data <= 16'h0031; 
        10'b0011101010: data <= 16'h0083; 
        10'b0011101011: data <= 16'h002a; 
        10'b0011101100: data <= 16'h0024; 
        10'b0011101101: data <= 16'h0040; 
        10'b0011101110: data <= 16'h0104; 
        10'b0011101111: data <= 16'h00d8; 
        10'b0011110000: data <= 16'h0032; 
        10'b0011110001: data <= 16'h0078; 
        10'b0011110010: data <= 16'h00ac; 
        10'b0011110011: data <= 16'h0070; 
        10'b0011110100: data <= 16'h00a4; 
        10'b0011110101: data <= 16'h0055; 
        10'b0011110110: data <= 16'hffd4; 
        10'b0011110111: data <= 16'hff12; 
        10'b0011111000: data <= 16'hff4e; 
        10'b0011111001: data <= 16'hffbf; 
        10'b0011111010: data <= 16'hffc9; 
        10'b0011111011: data <= 16'hffd8; 
        10'b0011111100: data <= 16'hffe1; 
        10'b0011111101: data <= 16'hffc3; 
        10'b0011111110: data <= 16'hffed; 
        10'b0011111111: data <= 16'h0028; 
        10'b0100000000: data <= 16'h006f; 
        10'b0100000001: data <= 16'h0093; 
        10'b0100000010: data <= 16'h007a; 
        10'b0100000011: data <= 16'h001e; 
        10'b0100000100: data <= 16'hfff1; 
        10'b0100000101: data <= 16'hff8f; 
        10'b0100000110: data <= 16'hff28; 
        10'b0100000111: data <= 16'hfe73; 
        10'b0100001000: data <= 16'hfebe; 
        10'b0100001001: data <= 16'hffd5; 
        10'b0100001010: data <= 16'h0136; 
        10'b0100001011: data <= 16'h01dc; 
        10'b0100001100: data <= 16'h0113; 
        10'b0100001101: data <= 16'h00a1; 
        10'b0100001110: data <= 16'h00af; 
        10'b0100001111: data <= 16'h00a2; 
        10'b0100010000: data <= 16'h00f2; 
        10'b0100010001: data <= 16'h009a; 
        10'b0100010010: data <= 16'hffd1; 
        10'b0100010011: data <= 16'hff14; 
        10'b0100010100: data <= 16'hff89; 
        10'b0100010101: data <= 16'hffbd; 
        10'b0100010110: data <= 16'hffce; 
        10'b0100010111: data <= 16'hffd6; 
        10'b0100011000: data <= 16'hfff9; 
        10'b0100011001: data <= 16'hfff6; 
        10'b0100011010: data <= 16'h0003; 
        10'b0100011011: data <= 16'h003c; 
        10'b0100011100: data <= 16'h0036; 
        10'b0100011101: data <= 16'h0017; 
        10'b0100011110: data <= 16'hffbb; 
        10'b0100011111: data <= 16'hff51; 
        10'b0100100000: data <= 16'hfebf; 
        10'b0100100001: data <= 16'hfe36; 
        10'b0100100010: data <= 16'hfdce; 
        10'b0100100011: data <= 16'hfdc0; 
        10'b0100100100: data <= 16'hfe58; 
        10'b0100100101: data <= 16'hff95; 
        10'b0100100110: data <= 16'h00fe; 
        10'b0100100111: data <= 16'h0126; 
        10'b0100101000: data <= 16'h00fa; 
        10'b0100101001: data <= 16'h00e9; 
        10'b0100101010: data <= 16'h0090; 
        10'b0100101011: data <= 16'h00f9; 
        10'b0100101100: data <= 16'h00e8; 
        10'b0100101101: data <= 16'h005d; 
        10'b0100101110: data <= 16'hffad; 
        10'b0100101111: data <= 16'hff67; 
        10'b0100110000: data <= 16'hffc7; 
        10'b0100110001: data <= 16'hffbf; 
        10'b0100110010: data <= 16'hffe5; 
        10'b0100110011: data <= 16'hfff9; 
        10'b0100110100: data <= 16'h0008; 
        10'b0100110101: data <= 16'hfff9; 
        10'b0100110110: data <= 16'hffcb; 
        10'b0100110111: data <= 16'h003a; 
        10'b0100111000: data <= 16'hffde; 
        10'b0100111001: data <= 16'hff4c; 
        10'b0100111010: data <= 16'hfef2; 
        10'b0100111011: data <= 16'hfe74; 
        10'b0100111100: data <= 16'hfe11; 
        10'b0100111101: data <= 16'hfe54; 
        10'b0100111110: data <= 16'hfeba; 
        10'b0100111111: data <= 16'hff66; 
        10'b0101000000: data <= 16'hffad; 
        10'b0101000001: data <= 16'h006c; 
        10'b0101000010: data <= 16'h00a9; 
        10'b0101000011: data <= 16'h00aa; 
        10'b0101000100: data <= 16'h004e; 
        10'b0101000101: data <= 16'h00b0; 
        10'b0101000110: data <= 16'h00da; 
        10'b0101000111: data <= 16'h00d4; 
        10'b0101001000: data <= 16'h00b9; 
        10'b0101001001: data <= 16'h0001; 
        10'b0101001010: data <= 16'hffae; 
        10'b0101001011: data <= 16'hffbc; 
        10'b0101001100: data <= 16'hffc4; 
        10'b0101001101: data <= 16'hffdc; 
        10'b0101001110: data <= 16'hffcf; 
        10'b0101001111: data <= 16'hffc9; 
        10'b0101010000: data <= 16'h0002; 
        10'b0101010001: data <= 16'hffd6; 
        10'b0101010010: data <= 16'hfff5; 
        10'b0101010011: data <= 16'hfffd; 
        10'b0101010100: data <= 16'hffbf; 
        10'b0101010101: data <= 16'hff4c; 
        10'b0101010110: data <= 16'hfec4; 
        10'b0101010111: data <= 16'hfe75; 
        10'b0101011000: data <= 16'hfe9b; 
        10'b0101011001: data <= 16'hff42; 
        10'b0101011010: data <= 16'h0004; 
        10'b0101011011: data <= 16'h0020; 
        10'b0101011100: data <= 16'h0032; 
        10'b0101011101: data <= 16'h0072; 
        10'b0101011110: data <= 16'h011b; 
        10'b0101011111: data <= 16'h0092; 
        10'b0101100000: data <= 16'h0064; 
        10'b0101100001: data <= 16'h008d; 
        10'b0101100010: data <= 16'h0071; 
        10'b0101100011: data <= 16'hfff6; 
        10'b0101100100: data <= 16'hff6e; 
        10'b0101100101: data <= 16'hff37; 
        10'b0101100110: data <= 16'hff2e; 
        10'b0101100111: data <= 16'hff7a; 
        10'b0101101000: data <= 16'hffe8; 
        10'b0101101001: data <= 16'hffd7; 
        10'b0101101010: data <= 16'hffea; 
        10'b0101101011: data <= 16'hfff1; 
        10'b0101101100: data <= 16'hffe3; 
        10'b0101101101: data <= 16'hffd5; 
        10'b0101101110: data <= 16'hffe5; 
        10'b0101101111: data <= 16'hffee; 
        10'b0101110000: data <= 16'hffac; 
        10'b0101110001: data <= 16'hff85; 
        10'b0101110010: data <= 16'hfeff; 
        10'b0101110011: data <= 16'hfed7; 
        10'b0101110100: data <= 16'hff37; 
        10'b0101110101: data <= 16'hffd8; 
        10'b0101110110: data <= 16'hffbf; 
        10'b0101110111: data <= 16'hff55; 
        10'b0101111000: data <= 16'h000e; 
        10'b0101111001: data <= 16'h00f3; 
        10'b0101111010: data <= 16'h00f6; 
        10'b0101111011: data <= 16'h002d; 
        10'b0101111100: data <= 16'h0070; 
        10'b0101111101: data <= 16'h0077; 
        10'b0101111110: data <= 16'h003f; 
        10'b0101111111: data <= 16'hffac; 
        10'b0110000000: data <= 16'hff20; 
        10'b0110000001: data <= 16'hff1e; 
        10'b0110000010: data <= 16'hff4e; 
        10'b0110000011: data <= 16'hff83; 
        10'b0110000100: data <= 16'hffb8; 
        10'b0110000101: data <= 16'hfffe; 
        10'b0110000110: data <= 16'hfff3; 
        10'b0110000111: data <= 16'hffda; 
        10'b0110001000: data <= 16'h0006; 
        10'b0110001001: data <= 16'hffcf; 
        10'b0110001010: data <= 16'hffe1; 
        10'b0110001011: data <= 16'hffec; 
        10'b0110001100: data <= 16'hfff1; 
        10'b0110001101: data <= 16'hff99; 
        10'b0110001110: data <= 16'hff18; 
        10'b0110001111: data <= 16'hff2e; 
        10'b0110010000: data <= 16'hff72; 
        10'b0110010001: data <= 16'hffec; 
        10'b0110010010: data <= 16'hff6b; 
        10'b0110010011: data <= 16'hff61; 
        10'b0110010100: data <= 16'h002d; 
        10'b0110010101: data <= 16'h0076; 
        10'b0110010110: data <= 16'h007e; 
        10'b0110010111: data <= 16'hffed; 
        10'b0110011000: data <= 16'hffcd; 
        10'b0110011001: data <= 16'hffda; 
        10'b0110011010: data <= 16'h0011; 
        10'b0110011011: data <= 16'hff9e; 
        10'b0110011100: data <= 16'hff7c; 
        10'b0110011101: data <= 16'hffc0; 
        10'b0110011110: data <= 16'hffa5; 
        10'b0110011111: data <= 16'hffc3; 
        10'b0110100000: data <= 16'hffaf; 
        10'b0110100001: data <= 16'hffb7; 
        10'b0110100010: data <= 16'h0002; 
        10'b0110100011: data <= 16'h0004; 
        10'b0110100100: data <= 16'h0005; 
        10'b0110100101: data <= 16'hffd0; 
        10'b0110100110: data <= 16'h0007; 
        10'b0110100111: data <= 16'h0012; 
        10'b0110101000: data <= 16'hffeb; 
        10'b0110101001: data <= 16'hff8c; 
        10'b0110101010: data <= 16'hff29; 
        10'b0110101011: data <= 16'hff1a; 
        10'b0110101100: data <= 16'hff54; 
        10'b0110101101: data <= 16'hff9b; 
        10'b0110101110: data <= 16'hff90; 
        10'b0110101111: data <= 16'hffda; 
        10'b0110110000: data <= 16'h002e; 
        10'b0110110001: data <= 16'h00bf; 
        10'b0110110010: data <= 16'h006e; 
        10'b0110110011: data <= 16'hfff5; 
        10'b0110110100: data <= 16'hff60; 
        10'b0110110101: data <= 16'hffd2; 
        10'b0110110110: data <= 16'hfff0; 
        10'b0110110111: data <= 16'h002a; 
        10'b0110111000: data <= 16'h0063; 
        10'b0110111001: data <= 16'h0061; 
        10'b0110111010: data <= 16'h0021; 
        10'b0110111011: data <= 16'h000d; 
        10'b0110111100: data <= 16'hffc3; 
        10'b0110111101: data <= 16'hfff2; 
        10'b0110111110: data <= 16'hffed; 
        10'b0110111111: data <= 16'hffd0; 
        10'b0111000000: data <= 16'hffee; 
        10'b0111000001: data <= 16'hfff6; 
        10'b0111000010: data <= 16'h002c; 
        10'b0111000011: data <= 16'h0008; 
        10'b0111000100: data <= 16'h0020; 
        10'b0111000101: data <= 16'hffca; 
        10'b0111000110: data <= 16'hffa8; 
        10'b0111000111: data <= 16'hff68; 
        10'b0111001000: data <= 16'hfeb5; 
        10'b0111001001: data <= 16'hfea3; 
        10'b0111001010: data <= 16'hfecb; 
        10'b0111001011: data <= 16'hffb2; 
        10'b0111001100: data <= 16'h005c; 
        10'b0111001101: data <= 16'h00ef; 
        10'b0111001110: data <= 16'hffe6; 
        10'b0111001111: data <= 16'hff52; 
        10'b0111010000: data <= 16'hff48; 
        10'b0111010001: data <= 16'hffc4; 
        10'b0111010010: data <= 16'h004e; 
        10'b0111010011: data <= 16'h00cc; 
        10'b0111010100: data <= 16'h008f; 
        10'b0111010101: data <= 16'h00b4; 
        10'b0111010110: data <= 16'h00af; 
        10'b0111010111: data <= 16'h004e; 
        10'b0111011000: data <= 16'hffe9; 
        10'b0111011001: data <= 16'hfff1; 
        10'b0111011010: data <= 16'hfffe; 
        10'b0111011011: data <= 16'hfffa; 
        10'b0111011100: data <= 16'hfff9; 
        10'b0111011101: data <= 16'h0007; 
        10'b0111011110: data <= 16'h0001; 
        10'b0111011111: data <= 16'h0070; 
        10'b0111100000: data <= 16'h003e; 
        10'b0111100001: data <= 16'h0013; 
        10'b0111100010: data <= 16'hffc5; 
        10'b0111100011: data <= 16'hff37; 
        10'b0111100100: data <= 16'hfe9a; 
        10'b0111100101: data <= 16'hfdc9; 
        10'b0111100110: data <= 16'hfd3e; 
        10'b0111100111: data <= 16'hfd7c; 
        10'b0111101000: data <= 16'hfe17; 
        10'b0111101001: data <= 16'hfee9; 
        10'b0111101010: data <= 16'hfefd; 
        10'b0111101011: data <= 16'hff19; 
        10'b0111101100: data <= 16'hfff7; 
        10'b0111101101: data <= 16'h0047; 
        10'b0111101110: data <= 16'h0083; 
        10'b0111101111: data <= 16'h00cf; 
        10'b0111110000: data <= 16'h002b; 
        10'b0111110001: data <= 16'h00fa; 
        10'b0111110010: data <= 16'h00fa; 
        10'b0111110011: data <= 16'h004b; 
        10'b0111110100: data <= 16'hffdb; 
        10'b0111110101: data <= 16'hffcb; 
        10'b0111110110: data <= 16'hffd0; 
        10'b0111110111: data <= 16'hffd4; 
        10'b0111111000: data <= 16'hffe5; 
        10'b0111111001: data <= 16'hffe6; 
        10'b0111111010: data <= 16'h0016; 
        10'b0111111011: data <= 16'h00a5; 
        10'b0111111100: data <= 16'h0077; 
        10'b0111111101: data <= 16'h0048; 
        10'b0111111110: data <= 16'h0026; 
        10'b0111111111: data <= 16'hffd4; 
        10'b1000000000: data <= 16'hff81; 
        10'b1000000001: data <= 16'hfe61; 
        10'b1000000010: data <= 16'hfd9c; 
        10'b1000000011: data <= 16'hfdbd; 
        10'b1000000100: data <= 16'hfd45; 
        10'b1000000101: data <= 16'hfdc6; 
        10'b1000000110: data <= 16'hfe97; 
        10'b1000000111: data <= 16'hffae; 
        10'b1000001000: data <= 16'h0092; 
        10'b1000001001: data <= 16'h00c4; 
        10'b1000001010: data <= 16'h00d4; 
        10'b1000001011: data <= 16'h00d1; 
        10'b1000001100: data <= 16'h0092; 
        10'b1000001101: data <= 16'h0124; 
        10'b1000001110: data <= 16'h0110; 
        10'b1000001111: data <= 16'h0068; 
        10'b1000010000: data <= 16'hffa0; 
        10'b1000010001: data <= 16'hffbf; 
        10'b1000010010: data <= 16'hffd1; 
        10'b1000010011: data <= 16'hfff8; 
        10'b1000010100: data <= 16'hfff9; 
        10'b1000010101: data <= 16'hffd0; 
        10'b1000010110: data <= 16'hffe1; 
        10'b1000010111: data <= 16'h00cf; 
        10'b1000011000: data <= 16'h00d3; 
        10'b1000011001: data <= 16'h00f8; 
        10'b1000011010: data <= 16'h00d6; 
        10'b1000011011: data <= 16'h004e; 
        10'b1000011100: data <= 16'h0018; 
        10'b1000011101: data <= 16'hffa9; 
        10'b1000011110: data <= 16'hffc1; 
        10'b1000011111: data <= 16'hff3b; 
        10'b1000100000: data <= 16'hfee0; 
        10'b1000100001: data <= 16'hfece; 
        10'b1000100010: data <= 16'hff2f; 
        10'b1000100011: data <= 16'h004a; 
        10'b1000100100: data <= 16'h00c5; 
        10'b1000100101: data <= 16'h00f6; 
        10'b1000100110: data <= 16'h0114; 
        10'b1000100111: data <= 16'h00f7; 
        10'b1000101000: data <= 16'h00db; 
        10'b1000101001: data <= 16'h00ff; 
        10'b1000101010: data <= 16'h0062; 
        10'b1000101011: data <= 16'h000b; 
        10'b1000101100: data <= 16'hffaf; 
        10'b1000101101: data <= 16'hfff1; 
        10'b1000101110: data <= 16'hfff8; 
        10'b1000101111: data <= 16'hffef; 
        10'b1000110000: data <= 16'hfff6; 
        10'b1000110001: data <= 16'hffc1; 
        10'b1000110010: data <= 16'h0025; 
        10'b1000110011: data <= 16'h00de; 
        10'b1000110100: data <= 16'h0111; 
        10'b1000110101: data <= 16'h0128; 
        10'b1000110110: data <= 16'h0139; 
        10'b1000110111: data <= 16'h009e; 
        10'b1000111000: data <= 16'h00ba; 
        10'b1000111001: data <= 16'h00d2; 
        10'b1000111010: data <= 16'h004e; 
        10'b1000111011: data <= 16'hffeb; 
        10'b1000111100: data <= 16'hffb9; 
        10'b1000111101: data <= 16'hff94; 
        10'b1000111110: data <= 16'h0021; 
        10'b1000111111: data <= 16'h003a; 
        10'b1001000000: data <= 16'h006f; 
        10'b1001000001: data <= 16'h00c6; 
        10'b1001000010: data <= 16'h00cf; 
        10'b1001000011: data <= 16'h008d; 
        10'b1001000100: data <= 16'h00f6; 
        10'b1001000101: data <= 16'h008c; 
        10'b1001000110: data <= 16'hffe6; 
        10'b1001000111: data <= 16'hffc8; 
        10'b1001001000: data <= 16'hffbf; 
        10'b1001001001: data <= 16'hffed; 
        10'b1001001010: data <= 16'hffec; 
        10'b1001001011: data <= 16'hffea; 
        10'b1001001100: data <= 16'hffd6; 
        10'b1001001101: data <= 16'hfffd; 
        10'b1001001110: data <= 16'hfff1; 
        10'b1001001111: data <= 16'h006e; 
        10'b1001010000: data <= 16'h0108; 
        10'b1001010001: data <= 16'h0107; 
        10'b1001010010: data <= 16'h00e6; 
        10'b1001010011: data <= 16'h0082; 
        10'b1001010100: data <= 16'h008a; 
        10'b1001010101: data <= 16'h002e; 
        10'b1001010110: data <= 16'hffee; 
        10'b1001010111: data <= 16'hffc2; 
        10'b1001011000: data <= 16'h0014; 
        10'b1001011001: data <= 16'hfff5; 
        10'b1001011010: data <= 16'hfff0; 
        10'b1001011011: data <= 16'hffe2; 
        10'b1001011100: data <= 16'h0041; 
        10'b1001011101: data <= 16'h0018; 
        10'b1001011110: data <= 16'h007f; 
        10'b1001011111: data <= 16'h00cc; 
        10'b1001100000: data <= 16'h0076; 
        10'b1001100001: data <= 16'h002d; 
        10'b1001100010: data <= 16'hffd2; 
        10'b1001100011: data <= 16'hff8a; 
        10'b1001100100: data <= 16'hffda; 
        10'b1001100101: data <= 16'hffcf; 
        10'b1001100110: data <= 16'hffc0; 
        10'b1001100111: data <= 16'hffc4; 
        10'b1001101000: data <= 16'hffe5; 
        10'b1001101001: data <= 16'hffee; 
        10'b1001101010: data <= 16'hfff4; 
        10'b1001101011: data <= 16'h0045; 
        10'b1001101100: data <= 16'h0084; 
        10'b1001101101: data <= 16'h00b4; 
        10'b1001101110: data <= 16'h00a1; 
        10'b1001101111: data <= 16'h005c; 
        10'b1001110000: data <= 16'h0007; 
        10'b1001110001: data <= 16'h0042; 
        10'b1001110010: data <= 16'h0050; 
        10'b1001110011: data <= 16'h0061; 
        10'b1001110100: data <= 16'h001b; 
        10'b1001110101: data <= 16'hffdd; 
        10'b1001110110: data <= 16'hffda; 
        10'b1001110111: data <= 16'hffca; 
        10'b1001111000: data <= 16'h002a; 
        10'b1001111001: data <= 16'h0020; 
        10'b1001111010: data <= 16'h001f; 
        10'b1001111011: data <= 16'h008d; 
        10'b1001111100: data <= 16'h0044; 
        10'b1001111101: data <= 16'hffe8; 
        10'b1001111110: data <= 16'hffe0; 
        10'b1001111111: data <= 16'hffd7; 
        10'b1010000000: data <= 16'hffa6; 
        10'b1010000001: data <= 16'hffbc; 
        10'b1010000010: data <= 16'hfff4; 
        10'b1010000011: data <= 16'hfffe; 
        10'b1010000100: data <= 16'hffed; 
        10'b1010000101: data <= 16'hffcd; 
        10'b1010000110: data <= 16'hffd6; 
        10'b1010000111: data <= 16'h002d; 
        10'b1010001000: data <= 16'h0091; 
        10'b1010001001: data <= 16'h00da; 
        10'b1010001010: data <= 16'h00a3; 
        10'b1010001011: data <= 16'h00ac; 
        10'b1010001100: data <= 16'h002a; 
        10'b1010001101: data <= 16'h006e; 
        10'b1010001110: data <= 16'h0046; 
        10'b1010001111: data <= 16'hffff; 
        10'b1010010000: data <= 16'hffc9; 
        10'b1010010001: data <= 16'h0009; 
        10'b1010010010: data <= 16'h0016; 
        10'b1010010011: data <= 16'h0037; 
        10'b1010010100: data <= 16'h0029; 
        10'b1010010101: data <= 16'h0055; 
        10'b1010010110: data <= 16'h0087; 
        10'b1010010111: data <= 16'hffe9; 
        10'b1010011000: data <= 16'hffa5; 
        10'b1010011001: data <= 16'hffa6; 
        10'b1010011010: data <= 16'hffd1; 
        10'b1010011011: data <= 16'hffc5; 
        10'b1010011100: data <= 16'hfffb; 
        10'b1010011101: data <= 16'hfff1; 
        10'b1010011110: data <= 16'hffc8; 
        10'b1010011111: data <= 16'hffcd; 
        10'b1010100000: data <= 16'hffd8; 
        10'b1010100001: data <= 16'h0006; 
        10'b1010100010: data <= 16'h0007; 
        10'b1010100011: data <= 16'h0001; 
        10'b1010100100: data <= 16'h005d; 
        10'b1010100101: data <= 16'h0096; 
        10'b1010100110: data <= 16'h00b0; 
        10'b1010100111: data <= 16'h00d0; 
        10'b1010101000: data <= 16'h00d3; 
        10'b1010101001: data <= 16'h00ad; 
        10'b1010101010: data <= 16'h00fd; 
        10'b1010101011: data <= 16'h010b; 
        10'b1010101100: data <= 16'h0111; 
        10'b1010101101: data <= 16'h00d7; 
        10'b1010101110: data <= 16'h00be; 
        10'b1010101111: data <= 16'h008c; 
        10'b1010110000: data <= 16'h0086; 
        10'b1010110001: data <= 16'hfff4; 
        10'b1010110010: data <= 16'hff93; 
        10'b1010110011: data <= 16'hff69; 
        10'b1010110100: data <= 16'hff79; 
        10'b1010110101: data <= 16'hffad; 
        10'b1010110110: data <= 16'hffb3; 
        10'b1010110111: data <= 16'hffe9; 
        10'b1010111000: data <= 16'hffda; 
        10'b1010111001: data <= 16'hffff; 
        10'b1010111010: data <= 16'hffd9; 
        10'b1010111011: data <= 16'h0007; 
        10'b1010111100: data <= 16'hfffa; 
        10'b1010111101: data <= 16'hffbf; 
        10'b1010111110: data <= 16'h0005; 
        10'b1010111111: data <= 16'h000a; 
        10'b1011000000: data <= 16'hfff0; 
        10'b1011000001: data <= 16'h003a; 
        10'b1011000010: data <= 16'h0058; 
        10'b1011000011: data <= 16'h0031; 
        10'b1011000100: data <= 16'h0076; 
        10'b1011000101: data <= 16'h0078; 
        10'b1011000110: data <= 16'h00e0; 
        10'b1011000111: data <= 16'h0100; 
        10'b1011001000: data <= 16'h0113; 
        10'b1011001001: data <= 16'h00d7; 
        10'b1011001010: data <= 16'h0099; 
        10'b1011001011: data <= 16'h003d; 
        10'b1011001100: data <= 16'hffe7; 
        10'b1011001101: data <= 16'hff9f; 
        10'b1011001110: data <= 16'hff9f; 
        10'b1011001111: data <= 16'hffb0; 
        10'b1011010000: data <= 16'hffb1; 
        10'b1011010001: data <= 16'hffd8; 
        10'b1011010010: data <= 16'hffd8; 
        10'b1011010011: data <= 16'hfffc; 
        10'b1011010100: data <= 16'hffd0; 
        10'b1011010101: data <= 16'h0006; 
        10'b1011010110: data <= 16'hffc0; 
        10'b1011010111: data <= 16'hfff7; 
        10'b1011011000: data <= 16'hffd2; 
        10'b1011011001: data <= 16'hffbf; 
        10'b1011011010: data <= 16'hffc2; 
        10'b1011011011: data <= 16'hfff0; 
        10'b1011011100: data <= 16'hfff1; 
        10'b1011011101: data <= 16'hffd5; 
        10'b1011011110: data <= 16'hffce; 
        10'b1011011111: data <= 16'hffef; 
        10'b1011100000: data <= 16'hfff0; 
        10'b1011100001: data <= 16'hffeb; 
        10'b1011100010: data <= 16'hffe3; 
        10'b1011100011: data <= 16'hffe7; 
        10'b1011100100: data <= 16'hffdc; 
        10'b1011100101: data <= 16'hffec; 
        10'b1011100110: data <= 16'hffdb; 
        10'b1011100111: data <= 16'hffb9; 
        10'b1011101000: data <= 16'hffd5; 
        10'b1011101001: data <= 16'hffeb; 
        10'b1011101010: data <= 16'hffe4; 
        10'b1011101011: data <= 16'hffed; 
        10'b1011101100: data <= 16'hffc3; 
        10'b1011101101: data <= 16'hffc4; 
        10'b1011101110: data <= 16'hfff7; 
        10'b1011101111: data <= 16'hffdd; 
        10'b1011110000: data <= 16'h0002; 
        10'b1011110001: data <= 16'hffd1; 
        10'b1011110010: data <= 16'hfffb; 
        10'b1011110011: data <= 16'h0007; 
        10'b1011110100: data <= 16'hffe1; 
        10'b1011110101: data <= 16'hffcf; 
        10'b1011110110: data <= 16'hffea; 
        10'b1011110111: data <= 16'hffc3; 
        10'b1011111000: data <= 16'h0003; 
        10'b1011111001: data <= 16'hffef; 
        10'b1011111010: data <= 16'hfffd; 
        10'b1011111011: data <= 16'hffed; 
        10'b1011111100: data <= 16'hfff6; 
        10'b1011111101: data <= 16'hffc2; 
        10'b1011111110: data <= 16'hffcd; 
        10'b1011111111: data <= 16'hfff3; 
        10'b1100000000: data <= 16'hffcd; 
        10'b1100000001: data <= 16'hfff6; 
        10'b1100000010: data <= 16'hffda; 
        10'b1100000011: data <= 16'hffea; 
        10'b1100000100: data <= 16'hffdc; 
        10'b1100000101: data <= 16'hffff; 
        10'b1100000110: data <= 16'hffc5; 
        10'b1100000111: data <= 16'hffcf; 
        10'b1100001000: data <= 16'hfffc; 
        10'b1100001001: data <= 16'hffeb; 
        10'b1100001010: data <= 16'hffcf; 
        10'b1100001011: data <= 16'hfff1; 
        10'b1100001100: data <= 16'hffc6; 
        10'b1100001101: data <= 16'hffc1; 
        10'b1100001110: data <= 16'hfffc; 
        10'b1100001111: data <= 16'hffe3; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 11) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 17'h1ffd8; 
        10'b0000000001: data <= 17'h1ff9c; 
        10'b0000000010: data <= 17'h1fffb; 
        10'b0000000011: data <= 17'h00005; 
        10'b0000000100: data <= 17'h0000a; 
        10'b0000000101: data <= 17'h1fff7; 
        10'b0000000110: data <= 17'h1ffda; 
        10'b0000000111: data <= 17'h0000a; 
        10'b0000001000: data <= 17'h1ffb0; 
        10'b0000001001: data <= 17'h00006; 
        10'b0000001010: data <= 17'h00007; 
        10'b0000001011: data <= 17'h1ffbb; 
        10'b0000001100: data <= 17'h1ffba; 
        10'b0000001101: data <= 17'h1ffb8; 
        10'b0000001110: data <= 17'h1ffbd; 
        10'b0000001111: data <= 17'h1ffc6; 
        10'b0000010000: data <= 17'h00001; 
        10'b0000010001: data <= 17'h00004; 
        10'b0000010010: data <= 17'h1ff9d; 
        10'b0000010011: data <= 17'h0000a; 
        10'b0000010100: data <= 17'h1ffe0; 
        10'b0000010101: data <= 17'h1ffe4; 
        10'b0000010110: data <= 17'h1ff7d; 
        10'b0000010111: data <= 17'h1fff9; 
        10'b0000011000: data <= 17'h1fffb; 
        10'b0000011001: data <= 17'h1ff85; 
        10'b0000011010: data <= 17'h1ffc4; 
        10'b0000011011: data <= 17'h00004; 
        10'b0000011100: data <= 17'h1ff99; 
        10'b0000011101: data <= 17'h1ffc0; 
        10'b0000011110: data <= 17'h1ff9b; 
        10'b0000011111: data <= 17'h1ffdd; 
        10'b0000100000: data <= 17'h1ff8c; 
        10'b0000100001: data <= 17'h1ffc9; 
        10'b0000100010: data <= 17'h0000d; 
        10'b0000100011: data <= 17'h00007; 
        10'b0000100100: data <= 17'h1ff84; 
        10'b0000100101: data <= 17'h1ff7f; 
        10'b0000100110: data <= 17'h1ff8c; 
        10'b0000100111: data <= 17'h1ffda; 
        10'b0000101000: data <= 17'h1ffe4; 
        10'b0000101001: data <= 17'h1ffc5; 
        10'b0000101010: data <= 17'h1ffbb; 
        10'b0000101011: data <= 17'h1ffa3; 
        10'b0000101100: data <= 17'h0000d; 
        10'b0000101101: data <= 17'h1ff9d; 
        10'b0000101110: data <= 17'h1ffea; 
        10'b0000101111: data <= 17'h1ffb4; 
        10'b0000110000: data <= 17'h1ffb6; 
        10'b0000110001: data <= 17'h1ff88; 
        10'b0000110010: data <= 17'h1ffce; 
        10'b0000110011: data <= 17'h1fff4; 
        10'b0000110100: data <= 17'h1ff94; 
        10'b0000110101: data <= 17'h1fffa; 
        10'b0000110110: data <= 17'h1ffd5; 
        10'b0000110111: data <= 17'h1ff95; 
        10'b0000111000: data <= 17'h1ffa6; 
        10'b0000111001: data <= 17'h1ffcd; 
        10'b0000111010: data <= 17'h1ffca; 
        10'b0000111011: data <= 17'h1ff9d; 
        10'b0000111100: data <= 17'h1ffe0; 
        10'b0000111101: data <= 17'h1ffeb; 
        10'b0000111110: data <= 17'h1ffab; 
        10'b0000111111: data <= 17'h1ffe9; 
        10'b0001000000: data <= 17'h1fff5; 
        10'b0001000001: data <= 17'h1ffc5; 
        10'b0001000010: data <= 17'h1ff92; 
        10'b0001000011: data <= 17'h1ff95; 
        10'b0001000100: data <= 17'h1ff87; 
        10'b0001000101: data <= 17'h1ff97; 
        10'b0001000110: data <= 17'h1ffbe; 
        10'b0001000111: data <= 17'h1ffb4; 
        10'b0001001000: data <= 17'h1ffaa; 
        10'b0001001001: data <= 17'h1ffa7; 
        10'b0001001010: data <= 17'h1ffe9; 
        10'b0001001011: data <= 17'h1fffd; 
        10'b0001001100: data <= 17'h1ffc2; 
        10'b0001001101: data <= 17'h1ff9a; 
        10'b0001001110: data <= 17'h0000b; 
        10'b0001001111: data <= 17'h1fff8; 
        10'b0001010000: data <= 17'h00000; 
        10'b0001010001: data <= 17'h1ffb1; 
        10'b0001010010: data <= 17'h1ff83; 
        10'b0001010011: data <= 17'h1ffc6; 
        10'b0001010100: data <= 17'h0000e; 
        10'b0001010101: data <= 17'h1ffe8; 
        10'b0001010110: data <= 17'h1ffc7; 
        10'b0001010111: data <= 17'h1fff1; 
        10'b0001011000: data <= 17'h1ffe7; 
        10'b0001011001: data <= 17'h00001; 
        10'b0001011010: data <= 17'h1ffda; 
        10'b0001011011: data <= 17'h1fff9; 
        10'b0001011100: data <= 17'h1fff1; 
        10'b0001011101: data <= 17'h1ffd0; 
        10'b0001011110: data <= 17'h0002c; 
        10'b0001011111: data <= 17'h00094; 
        10'b0001100000: data <= 17'h00139; 
        10'b0001100001: data <= 17'h00104; 
        10'b0001100010: data <= 17'h00109; 
        10'b0001100011: data <= 17'h00124; 
        10'b0001100100: data <= 17'h000cb; 
        10'b0001100101: data <= 17'h000e5; 
        10'b0001100110: data <= 17'h000b3; 
        10'b0001100111: data <= 17'h0000d; 
        10'b0001101000: data <= 17'h1ffee; 
        10'b0001101001: data <= 17'h1ff26; 
        10'b0001101010: data <= 17'h1ff82; 
        10'b0001101011: data <= 17'h1fff5; 
        10'b0001101100: data <= 17'h00006; 
        10'b0001101101: data <= 17'h1ffa0; 
        10'b0001101110: data <= 17'h1ffd4; 
        10'b0001101111: data <= 17'h1ffac; 
        10'b0001110000: data <= 17'h1ffd3; 
        10'b0001110001: data <= 17'h1fff9; 
        10'b0001110010: data <= 17'h1ffde; 
        10'b0001110011: data <= 17'h00004; 
        10'b0001110100: data <= 17'h00030; 
        10'b0001110101: data <= 17'h00000; 
        10'b0001110110: data <= 17'h000b8; 
        10'b0001110111: data <= 17'h0009b; 
        10'b0001111000: data <= 17'h001a7; 
        10'b0001111001: data <= 17'h0016b; 
        10'b0001111010: data <= 17'h001c3; 
        10'b0001111011: data <= 17'h0021e; 
        10'b0001111100: data <= 17'h00275; 
        10'b0001111101: data <= 17'h002a2; 
        10'b0001111110: data <= 17'h0025e; 
        10'b0001111111: data <= 17'h001bc; 
        10'b0010000000: data <= 17'h000fb; 
        10'b0010000001: data <= 17'h000c8; 
        10'b0010000010: data <= 17'h00148; 
        10'b0010000011: data <= 17'h00028; 
        10'b0010000100: data <= 17'h1ff20; 
        10'b0010000101: data <= 17'h1fea2; 
        10'b0010000110: data <= 17'h1fed5; 
        10'b0010000111: data <= 17'h1fedb; 
        10'b0010001000: data <= 17'h1ffdc; 
        10'b0010001001: data <= 17'h1ffcb; 
        10'b0010001010: data <= 17'h1ffb4; 
        10'b0010001011: data <= 17'h1ffec; 
        10'b0010001100: data <= 17'h1ff92; 
        10'b0010001101: data <= 17'h1ff82; 
        10'b0010001110: data <= 17'h1ffa2; 
        10'b0010001111: data <= 17'h1ffa2; 
        10'b0010010000: data <= 17'h00018; 
        10'b0010010001: data <= 17'h000bf; 
        10'b0010010010: data <= 17'h0015d; 
        10'b0010010011: data <= 17'h00117; 
        10'b0010010100: data <= 17'h00140; 
        10'b0010010101: data <= 17'h0011a; 
        10'b0010010110: data <= 17'h000ff; 
        10'b0010010111: data <= 17'h0014c; 
        10'b0010011000: data <= 17'h00151; 
        10'b0010011001: data <= 17'h00195; 
        10'b0010011010: data <= 17'h00045; 
        10'b0010011011: data <= 17'h0010e; 
        10'b0010011100: data <= 17'h00137; 
        10'b0010011101: data <= 17'h1ffe8; 
        10'b0010011110: data <= 17'h1ffef; 
        10'b0010011111: data <= 17'h1ff73; 
        10'b0010100000: data <= 17'h1ff3c; 
        10'b0010100001: data <= 17'h1fe60; 
        10'b0010100010: data <= 17'h1fdeb; 
        10'b0010100011: data <= 17'h1fe3d; 
        10'b0010100100: data <= 17'h1ff7d; 
        10'b0010100101: data <= 17'h00001; 
        10'b0010100110: data <= 17'h1ffa6; 
        10'b0010100111: data <= 17'h1ffc9; 
        10'b0010101000: data <= 17'h1ff9d; 
        10'b0010101001: data <= 17'h1ffb2; 
        10'b0010101010: data <= 17'h1ffaa; 
        10'b0010101011: data <= 17'h00028; 
        10'b0010101100: data <= 17'h000ed; 
        10'b0010101101: data <= 17'h001b8; 
        10'b0010101110: data <= 17'h00150; 
        10'b0010101111: data <= 17'h00102; 
        10'b0010110000: data <= 17'h00186; 
        10'b0010110001: data <= 17'h0013f; 
        10'b0010110010: data <= 17'h0011b; 
        10'b0010110011: data <= 17'h0010f; 
        10'b0010110100: data <= 17'h0016a; 
        10'b0010110101: data <= 17'h00208; 
        10'b0010110110: data <= 17'h00169; 
        10'b0010110111: data <= 17'h00082; 
        10'b0010111000: data <= 17'h00158; 
        10'b0010111001: data <= 17'h0013b; 
        10'b0010111010: data <= 17'h0012c; 
        10'b0010111011: data <= 17'h1ff7a; 
        10'b0010111100: data <= 17'h00080; 
        10'b0010111101: data <= 17'h1ff81; 
        10'b0010111110: data <= 17'h1fe37; 
        10'b0010111111: data <= 17'h1fe37; 
        10'b0011000000: data <= 17'h1fee8; 
        10'b0011000001: data <= 17'h1ffc8; 
        10'b0011000010: data <= 17'h1fff4; 
        10'b0011000011: data <= 17'h1ffd4; 
        10'b0011000100: data <= 17'h00005; 
        10'b0011000101: data <= 17'h1fff1; 
        10'b0011000110: data <= 17'h0001b; 
        10'b0011000111: data <= 17'h000c6; 
        10'b0011001000: data <= 17'h00207; 
        10'b0011001001: data <= 17'h00205; 
        10'b0011001010: data <= 17'h0016c; 
        10'b0011001011: data <= 17'h00066; 
        10'b0011001100: data <= 17'h0006e; 
        10'b0011001101: data <= 17'h000e7; 
        10'b0011001110: data <= 17'h00047; 
        10'b0011001111: data <= 17'h0006a; 
        10'b0011010000: data <= 17'h00131; 
        10'b0011010001: data <= 17'h00121; 
        10'b0011010010: data <= 17'h001de; 
        10'b0011010011: data <= 17'h00119; 
        10'b0011010100: data <= 17'h00056; 
        10'b0011010101: data <= 17'h000f0; 
        10'b0011010110: data <= 17'h000c7; 
        10'b0011010111: data <= 17'h000d8; 
        10'b0011011000: data <= 17'h000db; 
        10'b0011011001: data <= 17'h0001f; 
        10'b0011011010: data <= 17'h1ff23; 
        10'b0011011011: data <= 17'h1fdff; 
        10'b0011011100: data <= 17'h1fe90; 
        10'b0011011101: data <= 17'h1ff9f; 
        10'b0011011110: data <= 17'h1ff82; 
        10'b0011011111: data <= 17'h1ffbd; 
        10'b0011100000: data <= 17'h1ffcf; 
        10'b0011100001: data <= 17'h1ffb5; 
        10'b0011100010: data <= 17'h00016; 
        10'b0011100011: data <= 17'h000b8; 
        10'b0011100100: data <= 17'h001ac; 
        10'b0011100101: data <= 17'h00197; 
        10'b0011100110: data <= 17'h00132; 
        10'b0011100111: data <= 17'h0007d; 
        10'b0011101000: data <= 17'h000cf; 
        10'b0011101001: data <= 17'h00063; 
        10'b0011101010: data <= 17'h00106; 
        10'b0011101011: data <= 17'h00054; 
        10'b0011101100: data <= 17'h00047; 
        10'b0011101101: data <= 17'h00080; 
        10'b0011101110: data <= 17'h00208; 
        10'b0011101111: data <= 17'h001af; 
        10'b0011110000: data <= 17'h00064; 
        10'b0011110001: data <= 17'h000f0; 
        10'b0011110010: data <= 17'h00159; 
        10'b0011110011: data <= 17'h000e1; 
        10'b0011110100: data <= 17'h00149; 
        10'b0011110101: data <= 17'h000a9; 
        10'b0011110110: data <= 17'h1ffa8; 
        10'b0011110111: data <= 17'h1fe25; 
        10'b0011111000: data <= 17'h1fe9c; 
        10'b0011111001: data <= 17'h1ff7e; 
        10'b0011111010: data <= 17'h1ff92; 
        10'b0011111011: data <= 17'h1ffb1; 
        10'b0011111100: data <= 17'h1ffc2; 
        10'b0011111101: data <= 17'h1ff86; 
        10'b0011111110: data <= 17'h1ffd9; 
        10'b0011111111: data <= 17'h00050; 
        10'b0100000000: data <= 17'h000dd; 
        10'b0100000001: data <= 17'h00126; 
        10'b0100000010: data <= 17'h000f3; 
        10'b0100000011: data <= 17'h0003b; 
        10'b0100000100: data <= 17'h1ffe1; 
        10'b0100000101: data <= 17'h1ff1d; 
        10'b0100000110: data <= 17'h1fe50; 
        10'b0100000111: data <= 17'h1fce6; 
        10'b0100001000: data <= 17'h1fd7c; 
        10'b0100001001: data <= 17'h1ffaa; 
        10'b0100001010: data <= 17'h0026b; 
        10'b0100001011: data <= 17'h003b8; 
        10'b0100001100: data <= 17'h00226; 
        10'b0100001101: data <= 17'h00142; 
        10'b0100001110: data <= 17'h0015e; 
        10'b0100001111: data <= 17'h00143; 
        10'b0100010000: data <= 17'h001e4; 
        10'b0100010001: data <= 17'h00135; 
        10'b0100010010: data <= 17'h1ffa2; 
        10'b0100010011: data <= 17'h1fe28; 
        10'b0100010100: data <= 17'h1ff12; 
        10'b0100010101: data <= 17'h1ff7a; 
        10'b0100010110: data <= 17'h1ff9b; 
        10'b0100010111: data <= 17'h1ffac; 
        10'b0100011000: data <= 17'h1fff3; 
        10'b0100011001: data <= 17'h1ffec; 
        10'b0100011010: data <= 17'h00007; 
        10'b0100011011: data <= 17'h00077; 
        10'b0100011100: data <= 17'h0006b; 
        10'b0100011101: data <= 17'h0002e; 
        10'b0100011110: data <= 17'h1ff76; 
        10'b0100011111: data <= 17'h1fea1; 
        10'b0100100000: data <= 17'h1fd7f; 
        10'b0100100001: data <= 17'h1fc6b; 
        10'b0100100010: data <= 17'h1fb9d; 
        10'b0100100011: data <= 17'h1fb80; 
        10'b0100100100: data <= 17'h1fcaf; 
        10'b0100100101: data <= 17'h1ff2a; 
        10'b0100100110: data <= 17'h001fc; 
        10'b0100100111: data <= 17'h0024b; 
        10'b0100101000: data <= 17'h001f4; 
        10'b0100101001: data <= 17'h001d2; 
        10'b0100101010: data <= 17'h00120; 
        10'b0100101011: data <= 17'h001f3; 
        10'b0100101100: data <= 17'h001cf; 
        10'b0100101101: data <= 17'h000ba; 
        10'b0100101110: data <= 17'h1ff5a; 
        10'b0100101111: data <= 17'h1fece; 
        10'b0100110000: data <= 17'h1ff8e; 
        10'b0100110001: data <= 17'h1ff7e; 
        10'b0100110010: data <= 17'h1ffc9; 
        10'b0100110011: data <= 17'h1fff2; 
        10'b0100110100: data <= 17'h0000f; 
        10'b0100110101: data <= 17'h1fff2; 
        10'b0100110110: data <= 17'h1ff96; 
        10'b0100110111: data <= 17'h00074; 
        10'b0100111000: data <= 17'h1ffbb; 
        10'b0100111001: data <= 17'h1fe99; 
        10'b0100111010: data <= 17'h1fde5; 
        10'b0100111011: data <= 17'h1fce7; 
        10'b0100111100: data <= 17'h1fc21; 
        10'b0100111101: data <= 17'h1fca8; 
        10'b0100111110: data <= 17'h1fd74; 
        10'b0100111111: data <= 17'h1fecd; 
        10'b0101000000: data <= 17'h1ff5a; 
        10'b0101000001: data <= 17'h000d7; 
        10'b0101000010: data <= 17'h00152; 
        10'b0101000011: data <= 17'h00154; 
        10'b0101000100: data <= 17'h0009b; 
        10'b0101000101: data <= 17'h00160; 
        10'b0101000110: data <= 17'h001b3; 
        10'b0101000111: data <= 17'h001a9; 
        10'b0101001000: data <= 17'h00173; 
        10'b0101001001: data <= 17'h00002; 
        10'b0101001010: data <= 17'h1ff5d; 
        10'b0101001011: data <= 17'h1ff77; 
        10'b0101001100: data <= 17'h1ff88; 
        10'b0101001101: data <= 17'h1ffb9; 
        10'b0101001110: data <= 17'h1ff9d; 
        10'b0101001111: data <= 17'h1ff92; 
        10'b0101010000: data <= 17'h00004; 
        10'b0101010001: data <= 17'h1ffad; 
        10'b0101010010: data <= 17'h1ffeb; 
        10'b0101010011: data <= 17'h1fffa; 
        10'b0101010100: data <= 17'h1ff7d; 
        10'b0101010101: data <= 17'h1fe97; 
        10'b0101010110: data <= 17'h1fd88; 
        10'b0101010111: data <= 17'h1fcea; 
        10'b0101011000: data <= 17'h1fd35; 
        10'b0101011001: data <= 17'h1fe83; 
        10'b0101011010: data <= 17'h00007; 
        10'b0101011011: data <= 17'h0003f; 
        10'b0101011100: data <= 17'h00065; 
        10'b0101011101: data <= 17'h000e4; 
        10'b0101011110: data <= 17'h00236; 
        10'b0101011111: data <= 17'h00124; 
        10'b0101100000: data <= 17'h000c8; 
        10'b0101100001: data <= 17'h0011a; 
        10'b0101100010: data <= 17'h000e2; 
        10'b0101100011: data <= 17'h1ffec; 
        10'b0101100100: data <= 17'h1fedb; 
        10'b0101100101: data <= 17'h1fe6e; 
        10'b0101100110: data <= 17'h1fe5b; 
        10'b0101100111: data <= 17'h1fef4; 
        10'b0101101000: data <= 17'h1ffd1; 
        10'b0101101001: data <= 17'h1ffaf; 
        10'b0101101010: data <= 17'h1ffd4; 
        10'b0101101011: data <= 17'h1ffe1; 
        10'b0101101100: data <= 17'h1ffc7; 
        10'b0101101101: data <= 17'h1ffa9; 
        10'b0101101110: data <= 17'h1ffcb; 
        10'b0101101111: data <= 17'h1ffdc; 
        10'b0101110000: data <= 17'h1ff59; 
        10'b0101110001: data <= 17'h1ff09; 
        10'b0101110010: data <= 17'h1fdfe; 
        10'b0101110011: data <= 17'h1fdaf; 
        10'b0101110100: data <= 17'h1fe6e; 
        10'b0101110101: data <= 17'h1ffb1; 
        10'b0101110110: data <= 17'h1ff7d; 
        10'b0101110111: data <= 17'h1feab; 
        10'b0101111000: data <= 17'h0001b; 
        10'b0101111001: data <= 17'h001e7; 
        10'b0101111010: data <= 17'h001ec; 
        10'b0101111011: data <= 17'h0005a; 
        10'b0101111100: data <= 17'h000df; 
        10'b0101111101: data <= 17'h000ee; 
        10'b0101111110: data <= 17'h0007e; 
        10'b0101111111: data <= 17'h1ff58; 
        10'b0110000000: data <= 17'h1fe3f; 
        10'b0110000001: data <= 17'h1fe3d; 
        10'b0110000010: data <= 17'h1fe9c; 
        10'b0110000011: data <= 17'h1ff06; 
        10'b0110000100: data <= 17'h1ff70; 
        10'b0110000101: data <= 17'h1fffd; 
        10'b0110000110: data <= 17'h1ffe6; 
        10'b0110000111: data <= 17'h1ffb4; 
        10'b0110001000: data <= 17'h0000c; 
        10'b0110001001: data <= 17'h1ff9e; 
        10'b0110001010: data <= 17'h1ffc1; 
        10'b0110001011: data <= 17'h1ffd7; 
        10'b0110001100: data <= 17'h1ffe1; 
        10'b0110001101: data <= 17'h1ff32; 
        10'b0110001110: data <= 17'h1fe30; 
        10'b0110001111: data <= 17'h1fe5d; 
        10'b0110010000: data <= 17'h1fee3; 
        10'b0110010001: data <= 17'h1ffd8; 
        10'b0110010010: data <= 17'h1fed6; 
        10'b0110010011: data <= 17'h1fec2; 
        10'b0110010100: data <= 17'h0005a; 
        10'b0110010101: data <= 17'h000ec; 
        10'b0110010110: data <= 17'h000fc; 
        10'b0110010111: data <= 17'h1ffdb; 
        10'b0110011000: data <= 17'h1ff9a; 
        10'b0110011001: data <= 17'h1ffb4; 
        10'b0110011010: data <= 17'h00022; 
        10'b0110011011: data <= 17'h1ff3d; 
        10'b0110011100: data <= 17'h1fef8; 
        10'b0110011101: data <= 17'h1ff80; 
        10'b0110011110: data <= 17'h1ff4a; 
        10'b0110011111: data <= 17'h1ff85; 
        10'b0110100000: data <= 17'h1ff5e; 
        10'b0110100001: data <= 17'h1ff6f; 
        10'b0110100010: data <= 17'h00004; 
        10'b0110100011: data <= 17'h00007; 
        10'b0110100100: data <= 17'h0000b; 
        10'b0110100101: data <= 17'h1ffa0; 
        10'b0110100110: data <= 17'h0000e; 
        10'b0110100111: data <= 17'h00024; 
        10'b0110101000: data <= 17'h1ffd7; 
        10'b0110101001: data <= 17'h1ff18; 
        10'b0110101010: data <= 17'h1fe52; 
        10'b0110101011: data <= 17'h1fe34; 
        10'b0110101100: data <= 17'h1fea8; 
        10'b0110101101: data <= 17'h1ff36; 
        10'b0110101110: data <= 17'h1ff20; 
        10'b0110101111: data <= 17'h1ffb4; 
        10'b0110110000: data <= 17'h0005d; 
        10'b0110110001: data <= 17'h0017f; 
        10'b0110110010: data <= 17'h000dc; 
        10'b0110110011: data <= 17'h1ffea; 
        10'b0110110100: data <= 17'h1fec0; 
        10'b0110110101: data <= 17'h1ffa3; 
        10'b0110110110: data <= 17'h1ffe1; 
        10'b0110110111: data <= 17'h00054; 
        10'b0110111000: data <= 17'h000c6; 
        10'b0110111001: data <= 17'h000c2; 
        10'b0110111010: data <= 17'h00043; 
        10'b0110111011: data <= 17'h00019; 
        10'b0110111100: data <= 17'h1ff87; 
        10'b0110111101: data <= 17'h1ffe5; 
        10'b0110111110: data <= 17'h1ffda; 
        10'b0110111111: data <= 17'h1ff9f; 
        10'b0111000000: data <= 17'h1ffdc; 
        10'b0111000001: data <= 17'h1ffeb; 
        10'b0111000010: data <= 17'h00058; 
        10'b0111000011: data <= 17'h00010; 
        10'b0111000100: data <= 17'h00041; 
        10'b0111000101: data <= 17'h1ff95; 
        10'b0111000110: data <= 17'h1ff50; 
        10'b0111000111: data <= 17'h1fed0; 
        10'b0111001000: data <= 17'h1fd6a; 
        10'b0111001001: data <= 17'h1fd46; 
        10'b0111001010: data <= 17'h1fd96; 
        10'b0111001011: data <= 17'h1ff63; 
        10'b0111001100: data <= 17'h000b8; 
        10'b0111001101: data <= 17'h001de; 
        10'b0111001110: data <= 17'h1ffcc; 
        10'b0111001111: data <= 17'h1fea3; 
        10'b0111010000: data <= 17'h1fe8f; 
        10'b0111010001: data <= 17'h1ff88; 
        10'b0111010010: data <= 17'h0009b; 
        10'b0111010011: data <= 17'h00197; 
        10'b0111010100: data <= 17'h0011f; 
        10'b0111010101: data <= 17'h00169; 
        10'b0111010110: data <= 17'h0015e; 
        10'b0111010111: data <= 17'h0009b; 
        10'b0111011000: data <= 17'h1ffd2; 
        10'b0111011001: data <= 17'h1ffe1; 
        10'b0111011010: data <= 17'h1fffc; 
        10'b0111011011: data <= 17'h1fff4; 
        10'b0111011100: data <= 17'h1fff2; 
        10'b0111011101: data <= 17'h0000f; 
        10'b0111011110: data <= 17'h00002; 
        10'b0111011111: data <= 17'h000df; 
        10'b0111100000: data <= 17'h0007b; 
        10'b0111100001: data <= 17'h00027; 
        10'b0111100010: data <= 17'h1ff8a; 
        10'b0111100011: data <= 17'h1fe6e; 
        10'b0111100100: data <= 17'h1fd35; 
        10'b0111100101: data <= 17'h1fb92; 
        10'b0111100110: data <= 17'h1fa7c; 
        10'b0111100111: data <= 17'h1faf8; 
        10'b0111101000: data <= 17'h1fc2e; 
        10'b0111101001: data <= 17'h1fdd3; 
        10'b0111101010: data <= 17'h1fdfb; 
        10'b0111101011: data <= 17'h1fe32; 
        10'b0111101100: data <= 17'h1ffee; 
        10'b0111101101: data <= 17'h0008e; 
        10'b0111101110: data <= 17'h00105; 
        10'b0111101111: data <= 17'h0019d; 
        10'b0111110000: data <= 17'h00056; 
        10'b0111110001: data <= 17'h001f4; 
        10'b0111110010: data <= 17'h001f3; 
        10'b0111110011: data <= 17'h00096; 
        10'b0111110100: data <= 17'h1ffb6; 
        10'b0111110101: data <= 17'h1ff96; 
        10'b0111110110: data <= 17'h1ff9f; 
        10'b0111110111: data <= 17'h1ffa7; 
        10'b0111111000: data <= 17'h1ffc9; 
        10'b0111111001: data <= 17'h1ffcd; 
        10'b0111111010: data <= 17'h0002b; 
        10'b0111111011: data <= 17'h0014a; 
        10'b0111111100: data <= 17'h000ee; 
        10'b0111111101: data <= 17'h0008f; 
        10'b0111111110: data <= 17'h0004b; 
        10'b0111111111: data <= 17'h1ffa9; 
        10'b1000000000: data <= 17'h1ff02; 
        10'b1000000001: data <= 17'h1fcc2; 
        10'b1000000010: data <= 17'h1fb39; 
        10'b1000000011: data <= 17'h1fb7b; 
        10'b1000000100: data <= 17'h1fa8b; 
        10'b1000000101: data <= 17'h1fb8c; 
        10'b1000000110: data <= 17'h1fd2f; 
        10'b1000000111: data <= 17'h1ff5c; 
        10'b1000001000: data <= 17'h00123; 
        10'b1000001001: data <= 17'h00189; 
        10'b1000001010: data <= 17'h001a7; 
        10'b1000001011: data <= 17'h001a2; 
        10'b1000001100: data <= 17'h00125; 
        10'b1000001101: data <= 17'h00248; 
        10'b1000001110: data <= 17'h00221; 
        10'b1000001111: data <= 17'h000d0; 
        10'b1000010000: data <= 17'h1ff40; 
        10'b1000010001: data <= 17'h1ff7e; 
        10'b1000010010: data <= 17'h1ffa2; 
        10'b1000010011: data <= 17'h1fff1; 
        10'b1000010100: data <= 17'h1fff1; 
        10'b1000010101: data <= 17'h1ffa1; 
        10'b1000010110: data <= 17'h1ffc3; 
        10'b1000010111: data <= 17'h0019e; 
        10'b1000011000: data <= 17'h001a6; 
        10'b1000011001: data <= 17'h001f0; 
        10'b1000011010: data <= 17'h001ab; 
        10'b1000011011: data <= 17'h0009d; 
        10'b1000011100: data <= 17'h0002f; 
        10'b1000011101: data <= 17'h1ff52; 
        10'b1000011110: data <= 17'h1ff82; 
        10'b1000011111: data <= 17'h1fe76; 
        10'b1000100000: data <= 17'h1fdc0; 
        10'b1000100001: data <= 17'h1fd9b; 
        10'b1000100010: data <= 17'h1fe5f; 
        10'b1000100011: data <= 17'h00093; 
        10'b1000100100: data <= 17'h0018a; 
        10'b1000100101: data <= 17'h001ed; 
        10'b1000100110: data <= 17'h00228; 
        10'b1000100111: data <= 17'h001ee; 
        10'b1000101000: data <= 17'h001b5; 
        10'b1000101001: data <= 17'h001fe; 
        10'b1000101010: data <= 17'h000c3; 
        10'b1000101011: data <= 17'h00017; 
        10'b1000101100: data <= 17'h1ff5e; 
        10'b1000101101: data <= 17'h1ffe2; 
        10'b1000101110: data <= 17'h1fff0; 
        10'b1000101111: data <= 17'h1ffdd; 
        10'b1000110000: data <= 17'h1ffeb; 
        10'b1000110001: data <= 17'h1ff82; 
        10'b1000110010: data <= 17'h0004b; 
        10'b1000110011: data <= 17'h001bc; 
        10'b1000110100: data <= 17'h00222; 
        10'b1000110101: data <= 17'h0024f; 
        10'b1000110110: data <= 17'h00272; 
        10'b1000110111: data <= 17'h0013c; 
        10'b1000111000: data <= 17'h00174; 
        10'b1000111001: data <= 17'h001a5; 
        10'b1000111010: data <= 17'h0009b; 
        10'b1000111011: data <= 17'h1ffd6; 
        10'b1000111100: data <= 17'h1ff73; 
        10'b1000111101: data <= 17'h1ff28; 
        10'b1000111110: data <= 17'h00041; 
        10'b1000111111: data <= 17'h00074; 
        10'b1001000000: data <= 17'h000de; 
        10'b1001000001: data <= 17'h0018c; 
        10'b1001000010: data <= 17'h0019f; 
        10'b1001000011: data <= 17'h0011a; 
        10'b1001000100: data <= 17'h001ec; 
        10'b1001000101: data <= 17'h00117; 
        10'b1001000110: data <= 17'h1ffcc; 
        10'b1001000111: data <= 17'h1ff90; 
        10'b1001001000: data <= 17'h1ff7e; 
        10'b1001001001: data <= 17'h1ffda; 
        10'b1001001010: data <= 17'h1ffd8; 
        10'b1001001011: data <= 17'h1ffd3; 
        10'b1001001100: data <= 17'h1ffab; 
        10'b1001001101: data <= 17'h1fffa; 
        10'b1001001110: data <= 17'h1ffe1; 
        10'b1001001111: data <= 17'h000dd; 
        10'b1001010000: data <= 17'h0020f; 
        10'b1001010001: data <= 17'h0020f; 
        10'b1001010010: data <= 17'h001cc; 
        10'b1001010011: data <= 17'h00103; 
        10'b1001010100: data <= 17'h00115; 
        10'b1001010101: data <= 17'h0005c; 
        10'b1001010110: data <= 17'h1ffdc; 
        10'b1001010111: data <= 17'h1ff84; 
        10'b1001011000: data <= 17'h00028; 
        10'b1001011001: data <= 17'h1ffea; 
        10'b1001011010: data <= 17'h1ffdf; 
        10'b1001011011: data <= 17'h1ffc3; 
        10'b1001011100: data <= 17'h00081; 
        10'b1001011101: data <= 17'h0002f; 
        10'b1001011110: data <= 17'h000fd; 
        10'b1001011111: data <= 17'h00197; 
        10'b1001100000: data <= 17'h000ed; 
        10'b1001100001: data <= 17'h0005b; 
        10'b1001100010: data <= 17'h1ffa4; 
        10'b1001100011: data <= 17'h1ff13; 
        10'b1001100100: data <= 17'h1ffb3; 
        10'b1001100101: data <= 17'h1ff9e; 
        10'b1001100110: data <= 17'h1ff7f; 
        10'b1001100111: data <= 17'h1ff88; 
        10'b1001101000: data <= 17'h1ffcb; 
        10'b1001101001: data <= 17'h1ffdb; 
        10'b1001101010: data <= 17'h1ffe7; 
        10'b1001101011: data <= 17'h00089; 
        10'b1001101100: data <= 17'h00109; 
        10'b1001101101: data <= 17'h00168; 
        10'b1001101110: data <= 17'h00142; 
        10'b1001101111: data <= 17'h000b7; 
        10'b1001110000: data <= 17'h0000e; 
        10'b1001110001: data <= 17'h00084; 
        10'b1001110010: data <= 17'h000a0; 
        10'b1001110011: data <= 17'h000c2; 
        10'b1001110100: data <= 17'h00036; 
        10'b1001110101: data <= 17'h1ffb9; 
        10'b1001110110: data <= 17'h1ffb5; 
        10'b1001110111: data <= 17'h1ff95; 
        10'b1001111000: data <= 17'h00054; 
        10'b1001111001: data <= 17'h00040; 
        10'b1001111010: data <= 17'h0003f; 
        10'b1001111011: data <= 17'h00119; 
        10'b1001111100: data <= 17'h00089; 
        10'b1001111101: data <= 17'h1ffd0; 
        10'b1001111110: data <= 17'h1ffc1; 
        10'b1001111111: data <= 17'h1ffae; 
        10'b1010000000: data <= 17'h1ff4b; 
        10'b1010000001: data <= 17'h1ff78; 
        10'b1010000010: data <= 17'h1ffe7; 
        10'b1010000011: data <= 17'h1fffc; 
        10'b1010000100: data <= 17'h1ffda; 
        10'b1010000101: data <= 17'h1ff9a; 
        10'b1010000110: data <= 17'h1ffac; 
        10'b1010000111: data <= 17'h0005a; 
        10'b1010001000: data <= 17'h00121; 
        10'b1010001001: data <= 17'h001b5; 
        10'b1010001010: data <= 17'h00145; 
        10'b1010001011: data <= 17'h00158; 
        10'b1010001100: data <= 17'h00053; 
        10'b1010001101: data <= 17'h000dc; 
        10'b1010001110: data <= 17'h0008c; 
        10'b1010001111: data <= 17'h1fffe; 
        10'b1010010000: data <= 17'h1ff92; 
        10'b1010010001: data <= 17'h00012; 
        10'b1010010010: data <= 17'h0002d; 
        10'b1010010011: data <= 17'h0006e; 
        10'b1010010100: data <= 17'h00052; 
        10'b1010010101: data <= 17'h000aa; 
        10'b1010010110: data <= 17'h0010f; 
        10'b1010010111: data <= 17'h1ffd2; 
        10'b1010011000: data <= 17'h1ff4b; 
        10'b1010011001: data <= 17'h1ff4d; 
        10'b1010011010: data <= 17'h1ffa2; 
        10'b1010011011: data <= 17'h1ff8a; 
        10'b1010011100: data <= 17'h1fff6; 
        10'b1010011101: data <= 17'h1ffe1; 
        10'b1010011110: data <= 17'h1ff90; 
        10'b1010011111: data <= 17'h1ff99; 
        10'b1010100000: data <= 17'h1ffaf; 
        10'b1010100001: data <= 17'h0000d; 
        10'b1010100010: data <= 17'h0000e; 
        10'b1010100011: data <= 17'h00002; 
        10'b1010100100: data <= 17'h000ba; 
        10'b1010100101: data <= 17'h0012b; 
        10'b1010100110: data <= 17'h00161; 
        10'b1010100111: data <= 17'h001a0; 
        10'b1010101000: data <= 17'h001a7; 
        10'b1010101001: data <= 17'h0015b; 
        10'b1010101010: data <= 17'h001f9; 
        10'b1010101011: data <= 17'h00216; 
        10'b1010101100: data <= 17'h00223; 
        10'b1010101101: data <= 17'h001af; 
        10'b1010101110: data <= 17'h0017c; 
        10'b1010101111: data <= 17'h00119; 
        10'b1010110000: data <= 17'h0010c; 
        10'b1010110001: data <= 17'h1ffe9; 
        10'b1010110010: data <= 17'h1ff26; 
        10'b1010110011: data <= 17'h1fed3; 
        10'b1010110100: data <= 17'h1fef1; 
        10'b1010110101: data <= 17'h1ff5b; 
        10'b1010110110: data <= 17'h1ff66; 
        10'b1010110111: data <= 17'h1ffd2; 
        10'b1010111000: data <= 17'h1ffb3; 
        10'b1010111001: data <= 17'h1fffe; 
        10'b1010111010: data <= 17'h1ffb1; 
        10'b1010111011: data <= 17'h0000e; 
        10'b1010111100: data <= 17'h1fff4; 
        10'b1010111101: data <= 17'h1ff7e; 
        10'b1010111110: data <= 17'h0000a; 
        10'b1010111111: data <= 17'h00015; 
        10'b1011000000: data <= 17'h1ffe0; 
        10'b1011000001: data <= 17'h00075; 
        10'b1011000010: data <= 17'h000b0; 
        10'b1011000011: data <= 17'h00062; 
        10'b1011000100: data <= 17'h000ed; 
        10'b1011000101: data <= 17'h000f0; 
        10'b1011000110: data <= 17'h001c0; 
        10'b1011000111: data <= 17'h00200; 
        10'b1011001000: data <= 17'h00226; 
        10'b1011001001: data <= 17'h001ae; 
        10'b1011001010: data <= 17'h00132; 
        10'b1011001011: data <= 17'h0007b; 
        10'b1011001100: data <= 17'h1ffcf; 
        10'b1011001101: data <= 17'h1ff3e; 
        10'b1011001110: data <= 17'h1ff3d; 
        10'b1011001111: data <= 17'h1ff60; 
        10'b1011010000: data <= 17'h1ff62; 
        10'b1011010001: data <= 17'h1ffb0; 
        10'b1011010010: data <= 17'h1ffb0; 
        10'b1011010011: data <= 17'h1fff7; 
        10'b1011010100: data <= 17'h1ff9f; 
        10'b1011010101: data <= 17'h0000c; 
        10'b1011010110: data <= 17'h1ff81; 
        10'b1011010111: data <= 17'h1ffee; 
        10'b1011011000: data <= 17'h1ffa4; 
        10'b1011011001: data <= 17'h1ff7d; 
        10'b1011011010: data <= 17'h1ff83; 
        10'b1011011011: data <= 17'h1ffe0; 
        10'b1011011100: data <= 17'h1ffe2; 
        10'b1011011101: data <= 17'h1ffaa; 
        10'b1011011110: data <= 17'h1ff9c; 
        10'b1011011111: data <= 17'h1ffdd; 
        10'b1011100000: data <= 17'h1ffe0; 
        10'b1011100001: data <= 17'h1ffd6; 
        10'b1011100010: data <= 17'h1ffc5; 
        10'b1011100011: data <= 17'h1ffcf; 
        10'b1011100100: data <= 17'h1ffb7; 
        10'b1011100101: data <= 17'h1ffd9; 
        10'b1011100110: data <= 17'h1ffb7; 
        10'b1011100111: data <= 17'h1ff72; 
        10'b1011101000: data <= 17'h1ffa9; 
        10'b1011101001: data <= 17'h1ffd7; 
        10'b1011101010: data <= 17'h1ffc7; 
        10'b1011101011: data <= 17'h1ffdb; 
        10'b1011101100: data <= 17'h1ff86; 
        10'b1011101101: data <= 17'h1ff88; 
        10'b1011101110: data <= 17'h1ffee; 
        10'b1011101111: data <= 17'h1ffba; 
        10'b1011110000: data <= 17'h00003; 
        10'b1011110001: data <= 17'h1ffa2; 
        10'b1011110010: data <= 17'h1fff6; 
        10'b1011110011: data <= 17'h0000f; 
        10'b1011110100: data <= 17'h1ffc2; 
        10'b1011110101: data <= 17'h1ff9e; 
        10'b1011110110: data <= 17'h1ffd5; 
        10'b1011110111: data <= 17'h1ff85; 
        10'b1011111000: data <= 17'h00006; 
        10'b1011111001: data <= 17'h1ffdf; 
        10'b1011111010: data <= 17'h1fffa; 
        10'b1011111011: data <= 17'h1ffd9; 
        10'b1011111100: data <= 17'h1ffec; 
        10'b1011111101: data <= 17'h1ff84; 
        10'b1011111110: data <= 17'h1ff9a; 
        10'b1011111111: data <= 17'h1ffe5; 
        10'b1100000000: data <= 17'h1ff9a; 
        10'b1100000001: data <= 17'h1ffed; 
        10'b1100000010: data <= 17'h1ffb4; 
        10'b1100000011: data <= 17'h1ffd3; 
        10'b1100000100: data <= 17'h1ffb7; 
        10'b1100000101: data <= 17'h1fffe; 
        10'b1100000110: data <= 17'h1ff8b; 
        10'b1100000111: data <= 17'h1ff9f; 
        10'b1100001000: data <= 17'h1fff8; 
        10'b1100001001: data <= 17'h1ffd5; 
        10'b1100001010: data <= 17'h1ff9e; 
        10'b1100001011: data <= 17'h1ffe2; 
        10'b1100001100: data <= 17'h1ff8c; 
        10'b1100001101: data <= 17'h1ff82; 
        10'b1100001110: data <= 17'h1fff9; 
        10'b1100001111: data <= 17'h1ffc6; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 12) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 18'h3ffaf; 
        10'b0000000001: data <= 18'h3ff39; 
        10'b0000000010: data <= 18'h3fff6; 
        10'b0000000011: data <= 18'h00009; 
        10'b0000000100: data <= 18'h00014; 
        10'b0000000101: data <= 18'h3ffee; 
        10'b0000000110: data <= 18'h3ffb4; 
        10'b0000000111: data <= 18'h00015; 
        10'b0000001000: data <= 18'h3ff5f; 
        10'b0000001001: data <= 18'h0000d; 
        10'b0000001010: data <= 18'h0000e; 
        10'b0000001011: data <= 18'h3ff77; 
        10'b0000001100: data <= 18'h3ff73; 
        10'b0000001101: data <= 18'h3ff70; 
        10'b0000001110: data <= 18'h3ff7b; 
        10'b0000001111: data <= 18'h3ff8c; 
        10'b0000010000: data <= 18'h00003; 
        10'b0000010001: data <= 18'h00009; 
        10'b0000010010: data <= 18'h3ff39; 
        10'b0000010011: data <= 18'h00014; 
        10'b0000010100: data <= 18'h3ffbf; 
        10'b0000010101: data <= 18'h3ffc8; 
        10'b0000010110: data <= 18'h3fefb; 
        10'b0000010111: data <= 18'h3fff2; 
        10'b0000011000: data <= 18'h3fff6; 
        10'b0000011001: data <= 18'h3ff0a; 
        10'b0000011010: data <= 18'h3ff87; 
        10'b0000011011: data <= 18'h00007; 
        10'b0000011100: data <= 18'h3ff32; 
        10'b0000011101: data <= 18'h3ff7f; 
        10'b0000011110: data <= 18'h3ff36; 
        10'b0000011111: data <= 18'h3ffba; 
        10'b0000100000: data <= 18'h3ff18; 
        10'b0000100001: data <= 18'h3ff91; 
        10'b0000100010: data <= 18'h0001b; 
        10'b0000100011: data <= 18'h0000f; 
        10'b0000100100: data <= 18'h3ff09; 
        10'b0000100101: data <= 18'h3fefe; 
        10'b0000100110: data <= 18'h3ff18; 
        10'b0000100111: data <= 18'h3ffb4; 
        10'b0000101000: data <= 18'h3ffc9; 
        10'b0000101001: data <= 18'h3ff8a; 
        10'b0000101010: data <= 18'h3ff76; 
        10'b0000101011: data <= 18'h3ff46; 
        10'b0000101100: data <= 18'h00019; 
        10'b0000101101: data <= 18'h3ff39; 
        10'b0000101110: data <= 18'h3ffd4; 
        10'b0000101111: data <= 18'h3ff69; 
        10'b0000110000: data <= 18'h3ff6c; 
        10'b0000110001: data <= 18'h3ff10; 
        10'b0000110010: data <= 18'h3ff9c; 
        10'b0000110011: data <= 18'h3ffe8; 
        10'b0000110100: data <= 18'h3ff27; 
        10'b0000110101: data <= 18'h3fff3; 
        10'b0000110110: data <= 18'h3ffaa; 
        10'b0000110111: data <= 18'h3ff29; 
        10'b0000111000: data <= 18'h3ff4b; 
        10'b0000111001: data <= 18'h3ff9b; 
        10'b0000111010: data <= 18'h3ff94; 
        10'b0000111011: data <= 18'h3ff3a; 
        10'b0000111100: data <= 18'h3ffc1; 
        10'b0000111101: data <= 18'h3ffd5; 
        10'b0000111110: data <= 18'h3ff57; 
        10'b0000111111: data <= 18'h3ffd2; 
        10'b0001000000: data <= 18'h3ffea; 
        10'b0001000001: data <= 18'h3ff8a; 
        10'b0001000010: data <= 18'h3ff23; 
        10'b0001000011: data <= 18'h3ff29; 
        10'b0001000100: data <= 18'h3ff0e; 
        10'b0001000101: data <= 18'h3ff2e; 
        10'b0001000110: data <= 18'h3ff7b; 
        10'b0001000111: data <= 18'h3ff68; 
        10'b0001001000: data <= 18'h3ff54; 
        10'b0001001001: data <= 18'h3ff4e; 
        10'b0001001010: data <= 18'h3ffd2; 
        10'b0001001011: data <= 18'h3fffb; 
        10'b0001001100: data <= 18'h3ff85; 
        10'b0001001101: data <= 18'h3ff35; 
        10'b0001001110: data <= 18'h00016; 
        10'b0001001111: data <= 18'h3ffef; 
        10'b0001010000: data <= 18'h00001; 
        10'b0001010001: data <= 18'h3ff61; 
        10'b0001010010: data <= 18'h3ff05; 
        10'b0001010011: data <= 18'h3ff8b; 
        10'b0001010100: data <= 18'h0001c; 
        10'b0001010101: data <= 18'h3ffd0; 
        10'b0001010110: data <= 18'h3ff8e; 
        10'b0001010111: data <= 18'h3ffe2; 
        10'b0001011000: data <= 18'h3ffcd; 
        10'b0001011001: data <= 18'h00001; 
        10'b0001011010: data <= 18'h3ffb5; 
        10'b0001011011: data <= 18'h3fff2; 
        10'b0001011100: data <= 18'h3ffe3; 
        10'b0001011101: data <= 18'h3ffa0; 
        10'b0001011110: data <= 18'h00059; 
        10'b0001011111: data <= 18'h00128; 
        10'b0001100000: data <= 18'h00272; 
        10'b0001100001: data <= 18'h00208; 
        10'b0001100010: data <= 18'h00212; 
        10'b0001100011: data <= 18'h00249; 
        10'b0001100100: data <= 18'h00196; 
        10'b0001100101: data <= 18'h001c9; 
        10'b0001100110: data <= 18'h00165; 
        10'b0001100111: data <= 18'h0001b; 
        10'b0001101000: data <= 18'h3ffdc; 
        10'b0001101001: data <= 18'h3fe4c; 
        10'b0001101010: data <= 18'h3ff04; 
        10'b0001101011: data <= 18'h3ffea; 
        10'b0001101100: data <= 18'h0000c; 
        10'b0001101101: data <= 18'h3ff40; 
        10'b0001101110: data <= 18'h3ffa9; 
        10'b0001101111: data <= 18'h3ff58; 
        10'b0001110000: data <= 18'h3ffa6; 
        10'b0001110001: data <= 18'h3fff1; 
        10'b0001110010: data <= 18'h3ffbc; 
        10'b0001110011: data <= 18'h00008; 
        10'b0001110100: data <= 18'h0005f; 
        10'b0001110101: data <= 18'h3ffff; 
        10'b0001110110: data <= 18'h00170; 
        10'b0001110111: data <= 18'h00136; 
        10'b0001111000: data <= 18'h0034e; 
        10'b0001111001: data <= 18'h002d7; 
        10'b0001111010: data <= 18'h00385; 
        10'b0001111011: data <= 18'h0043c; 
        10'b0001111100: data <= 18'h004ea; 
        10'b0001111101: data <= 18'h00544; 
        10'b0001111110: data <= 18'h004bc; 
        10'b0001111111: data <= 18'h00379; 
        10'b0010000000: data <= 18'h001f5; 
        10'b0010000001: data <= 18'h00191; 
        10'b0010000010: data <= 18'h0028f; 
        10'b0010000011: data <= 18'h00050; 
        10'b0010000100: data <= 18'h3fe3f; 
        10'b0010000101: data <= 18'h3fd44; 
        10'b0010000110: data <= 18'h3fdaa; 
        10'b0010000111: data <= 18'h3fdb7; 
        10'b0010001000: data <= 18'h3ffb9; 
        10'b0010001001: data <= 18'h3ff96; 
        10'b0010001010: data <= 18'h3ff67; 
        10'b0010001011: data <= 18'h3ffd8; 
        10'b0010001100: data <= 18'h3ff23; 
        10'b0010001101: data <= 18'h3ff03; 
        10'b0010001110: data <= 18'h3ff43; 
        10'b0010001111: data <= 18'h3ff44; 
        10'b0010010000: data <= 18'h0002f; 
        10'b0010010001: data <= 18'h0017e; 
        10'b0010010010: data <= 18'h002bb; 
        10'b0010010011: data <= 18'h0022e; 
        10'b0010010100: data <= 18'h0027f; 
        10'b0010010101: data <= 18'h00234; 
        10'b0010010110: data <= 18'h001fe; 
        10'b0010010111: data <= 18'h00298; 
        10'b0010011000: data <= 18'h002a3; 
        10'b0010011001: data <= 18'h00329; 
        10'b0010011010: data <= 18'h0008a; 
        10'b0010011011: data <= 18'h0021b; 
        10'b0010011100: data <= 18'h0026f; 
        10'b0010011101: data <= 18'h3ffd0; 
        10'b0010011110: data <= 18'h3ffdf; 
        10'b0010011111: data <= 18'h3fee6; 
        10'b0010100000: data <= 18'h3fe78; 
        10'b0010100001: data <= 18'h3fcbf; 
        10'b0010100010: data <= 18'h3fbd7; 
        10'b0010100011: data <= 18'h3fc7b; 
        10'b0010100100: data <= 18'h3fefb; 
        10'b0010100101: data <= 18'h00001; 
        10'b0010100110: data <= 18'h3ff4c; 
        10'b0010100111: data <= 18'h3ff92; 
        10'b0010101000: data <= 18'h3ff3a; 
        10'b0010101001: data <= 18'h3ff64; 
        10'b0010101010: data <= 18'h3ff54; 
        10'b0010101011: data <= 18'h00051; 
        10'b0010101100: data <= 18'h001d9; 
        10'b0010101101: data <= 18'h00370; 
        10'b0010101110: data <= 18'h002a1; 
        10'b0010101111: data <= 18'h00204; 
        10'b0010110000: data <= 18'h0030d; 
        10'b0010110001: data <= 18'h0027d; 
        10'b0010110010: data <= 18'h00236; 
        10'b0010110011: data <= 18'h0021e; 
        10'b0010110100: data <= 18'h002d5; 
        10'b0010110101: data <= 18'h0040f; 
        10'b0010110110: data <= 18'h002d3; 
        10'b0010110111: data <= 18'h00105; 
        10'b0010111000: data <= 18'h002b0; 
        10'b0010111001: data <= 18'h00276; 
        10'b0010111010: data <= 18'h00258; 
        10'b0010111011: data <= 18'h3fef4; 
        10'b0010111100: data <= 18'h00100; 
        10'b0010111101: data <= 18'h3ff02; 
        10'b0010111110: data <= 18'h3fc6e; 
        10'b0010111111: data <= 18'h3fc6e; 
        10'b0011000000: data <= 18'h3fdd0; 
        10'b0011000001: data <= 18'h3ff8f; 
        10'b0011000010: data <= 18'h3ffe7; 
        10'b0011000011: data <= 18'h3ffa8; 
        10'b0011000100: data <= 18'h0000b; 
        10'b0011000101: data <= 18'h3ffe1; 
        10'b0011000110: data <= 18'h00036; 
        10'b0011000111: data <= 18'h0018b; 
        10'b0011001000: data <= 18'h0040f; 
        10'b0011001001: data <= 18'h0040a; 
        10'b0011001010: data <= 18'h002d8; 
        10'b0011001011: data <= 18'h000cd; 
        10'b0011001100: data <= 18'h000dc; 
        10'b0011001101: data <= 18'h001cf; 
        10'b0011001110: data <= 18'h0008e; 
        10'b0011001111: data <= 18'h000d3; 
        10'b0011010000: data <= 18'h00262; 
        10'b0011010001: data <= 18'h00241; 
        10'b0011010010: data <= 18'h003bc; 
        10'b0011010011: data <= 18'h00232; 
        10'b0011010100: data <= 18'h000ac; 
        10'b0011010101: data <= 18'h001e0; 
        10'b0011010110: data <= 18'h0018e; 
        10'b0011010111: data <= 18'h001b0; 
        10'b0011011000: data <= 18'h001b6; 
        10'b0011011001: data <= 18'h0003e; 
        10'b0011011010: data <= 18'h3fe47; 
        10'b0011011011: data <= 18'h3fbfe; 
        10'b0011011100: data <= 18'h3fd20; 
        10'b0011011101: data <= 18'h3ff3f; 
        10'b0011011110: data <= 18'h3ff04; 
        10'b0011011111: data <= 18'h3ff7a; 
        10'b0011100000: data <= 18'h3ff9e; 
        10'b0011100001: data <= 18'h3ff69; 
        10'b0011100010: data <= 18'h0002c; 
        10'b0011100011: data <= 18'h00171; 
        10'b0011100100: data <= 18'h00359; 
        10'b0011100101: data <= 18'h0032e; 
        10'b0011100110: data <= 18'h00264; 
        10'b0011100111: data <= 18'h000fa; 
        10'b0011101000: data <= 18'h0019e; 
        10'b0011101001: data <= 18'h000c5; 
        10'b0011101010: data <= 18'h0020b; 
        10'b0011101011: data <= 18'h000a8; 
        10'b0011101100: data <= 18'h0008f; 
        10'b0011101101: data <= 18'h00100; 
        10'b0011101110: data <= 18'h00410; 
        10'b0011101111: data <= 18'h0035f; 
        10'b0011110000: data <= 18'h000c7; 
        10'b0011110001: data <= 18'h001df; 
        10'b0011110010: data <= 18'h002b1; 
        10'b0011110011: data <= 18'h001c1; 
        10'b0011110100: data <= 18'h00291; 
        10'b0011110101: data <= 18'h00152; 
        10'b0011110110: data <= 18'h3ff50; 
        10'b0011110111: data <= 18'h3fc49; 
        10'b0011111000: data <= 18'h3fd38; 
        10'b0011111001: data <= 18'h3fefc; 
        10'b0011111010: data <= 18'h3ff23; 
        10'b0011111011: data <= 18'h3ff61; 
        10'b0011111100: data <= 18'h3ff83; 
        10'b0011111101: data <= 18'h3ff0c; 
        10'b0011111110: data <= 18'h3ffb2; 
        10'b0011111111: data <= 18'h0009f; 
        10'b0100000000: data <= 18'h001bb; 
        10'b0100000001: data <= 18'h0024b; 
        10'b0100000010: data <= 18'h001e6; 
        10'b0100000011: data <= 18'h00076; 
        10'b0100000100: data <= 18'h3ffc2; 
        10'b0100000101: data <= 18'h3fe3a; 
        10'b0100000110: data <= 18'h3fc9f; 
        10'b0100000111: data <= 18'h3f9cc; 
        10'b0100001000: data <= 18'h3faf8; 
        10'b0100001001: data <= 18'h3ff54; 
        10'b0100001010: data <= 18'h004d7; 
        10'b0100001011: data <= 18'h00770; 
        10'b0100001100: data <= 18'h0044c; 
        10'b0100001101: data <= 18'h00283; 
        10'b0100001110: data <= 18'h002bb; 
        10'b0100001111: data <= 18'h00286; 
        10'b0100010000: data <= 18'h003c8; 
        10'b0100010001: data <= 18'h0026a; 
        10'b0100010010: data <= 18'h3ff45; 
        10'b0100010011: data <= 18'h3fc50; 
        10'b0100010100: data <= 18'h3fe25; 
        10'b0100010101: data <= 18'h3fef4; 
        10'b0100010110: data <= 18'h3ff36; 
        10'b0100010111: data <= 18'h3ff58; 
        10'b0100011000: data <= 18'h3ffe5; 
        10'b0100011001: data <= 18'h3ffd8; 
        10'b0100011010: data <= 18'h0000d; 
        10'b0100011011: data <= 18'h000ef; 
        10'b0100011100: data <= 18'h000d7; 
        10'b0100011101: data <= 18'h0005b; 
        10'b0100011110: data <= 18'h3feeb; 
        10'b0100011111: data <= 18'h3fd43; 
        10'b0100100000: data <= 18'h3fafd; 
        10'b0100100001: data <= 18'h3f8d7; 
        10'b0100100010: data <= 18'h3f739; 
        10'b0100100011: data <= 18'h3f700; 
        10'b0100100100: data <= 18'h3f95f; 
        10'b0100100101: data <= 18'h3fe54; 
        10'b0100100110: data <= 18'h003f8; 
        10'b0100100111: data <= 18'h00496; 
        10'b0100101000: data <= 18'h003e8; 
        10'b0100101001: data <= 18'h003a4; 
        10'b0100101010: data <= 18'h0023f; 
        10'b0100101011: data <= 18'h003e6; 
        10'b0100101100: data <= 18'h0039e; 
        10'b0100101101: data <= 18'h00173; 
        10'b0100101110: data <= 18'h3feb4; 
        10'b0100101111: data <= 18'h3fd9b; 
        10'b0100110000: data <= 18'h3ff1b; 
        10'b0100110001: data <= 18'h3fefd; 
        10'b0100110010: data <= 18'h3ff92; 
        10'b0100110011: data <= 18'h3ffe4; 
        10'b0100110100: data <= 18'h0001e; 
        10'b0100110101: data <= 18'h3ffe4; 
        10'b0100110110: data <= 18'h3ff2c; 
        10'b0100110111: data <= 18'h000e8; 
        10'b0100111000: data <= 18'h3ff76; 
        10'b0100111001: data <= 18'h3fd31; 
        10'b0100111010: data <= 18'h3fbca; 
        10'b0100111011: data <= 18'h3f9cf; 
        10'b0100111100: data <= 18'h3f842; 
        10'b0100111101: data <= 18'h3f950; 
        10'b0100111110: data <= 18'h3fae8; 
        10'b0100111111: data <= 18'h3fd99; 
        10'b0101000000: data <= 18'h3feb3; 
        10'b0101000001: data <= 18'h001ae; 
        10'b0101000010: data <= 18'h002a4; 
        10'b0101000011: data <= 18'h002a7; 
        10'b0101000100: data <= 18'h00136; 
        10'b0101000101: data <= 18'h002c0; 
        10'b0101000110: data <= 18'h00367; 
        10'b0101000111: data <= 18'h00351; 
        10'b0101001000: data <= 18'h002e5; 
        10'b0101001001: data <= 18'h00003; 
        10'b0101001010: data <= 18'h3feba; 
        10'b0101001011: data <= 18'h3feef; 
        10'b0101001100: data <= 18'h3ff10; 
        10'b0101001101: data <= 18'h3ff72; 
        10'b0101001110: data <= 18'h3ff3b; 
        10'b0101001111: data <= 18'h3ff23; 
        10'b0101010000: data <= 18'h00009; 
        10'b0101010001: data <= 18'h3ff5a; 
        10'b0101010010: data <= 18'h3ffd6; 
        10'b0101010011: data <= 18'h3fff3; 
        10'b0101010100: data <= 18'h3fefb; 
        10'b0101010101: data <= 18'h3fd2e; 
        10'b0101010110: data <= 18'h3fb11; 
        10'b0101010111: data <= 18'h3f9d4; 
        10'b0101011000: data <= 18'h3fa6b; 
        10'b0101011001: data <= 18'h3fd07; 
        10'b0101011010: data <= 18'h0000f; 
        10'b0101011011: data <= 18'h0007f; 
        10'b0101011100: data <= 18'h000c9; 
        10'b0101011101: data <= 18'h001c9; 
        10'b0101011110: data <= 18'h0046b; 
        10'b0101011111: data <= 18'h00249; 
        10'b0101100000: data <= 18'h0018f; 
        10'b0101100001: data <= 18'h00235; 
        10'b0101100010: data <= 18'h001c4; 
        10'b0101100011: data <= 18'h3ffd9; 
        10'b0101100100: data <= 18'h3fdb6; 
        10'b0101100101: data <= 18'h3fcdc; 
        10'b0101100110: data <= 18'h3fcb6; 
        10'b0101100111: data <= 18'h3fde9; 
        10'b0101101000: data <= 18'h3ffa2; 
        10'b0101101001: data <= 18'h3ff5e; 
        10'b0101101010: data <= 18'h3ffa9; 
        10'b0101101011: data <= 18'h3ffc2; 
        10'b0101101100: data <= 18'h3ff8e; 
        10'b0101101101: data <= 18'h3ff53; 
        10'b0101101110: data <= 18'h3ff96; 
        10'b0101101111: data <= 18'h3ffb9; 
        10'b0101110000: data <= 18'h3feb2; 
        10'b0101110001: data <= 18'h3fe13; 
        10'b0101110010: data <= 18'h3fbfd; 
        10'b0101110011: data <= 18'h3fb5e; 
        10'b0101110100: data <= 18'h3fcdb; 
        10'b0101110101: data <= 18'h3ff62; 
        10'b0101110110: data <= 18'h3fefa; 
        10'b0101110111: data <= 18'h3fd56; 
        10'b0101111000: data <= 18'h00036; 
        10'b0101111001: data <= 18'h003ce; 
        10'b0101111010: data <= 18'h003d8; 
        10'b0101111011: data <= 18'h000b4; 
        10'b0101111100: data <= 18'h001be; 
        10'b0101111101: data <= 18'h001dc; 
        10'b0101111110: data <= 18'h000fd; 
        10'b0101111111: data <= 18'h3feb1; 
        10'b0110000000: data <= 18'h3fc7e; 
        10'b0110000001: data <= 18'h3fc7a; 
        10'b0110000010: data <= 18'h3fd38; 
        10'b0110000011: data <= 18'h3fe0c; 
        10'b0110000100: data <= 18'h3fee1; 
        10'b0110000101: data <= 18'h3fffa; 
        10'b0110000110: data <= 18'h3ffcc; 
        10'b0110000111: data <= 18'h3ff67; 
        10'b0110001000: data <= 18'h00018; 
        10'b0110001001: data <= 18'h3ff3d; 
        10'b0110001010: data <= 18'h3ff83; 
        10'b0110001011: data <= 18'h3ffaf; 
        10'b0110001100: data <= 18'h3ffc2; 
        10'b0110001101: data <= 18'h3fe63; 
        10'b0110001110: data <= 18'h3fc61; 
        10'b0110001111: data <= 18'h3fcba; 
        10'b0110010000: data <= 18'h3fdc7; 
        10'b0110010001: data <= 18'h3ffb1; 
        10'b0110010010: data <= 18'h3fdab; 
        10'b0110010011: data <= 18'h3fd84; 
        10'b0110010100: data <= 18'h000b4; 
        10'b0110010101: data <= 18'h001d7; 
        10'b0110010110: data <= 18'h001f7; 
        10'b0110010111: data <= 18'h3ffb5; 
        10'b0110011000: data <= 18'h3ff34; 
        10'b0110011001: data <= 18'h3ff68; 
        10'b0110011010: data <= 18'h00045; 
        10'b0110011011: data <= 18'h3fe7a; 
        10'b0110011100: data <= 18'h3fdf0; 
        10'b0110011101: data <= 18'h3ff00; 
        10'b0110011110: data <= 18'h3fe94; 
        10'b0110011111: data <= 18'h3ff0b; 
        10'b0110100000: data <= 18'h3febd; 
        10'b0110100001: data <= 18'h3fedd; 
        10'b0110100010: data <= 18'h00007; 
        10'b0110100011: data <= 18'h0000e; 
        10'b0110100100: data <= 18'h00015; 
        10'b0110100101: data <= 18'h3ff40; 
        10'b0110100110: data <= 18'h0001d; 
        10'b0110100111: data <= 18'h00047; 
        10'b0110101000: data <= 18'h3ffad; 
        10'b0110101001: data <= 18'h3fe31; 
        10'b0110101010: data <= 18'h3fca4; 
        10'b0110101011: data <= 18'h3fc68; 
        10'b0110101100: data <= 18'h3fd4f; 
        10'b0110101101: data <= 18'h3fe6c; 
        10'b0110101110: data <= 18'h3fe41; 
        10'b0110101111: data <= 18'h3ff69; 
        10'b0110110000: data <= 18'h000ba; 
        10'b0110110001: data <= 18'h002fe; 
        10'b0110110010: data <= 18'h001b8; 
        10'b0110110011: data <= 18'h3ffd5; 
        10'b0110110100: data <= 18'h3fd81; 
        10'b0110110101: data <= 18'h3ff46; 
        10'b0110110110: data <= 18'h3ffc1; 
        10'b0110110111: data <= 18'h000a8; 
        10'b0110111000: data <= 18'h0018d; 
        10'b0110111001: data <= 18'h00184; 
        10'b0110111010: data <= 18'h00086; 
        10'b0110111011: data <= 18'h00033; 
        10'b0110111100: data <= 18'h3ff0d; 
        10'b0110111101: data <= 18'h3ffca; 
        10'b0110111110: data <= 18'h3ffb3; 
        10'b0110111111: data <= 18'h3ff3f; 
        10'b0111000000: data <= 18'h3ffb7; 
        10'b0111000001: data <= 18'h3ffd7; 
        10'b0111000010: data <= 18'h000b0; 
        10'b0111000011: data <= 18'h0001f; 
        10'b0111000100: data <= 18'h00081; 
        10'b0111000101: data <= 18'h3ff2a; 
        10'b0111000110: data <= 18'h3fea1; 
        10'b0111000111: data <= 18'h3fda0; 
        10'b0111001000: data <= 18'h3fad4; 
        10'b0111001001: data <= 18'h3fa8d; 
        10'b0111001010: data <= 18'h3fb2b; 
        10'b0111001011: data <= 18'h3fec7; 
        10'b0111001100: data <= 18'h00171; 
        10'b0111001101: data <= 18'h003bb; 
        10'b0111001110: data <= 18'h3ff99; 
        10'b0111001111: data <= 18'h3fd47; 
        10'b0111010000: data <= 18'h3fd1f; 
        10'b0111010001: data <= 18'h3ff10; 
        10'b0111010010: data <= 18'h00137; 
        10'b0111010011: data <= 18'h0032f; 
        10'b0111010100: data <= 18'h0023d; 
        10'b0111010101: data <= 18'h002d2; 
        10'b0111010110: data <= 18'h002bd; 
        10'b0111010111: data <= 18'h00136; 
        10'b0111011000: data <= 18'h3ffa4; 
        10'b0111011001: data <= 18'h3ffc2; 
        10'b0111011010: data <= 18'h3fff8; 
        10'b0111011011: data <= 18'h3ffe9; 
        10'b0111011100: data <= 18'h3ffe4; 
        10'b0111011101: data <= 18'h0001e; 
        10'b0111011110: data <= 18'h00004; 
        10'b0111011111: data <= 18'h001be; 
        10'b0111100000: data <= 18'h000f7; 
        10'b0111100001: data <= 18'h0004d; 
        10'b0111100010: data <= 18'h3ff14; 
        10'b0111100011: data <= 18'h3fcdd; 
        10'b0111100100: data <= 18'h3fa69; 
        10'b0111100101: data <= 18'h3f723; 
        10'b0111100110: data <= 18'h3f4f9; 
        10'b0111100111: data <= 18'h3f5ef; 
        10'b0111101000: data <= 18'h3f85b; 
        10'b0111101001: data <= 18'h3fba5; 
        10'b0111101010: data <= 18'h3fbf6; 
        10'b0111101011: data <= 18'h3fc65; 
        10'b0111101100: data <= 18'h3ffdb; 
        10'b0111101101: data <= 18'h0011d; 
        10'b0111101110: data <= 18'h0020a; 
        10'b0111101111: data <= 18'h0033a; 
        10'b0111110000: data <= 18'h000ab; 
        10'b0111110001: data <= 18'h003e8; 
        10'b0111110010: data <= 18'h003e6; 
        10'b0111110011: data <= 18'h0012c; 
        10'b0111110100: data <= 18'h3ff6c; 
        10'b0111110101: data <= 18'h3ff2b; 
        10'b0111110110: data <= 18'h3ff3e; 
        10'b0111110111: data <= 18'h3ff4f; 
        10'b0111111000: data <= 18'h3ff93; 
        10'b0111111001: data <= 18'h3ff99; 
        10'b0111111010: data <= 18'h00057; 
        10'b0111111011: data <= 18'h00294; 
        10'b0111111100: data <= 18'h001dc; 
        10'b0111111101: data <= 18'h0011f; 
        10'b0111111110: data <= 18'h00096; 
        10'b0111111111: data <= 18'h3ff52; 
        10'b1000000000: data <= 18'h3fe03; 
        10'b1000000001: data <= 18'h3f983; 
        10'b1000000010: data <= 18'h3f672; 
        10'b1000000011: data <= 18'h3f6f6; 
        10'b1000000100: data <= 18'h3f515; 
        10'b1000000101: data <= 18'h3f717; 
        10'b1000000110: data <= 18'h3fa5d; 
        10'b1000000111: data <= 18'h3feb8; 
        10'b1000001000: data <= 18'h00246; 
        10'b1000001001: data <= 18'h00311; 
        10'b1000001010: data <= 18'h0034e; 
        10'b1000001011: data <= 18'h00345; 
        10'b1000001100: data <= 18'h0024a; 
        10'b1000001101: data <= 18'h00490; 
        10'b1000001110: data <= 18'h00442; 
        10'b1000001111: data <= 18'h001a0; 
        10'b1000010000: data <= 18'h3fe80; 
        10'b1000010001: data <= 18'h3fefc; 
        10'b1000010010: data <= 18'h3ff43; 
        10'b1000010011: data <= 18'h3ffe2; 
        10'b1000010100: data <= 18'h3ffe2; 
        10'b1000010101: data <= 18'h3ff41; 
        10'b1000010110: data <= 18'h3ff86; 
        10'b1000010111: data <= 18'h0033c; 
        10'b1000011000: data <= 18'h0034d; 
        10'b1000011001: data <= 18'h003e0; 
        10'b1000011010: data <= 18'h00357; 
        10'b1000011011: data <= 18'h0013a; 
        10'b1000011100: data <= 18'h0005e; 
        10'b1000011101: data <= 18'h3fea3; 
        10'b1000011110: data <= 18'h3ff05; 
        10'b1000011111: data <= 18'h3fcec; 
        10'b1000100000: data <= 18'h3fb80; 
        10'b1000100001: data <= 18'h3fb37; 
        10'b1000100010: data <= 18'h3fcbd; 
        10'b1000100011: data <= 18'h00126; 
        10'b1000100100: data <= 18'h00314; 
        10'b1000100101: data <= 18'h003da; 
        10'b1000100110: data <= 18'h00451; 
        10'b1000100111: data <= 18'h003dc; 
        10'b1000101000: data <= 18'h0036a; 
        10'b1000101001: data <= 18'h003fc; 
        10'b1000101010: data <= 18'h00187; 
        10'b1000101011: data <= 18'h0002e; 
        10'b1000101100: data <= 18'h3febc; 
        10'b1000101101: data <= 18'h3ffc4; 
        10'b1000101110: data <= 18'h3ffe0; 
        10'b1000101111: data <= 18'h3ffbb; 
        10'b1000110000: data <= 18'h3ffd6; 
        10'b1000110001: data <= 18'h3ff04; 
        10'b1000110010: data <= 18'h00095; 
        10'b1000110011: data <= 18'h00379; 
        10'b1000110100: data <= 18'h00444; 
        10'b1000110101: data <= 18'h0049e; 
        10'b1000110110: data <= 18'h004e4; 
        10'b1000110111: data <= 18'h00278; 
        10'b1000111000: data <= 18'h002e7; 
        10'b1000111001: data <= 18'h00349; 
        10'b1000111010: data <= 18'h00136; 
        10'b1000111011: data <= 18'h3ffab; 
        10'b1000111100: data <= 18'h3fee6; 
        10'b1000111101: data <= 18'h3fe50; 
        10'b1000111110: data <= 18'h00083; 
        10'b1000111111: data <= 18'h000e9; 
        10'b1001000000: data <= 18'h001bd; 
        10'b1001000001: data <= 18'h00318; 
        10'b1001000010: data <= 18'h0033e; 
        10'b1001000011: data <= 18'h00235; 
        10'b1001000100: data <= 18'h003d7; 
        10'b1001000101: data <= 18'h0022f; 
        10'b1001000110: data <= 18'h3ff98; 
        10'b1001000111: data <= 18'h3ff20; 
        10'b1001001000: data <= 18'h3fefc; 
        10'b1001001001: data <= 18'h3ffb3; 
        10'b1001001010: data <= 18'h3ffb0; 
        10'b1001001011: data <= 18'h3ffa7; 
        10'b1001001100: data <= 18'h3ff56; 
        10'b1001001101: data <= 18'h3fff4; 
        10'b1001001110: data <= 18'h3ffc2; 
        10'b1001001111: data <= 18'h001ba; 
        10'b1001010000: data <= 18'h0041e; 
        10'b1001010001: data <= 18'h0041d; 
        10'b1001010010: data <= 18'h00398; 
        10'b1001010011: data <= 18'h00207; 
        10'b1001010100: data <= 18'h0022a; 
        10'b1001010101: data <= 18'h000b7; 
        10'b1001010110: data <= 18'h3ffb7; 
        10'b1001010111: data <= 18'h3ff07; 
        10'b1001011000: data <= 18'h00050; 
        10'b1001011001: data <= 18'h3ffd3; 
        10'b1001011010: data <= 18'h3ffbf; 
        10'b1001011011: data <= 18'h3ff87; 
        10'b1001011100: data <= 18'h00102; 
        10'b1001011101: data <= 18'h0005e; 
        10'b1001011110: data <= 18'h001fa; 
        10'b1001011111: data <= 18'h0032e; 
        10'b1001100000: data <= 18'h001da; 
        10'b1001100001: data <= 18'h000b5; 
        10'b1001100010: data <= 18'h3ff48; 
        10'b1001100011: data <= 18'h3fe27; 
        10'b1001100100: data <= 18'h3ff66; 
        10'b1001100101: data <= 18'h3ff3d; 
        10'b1001100110: data <= 18'h3feff; 
        10'b1001100111: data <= 18'h3ff0f; 
        10'b1001101000: data <= 18'h3ff96; 
        10'b1001101001: data <= 18'h3ffb6; 
        10'b1001101010: data <= 18'h3ffcf; 
        10'b1001101011: data <= 18'h00113; 
        10'b1001101100: data <= 18'h00212; 
        10'b1001101101: data <= 18'h002d1; 
        10'b1001101110: data <= 18'h00283; 
        10'b1001101111: data <= 18'h0016e; 
        10'b1001110000: data <= 18'h0001c; 
        10'b1001110001: data <= 18'h00109; 
        10'b1001110010: data <= 18'h00140; 
        10'b1001110011: data <= 18'h00185; 
        10'b1001110100: data <= 18'h0006c; 
        10'b1001110101: data <= 18'h3ff72; 
        10'b1001110110: data <= 18'h3ff69; 
        10'b1001110111: data <= 18'h3ff2a; 
        10'b1001111000: data <= 18'h000a8; 
        10'b1001111001: data <= 18'h00080; 
        10'b1001111010: data <= 18'h0007e; 
        10'b1001111011: data <= 18'h00233; 
        10'b1001111100: data <= 18'h00111; 
        10'b1001111101: data <= 18'h3ff9f; 
        10'b1001111110: data <= 18'h3ff82; 
        10'b1001111111: data <= 18'h3ff5b; 
        10'b1010000000: data <= 18'h3fe96; 
        10'b1010000001: data <= 18'h3fef1; 
        10'b1010000010: data <= 18'h3ffcf; 
        10'b1010000011: data <= 18'h3fff8; 
        10'b1010000100: data <= 18'h3ffb5; 
        10'b1010000101: data <= 18'h3ff35; 
        10'b1010000110: data <= 18'h3ff57; 
        10'b1010000111: data <= 18'h000b5; 
        10'b1010001000: data <= 18'h00242; 
        10'b1010001001: data <= 18'h00369; 
        10'b1010001010: data <= 18'h0028b; 
        10'b1010001011: data <= 18'h002af; 
        10'b1010001100: data <= 18'h000a6; 
        10'b1010001101: data <= 18'h001b8; 
        10'b1010001110: data <= 18'h00118; 
        10'b1010001111: data <= 18'h3fffc; 
        10'b1010010000: data <= 18'h3ff23; 
        10'b1010010001: data <= 18'h00023; 
        10'b1010010010: data <= 18'h00059; 
        10'b1010010011: data <= 18'h000dc; 
        10'b1010010100: data <= 18'h000a4; 
        10'b1010010101: data <= 18'h00154; 
        10'b1010010110: data <= 18'h0021e; 
        10'b1010010111: data <= 18'h3ffa5; 
        10'b1010011000: data <= 18'h3fe96; 
        10'b1010011001: data <= 18'h3fe99; 
        10'b1010011010: data <= 18'h3ff43; 
        10'b1010011011: data <= 18'h3ff13; 
        10'b1010011100: data <= 18'h3ffeb; 
        10'b1010011101: data <= 18'h3ffc3; 
        10'b1010011110: data <= 18'h3ff1f; 
        10'b1010011111: data <= 18'h3ff33; 
        10'b1010100000: data <= 18'h3ff5e; 
        10'b1010100001: data <= 18'h0001a; 
        10'b1010100010: data <= 18'h0001b; 
        10'b1010100011: data <= 18'h00003; 
        10'b1010100100: data <= 18'h00174; 
        10'b1010100101: data <= 18'h00257; 
        10'b1010100110: data <= 18'h002c1; 
        10'b1010100111: data <= 18'h00340; 
        10'b1010101000: data <= 18'h0034e; 
        10'b1010101001: data <= 18'h002b6; 
        10'b1010101010: data <= 18'h003f3; 
        10'b1010101011: data <= 18'h0042b; 
        10'b1010101100: data <= 18'h00445; 
        10'b1010101101: data <= 18'h0035d; 
        10'b1010101110: data <= 18'h002f7; 
        10'b1010101111: data <= 18'h00232; 
        10'b1010110000: data <= 18'h00218; 
        10'b1010110001: data <= 18'h3ffd1; 
        10'b1010110010: data <= 18'h3fe4c; 
        10'b1010110011: data <= 18'h3fda5; 
        10'b1010110100: data <= 18'h3fde2; 
        10'b1010110101: data <= 18'h3feb5; 
        10'b1010110110: data <= 18'h3fecb; 
        10'b1010110111: data <= 18'h3ffa5; 
        10'b1010111000: data <= 18'h3ff66; 
        10'b1010111001: data <= 18'h3fffc; 
        10'b1010111010: data <= 18'h3ff63; 
        10'b1010111011: data <= 18'h0001c; 
        10'b1010111100: data <= 18'h3ffe8; 
        10'b1010111101: data <= 18'h3fefd; 
        10'b1010111110: data <= 18'h00014; 
        10'b1010111111: data <= 18'h0002a; 
        10'b1011000000: data <= 18'h3ffc0; 
        10'b1011000001: data <= 18'h000ea; 
        10'b1011000010: data <= 18'h00160; 
        10'b1011000011: data <= 18'h000c5; 
        10'b1011000100: data <= 18'h001da; 
        10'b1011000101: data <= 18'h001df; 
        10'b1011000110: data <= 18'h00380; 
        10'b1011000111: data <= 18'h00400; 
        10'b1011001000: data <= 18'h0044b; 
        10'b1011001001: data <= 18'h0035d; 
        10'b1011001010: data <= 18'h00264; 
        10'b1011001011: data <= 18'h000f6; 
        10'b1011001100: data <= 18'h3ff9d; 
        10'b1011001101: data <= 18'h3fe7c; 
        10'b1011001110: data <= 18'h3fe7a; 
        10'b1011001111: data <= 18'h3fec1; 
        10'b1011010000: data <= 18'h3fec3; 
        10'b1011010001: data <= 18'h3ff60; 
        10'b1011010010: data <= 18'h3ff60; 
        10'b1011010011: data <= 18'h3ffef; 
        10'b1011010100: data <= 18'h3ff3e; 
        10'b1011010101: data <= 18'h00019; 
        10'b1011010110: data <= 18'h3ff02; 
        10'b1011010111: data <= 18'h3ffdc; 
        10'b1011011000: data <= 18'h3ff48; 
        10'b1011011001: data <= 18'h3fefa; 
        10'b1011011010: data <= 18'h3ff06; 
        10'b1011011011: data <= 18'h3ffc0; 
        10'b1011011100: data <= 18'h3ffc4; 
        10'b1011011101: data <= 18'h3ff53; 
        10'b1011011110: data <= 18'h3ff37; 
        10'b1011011111: data <= 18'h3ffba; 
        10'b1011100000: data <= 18'h3ffc0; 
        10'b1011100001: data <= 18'h3ffac; 
        10'b1011100010: data <= 18'h3ff8b; 
        10'b1011100011: data <= 18'h3ff9e; 
        10'b1011100100: data <= 18'h3ff6f; 
        10'b1011100101: data <= 18'h3ffb2; 
        10'b1011100110: data <= 18'h3ff6d; 
        10'b1011100111: data <= 18'h3fee5; 
        10'b1011101000: data <= 18'h3ff52; 
        10'b1011101001: data <= 18'h3ffae; 
        10'b1011101010: data <= 18'h3ff8e; 
        10'b1011101011: data <= 18'h3ffb6; 
        10'b1011101100: data <= 18'h3ff0b; 
        10'b1011101101: data <= 18'h3ff10; 
        10'b1011101110: data <= 18'h3ffdb; 
        10'b1011101111: data <= 18'h3ff74; 
        10'b1011110000: data <= 18'h00006; 
        10'b1011110001: data <= 18'h3ff44; 
        10'b1011110010: data <= 18'h3ffeb; 
        10'b1011110011: data <= 18'h0001d; 
        10'b1011110100: data <= 18'h3ff83; 
        10'b1011110101: data <= 18'h3ff3c; 
        10'b1011110110: data <= 18'h3ffaa; 
        10'b1011110111: data <= 18'h3ff0b; 
        10'b1011111000: data <= 18'h0000d; 
        10'b1011111001: data <= 18'h3ffbd; 
        10'b1011111010: data <= 18'h3fff3; 
        10'b1011111011: data <= 18'h3ffb2; 
        10'b1011111100: data <= 18'h3ffd8; 
        10'b1011111101: data <= 18'h3ff07; 
        10'b1011111110: data <= 18'h3ff34; 
        10'b1011111111: data <= 18'h3ffca; 
        10'b1100000000: data <= 18'h3ff33; 
        10'b1100000001: data <= 18'h3ffda; 
        10'b1100000010: data <= 18'h3ff67; 
        10'b1100000011: data <= 18'h3ffa6; 
        10'b1100000100: data <= 18'h3ff6e; 
        10'b1100000101: data <= 18'h3fffb; 
        10'b1100000110: data <= 18'h3ff15; 
        10'b1100000111: data <= 18'h3ff3e; 
        10'b1100001000: data <= 18'h3fff0; 
        10'b1100001001: data <= 18'h3ffab; 
        10'b1100001010: data <= 18'h3ff3c; 
        10'b1100001011: data <= 18'h3ffc3; 
        10'b1100001100: data <= 18'h3ff18; 
        10'b1100001101: data <= 18'h3ff05; 
        10'b1100001110: data <= 18'h3fff2; 
        10'b1100001111: data <= 18'h3ff8b; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 13) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 19'h7ff5f; 
        10'b0000000001: data <= 19'h7fe71; 
        10'b0000000010: data <= 19'h7ffec; 
        10'b0000000011: data <= 19'h00012; 
        10'b0000000100: data <= 19'h00028; 
        10'b0000000101: data <= 19'h7ffdd; 
        10'b0000000110: data <= 19'h7ff68; 
        10'b0000000111: data <= 19'h00029; 
        10'b0000001000: data <= 19'h7febe; 
        10'b0000001001: data <= 19'h00019; 
        10'b0000001010: data <= 19'h0001b; 
        10'b0000001011: data <= 19'h7feee; 
        10'b0000001100: data <= 19'h7fee7; 
        10'b0000001101: data <= 19'h7fee0; 
        10'b0000001110: data <= 19'h7fef6; 
        10'b0000001111: data <= 19'h7ff18; 
        10'b0000010000: data <= 19'h00005; 
        10'b0000010001: data <= 19'h00012; 
        10'b0000010010: data <= 19'h7fe72; 
        10'b0000010011: data <= 19'h00029; 
        10'b0000010100: data <= 19'h7ff7f; 
        10'b0000010101: data <= 19'h7ff90; 
        10'b0000010110: data <= 19'h7fdf6; 
        10'b0000010111: data <= 19'h7ffe3; 
        10'b0000011000: data <= 19'h7ffed; 
        10'b0000011001: data <= 19'h7fe15; 
        10'b0000011010: data <= 19'h7ff0e; 
        10'b0000011011: data <= 19'h0000e; 
        10'b0000011100: data <= 19'h7fe65; 
        10'b0000011101: data <= 19'h7fefe; 
        10'b0000011110: data <= 19'h7fe6c; 
        10'b0000011111: data <= 19'h7ff73; 
        10'b0000100000: data <= 19'h7fe30; 
        10'b0000100001: data <= 19'h7ff22; 
        10'b0000100010: data <= 19'h00035; 
        10'b0000100011: data <= 19'h0001d; 
        10'b0000100100: data <= 19'h7fe12; 
        10'b0000100101: data <= 19'h7fdfb; 
        10'b0000100110: data <= 19'h7fe30; 
        10'b0000100111: data <= 19'h7ff67; 
        10'b0000101000: data <= 19'h7ff92; 
        10'b0000101001: data <= 19'h7ff14; 
        10'b0000101010: data <= 19'h7feec; 
        10'b0000101011: data <= 19'h7fe8c; 
        10'b0000101100: data <= 19'h00033; 
        10'b0000101101: data <= 19'h7fe73; 
        10'b0000101110: data <= 19'h7ffa8; 
        10'b0000101111: data <= 19'h7fed1; 
        10'b0000110000: data <= 19'h7fed8; 
        10'b0000110001: data <= 19'h7fe20; 
        10'b0000110010: data <= 19'h7ff38; 
        10'b0000110011: data <= 19'h7ffd0; 
        10'b0000110100: data <= 19'h7fe4e; 
        10'b0000110101: data <= 19'h7ffe7; 
        10'b0000110110: data <= 19'h7ff55; 
        10'b0000110111: data <= 19'h7fe52; 
        10'b0000111000: data <= 19'h7fe96; 
        10'b0000111001: data <= 19'h7ff35; 
        10'b0000111010: data <= 19'h7ff27; 
        10'b0000111011: data <= 19'h7fe73; 
        10'b0000111100: data <= 19'h7ff82; 
        10'b0000111101: data <= 19'h7ffab; 
        10'b0000111110: data <= 19'h7feae; 
        10'b0000111111: data <= 19'h7ffa4; 
        10'b0001000000: data <= 19'h7ffd3; 
        10'b0001000001: data <= 19'h7ff14; 
        10'b0001000010: data <= 19'h7fe46; 
        10'b0001000011: data <= 19'h7fe52; 
        10'b0001000100: data <= 19'h7fe1c; 
        10'b0001000101: data <= 19'h7fe5c; 
        10'b0001000110: data <= 19'h7fef6; 
        10'b0001000111: data <= 19'h7fed0; 
        10'b0001001000: data <= 19'h7fea8; 
        10'b0001001001: data <= 19'h7fe9c; 
        10'b0001001010: data <= 19'h7ffa4; 
        10'b0001001011: data <= 19'h7fff5; 
        10'b0001001100: data <= 19'h7ff09; 
        10'b0001001101: data <= 19'h7fe69; 
        10'b0001001110: data <= 19'h0002d; 
        10'b0001001111: data <= 19'h7ffdf; 
        10'b0001010000: data <= 19'h00001; 
        10'b0001010001: data <= 19'h7fec2; 
        10'b0001010010: data <= 19'h7fe0a; 
        10'b0001010011: data <= 19'h7ff16; 
        10'b0001010100: data <= 19'h00038; 
        10'b0001010101: data <= 19'h7ffa0; 
        10'b0001010110: data <= 19'h7ff1d; 
        10'b0001010111: data <= 19'h7ffc3; 
        10'b0001011000: data <= 19'h7ff9a; 
        10'b0001011001: data <= 19'h00002; 
        10'b0001011010: data <= 19'h7ff6a; 
        10'b0001011011: data <= 19'h7ffe4; 
        10'b0001011100: data <= 19'h7ffc6; 
        10'b0001011101: data <= 19'h7ff41; 
        10'b0001011110: data <= 19'h000b2; 
        10'b0001011111: data <= 19'h00251; 
        10'b0001100000: data <= 19'h004e4; 
        10'b0001100001: data <= 19'h00410; 
        10'b0001100010: data <= 19'h00424; 
        10'b0001100011: data <= 19'h00492; 
        10'b0001100100: data <= 19'h0032b; 
        10'b0001100101: data <= 19'h00393; 
        10'b0001100110: data <= 19'h002cb; 
        10'b0001100111: data <= 19'h00036; 
        10'b0001101000: data <= 19'h7ffb9; 
        10'b0001101001: data <= 19'h7fc97; 
        10'b0001101010: data <= 19'h7fe07; 
        10'b0001101011: data <= 19'h7ffd4; 
        10'b0001101100: data <= 19'h00018; 
        10'b0001101101: data <= 19'h7fe81; 
        10'b0001101110: data <= 19'h7ff52; 
        10'b0001101111: data <= 19'h7feb0; 
        10'b0001110000: data <= 19'h7ff4c; 
        10'b0001110001: data <= 19'h7ffe3; 
        10'b0001110010: data <= 19'h7ff78; 
        10'b0001110011: data <= 19'h0000f; 
        10'b0001110100: data <= 19'h000be; 
        10'b0001110101: data <= 19'h7fffe; 
        10'b0001110110: data <= 19'h002df; 
        10'b0001110111: data <= 19'h0026d; 
        10'b0001111000: data <= 19'h0069c; 
        10'b0001111001: data <= 19'h005ae; 
        10'b0001111010: data <= 19'h0070b; 
        10'b0001111011: data <= 19'h00879; 
        10'b0001111100: data <= 19'h009d4; 
        10'b0001111101: data <= 19'h00a88; 
        10'b0001111110: data <= 19'h00978; 
        10'b0001111111: data <= 19'h006f1; 
        10'b0010000000: data <= 19'h003ea; 
        10'b0010000001: data <= 19'h00322; 
        10'b0010000010: data <= 19'h0051f; 
        10'b0010000011: data <= 19'h000a1; 
        10'b0010000100: data <= 19'h7fc7f; 
        10'b0010000101: data <= 19'h7fa88; 
        10'b0010000110: data <= 19'h7fb54; 
        10'b0010000111: data <= 19'h7fb6d; 
        10'b0010001000: data <= 19'h7ff72; 
        10'b0010001001: data <= 19'h7ff2b; 
        10'b0010001010: data <= 19'h7fecf; 
        10'b0010001011: data <= 19'h7ffb0; 
        10'b0010001100: data <= 19'h7fe47; 
        10'b0010001101: data <= 19'h7fe07; 
        10'b0010001110: data <= 19'h7fe87; 
        10'b0010001111: data <= 19'h7fe87; 
        10'b0010010000: data <= 19'h0005e; 
        10'b0010010001: data <= 19'h002fd; 
        10'b0010010010: data <= 19'h00576; 
        10'b0010010011: data <= 19'h0045d; 
        10'b0010010100: data <= 19'h004fe; 
        10'b0010010101: data <= 19'h00468; 
        10'b0010010110: data <= 19'h003fd; 
        10'b0010010111: data <= 19'h00531; 
        10'b0010011000: data <= 19'h00545; 
        10'b0010011001: data <= 19'h00653; 
        10'b0010011010: data <= 19'h00115; 
        10'b0010011011: data <= 19'h00436; 
        10'b0010011100: data <= 19'h004dd; 
        10'b0010011101: data <= 19'h7ffa0; 
        10'b0010011110: data <= 19'h7ffbe; 
        10'b0010011111: data <= 19'h7fdcc; 
        10'b0010100000: data <= 19'h7fcef; 
        10'b0010100001: data <= 19'h7f97e; 
        10'b0010100010: data <= 19'h7f7ae; 
        10'b0010100011: data <= 19'h7f8f5; 
        10'b0010100100: data <= 19'h7fdf5; 
        10'b0010100101: data <= 19'h00002; 
        10'b0010100110: data <= 19'h7fe99; 
        10'b0010100111: data <= 19'h7ff23; 
        10'b0010101000: data <= 19'h7fe74; 
        10'b0010101001: data <= 19'h7fec9; 
        10'b0010101010: data <= 19'h7fea7; 
        10'b0010101011: data <= 19'h000a1; 
        10'b0010101100: data <= 19'h003b3; 
        10'b0010101101: data <= 19'h006e0; 
        10'b0010101110: data <= 19'h00542; 
        10'b0010101111: data <= 19'h00407; 
        10'b0010110000: data <= 19'h0061a; 
        10'b0010110001: data <= 19'h004fa; 
        10'b0010110010: data <= 19'h0046d; 
        10'b0010110011: data <= 19'h0043c; 
        10'b0010110100: data <= 19'h005a9; 
        10'b0010110101: data <= 19'h0081f; 
        10'b0010110110: data <= 19'h005a5; 
        10'b0010110111: data <= 19'h0020a; 
        10'b0010111000: data <= 19'h0055f; 
        10'b0010111001: data <= 19'h004ed; 
        10'b0010111010: data <= 19'h004b0; 
        10'b0010111011: data <= 19'h7fde7; 
        10'b0010111100: data <= 19'h00200; 
        10'b0010111101: data <= 19'h7fe04; 
        10'b0010111110: data <= 19'h7f8dc; 
        10'b0010111111: data <= 19'h7f8dc; 
        10'b0011000000: data <= 19'h7fba0; 
        10'b0011000001: data <= 19'h7ff1f; 
        10'b0011000010: data <= 19'h7ffce; 
        10'b0011000011: data <= 19'h7ff50; 
        10'b0011000100: data <= 19'h00016; 
        10'b0011000101: data <= 19'h7ffc2; 
        10'b0011000110: data <= 19'h0006b; 
        10'b0011000111: data <= 19'h00316; 
        10'b0011001000: data <= 19'h0081e; 
        10'b0011001001: data <= 19'h00813; 
        10'b0011001010: data <= 19'h005b1; 
        10'b0011001011: data <= 19'h00199; 
        10'b0011001100: data <= 19'h001b7; 
        10'b0011001101: data <= 19'h0039e; 
        10'b0011001110: data <= 19'h0011c; 
        10'b0011001111: data <= 19'h001a6; 
        10'b0011010000: data <= 19'h004c3; 
        10'b0011010001: data <= 19'h00482; 
        10'b0011010010: data <= 19'h00779; 
        10'b0011010011: data <= 19'h00464; 
        10'b0011010100: data <= 19'h00158; 
        10'b0011010101: data <= 19'h003c0; 
        10'b0011010110: data <= 19'h0031c; 
        10'b0011010111: data <= 19'h00361; 
        10'b0011011000: data <= 19'h0036c; 
        10'b0011011001: data <= 19'h0007c; 
        10'b0011011010: data <= 19'h7fc8d; 
        10'b0011011011: data <= 19'h7f7fc; 
        10'b0011011100: data <= 19'h7fa41; 
        10'b0011011101: data <= 19'h7fe7e; 
        10'b0011011110: data <= 19'h7fe09; 
        10'b0011011111: data <= 19'h7fef4; 
        10'b0011100000: data <= 19'h7ff3d; 
        10'b0011100001: data <= 19'h7fed3; 
        10'b0011100010: data <= 19'h00057; 
        10'b0011100011: data <= 19'h002e2; 
        10'b0011100100: data <= 19'h006b1; 
        10'b0011100101: data <= 19'h0065c; 
        10'b0011100110: data <= 19'h004c7; 
        10'b0011100111: data <= 19'h001f4; 
        10'b0011101000: data <= 19'h0033c; 
        10'b0011101001: data <= 19'h0018b; 
        10'b0011101010: data <= 19'h00416; 
        10'b0011101011: data <= 19'h00150; 
        10'b0011101100: data <= 19'h0011e; 
        10'b0011101101: data <= 19'h00200; 
        10'b0011101110: data <= 19'h00820; 
        10'b0011101111: data <= 19'h006be; 
        10'b0011110000: data <= 19'h0018e; 
        10'b0011110001: data <= 19'h003bf; 
        10'b0011110010: data <= 19'h00562; 
        10'b0011110011: data <= 19'h00382; 
        10'b0011110100: data <= 19'h00522; 
        10'b0011110101: data <= 19'h002a5; 
        10'b0011110110: data <= 19'h7fea0; 
        10'b0011110111: data <= 19'h7f893; 
        10'b0011111000: data <= 19'h7fa70; 
        10'b0011111001: data <= 19'h7fdf8; 
        10'b0011111010: data <= 19'h7fe46; 
        10'b0011111011: data <= 19'h7fec2; 
        10'b0011111100: data <= 19'h7ff07; 
        10'b0011111101: data <= 19'h7fe18; 
        10'b0011111110: data <= 19'h7ff64; 
        10'b0011111111: data <= 19'h0013e; 
        10'b0100000000: data <= 19'h00375; 
        10'b0100000001: data <= 19'h00496; 
        10'b0100000010: data <= 19'h003cd; 
        10'b0100000011: data <= 19'h000ec; 
        10'b0100000100: data <= 19'h7ff85; 
        10'b0100000101: data <= 19'h7fc75; 
        10'b0100000110: data <= 19'h7f93f; 
        10'b0100000111: data <= 19'h7f398; 
        10'b0100001000: data <= 19'h7f5ef; 
        10'b0100001001: data <= 19'h7fea9; 
        10'b0100001010: data <= 19'h009ad; 
        10'b0100001011: data <= 19'h00ee0; 
        10'b0100001100: data <= 19'h00898; 
        10'b0100001101: data <= 19'h00506; 
        10'b0100001110: data <= 19'h00576; 
        10'b0100001111: data <= 19'h0050c; 
        10'b0100010000: data <= 19'h00790; 
        10'b0100010001: data <= 19'h004d3; 
        10'b0100010010: data <= 19'h7fe8a; 
        10'b0100010011: data <= 19'h7f8a0; 
        10'b0100010100: data <= 19'h7fc4a; 
        10'b0100010101: data <= 19'h7fde8; 
        10'b0100010110: data <= 19'h7fe6d; 
        10'b0100010111: data <= 19'h7feb0; 
        10'b0100011000: data <= 19'h7ffca; 
        10'b0100011001: data <= 19'h7ffaf; 
        10'b0100011010: data <= 19'h0001a; 
        10'b0100011011: data <= 19'h001dd; 
        10'b0100011100: data <= 19'h001ad; 
        10'b0100011101: data <= 19'h000b7; 
        10'b0100011110: data <= 19'h7fdd6; 
        10'b0100011111: data <= 19'h7fa86; 
        10'b0100100000: data <= 19'h7f5fb; 
        10'b0100100001: data <= 19'h7f1ad; 
        10'b0100100010: data <= 19'h7ee73; 
        10'b0100100011: data <= 19'h7ee00; 
        10'b0100100100: data <= 19'h7f2bd; 
        10'b0100100101: data <= 19'h7fca7; 
        10'b0100100110: data <= 19'h007ef; 
        10'b0100100111: data <= 19'h0092c; 
        10'b0100101000: data <= 19'h007cf; 
        10'b0100101001: data <= 19'h00748; 
        10'b0100101010: data <= 19'h0047e; 
        10'b0100101011: data <= 19'h007cc; 
        10'b0100101100: data <= 19'h0073c; 
        10'b0100101101: data <= 19'h002e6; 
        10'b0100101110: data <= 19'h7fd68; 
        10'b0100101111: data <= 19'h7fb37; 
        10'b0100110000: data <= 19'h7fe36; 
        10'b0100110001: data <= 19'h7fdf9; 
        10'b0100110010: data <= 19'h7ff24; 
        10'b0100110011: data <= 19'h7ffc8; 
        10'b0100110100: data <= 19'h0003c; 
        10'b0100110101: data <= 19'h7ffc8; 
        10'b0100110110: data <= 19'h7fe58; 
        10'b0100110111: data <= 19'h001d1; 
        10'b0100111000: data <= 19'h7feed; 
        10'b0100111001: data <= 19'h7fa62; 
        10'b0100111010: data <= 19'h7f793; 
        10'b0100111011: data <= 19'h7f39e; 
        10'b0100111100: data <= 19'h7f085; 
        10'b0100111101: data <= 19'h7f29f; 
        10'b0100111110: data <= 19'h7f5d0; 
        10'b0100111111: data <= 19'h7fb33; 
        10'b0101000000: data <= 19'h7fd66; 
        10'b0101000001: data <= 19'h0035d; 
        10'b0101000010: data <= 19'h00548; 
        10'b0101000011: data <= 19'h0054f; 
        10'b0101000100: data <= 19'h0026c; 
        10'b0101000101: data <= 19'h0057f; 
        10'b0101000110: data <= 19'h006cd; 
        10'b0101000111: data <= 19'h006a2; 
        10'b0101001000: data <= 19'h005ca; 
        10'b0101001001: data <= 19'h00007; 
        10'b0101001010: data <= 19'h7fd73; 
        10'b0101001011: data <= 19'h7fdde; 
        10'b0101001100: data <= 19'h7fe1f; 
        10'b0101001101: data <= 19'h7fee3; 
        10'b0101001110: data <= 19'h7fe76; 
        10'b0101001111: data <= 19'h7fe46; 
        10'b0101010000: data <= 19'h00011; 
        10'b0101010001: data <= 19'h7feb3; 
        10'b0101010010: data <= 19'h7ffab; 
        10'b0101010011: data <= 19'h7ffe6; 
        10'b0101010100: data <= 19'h7fdf5; 
        10'b0101010101: data <= 19'h7fa5d; 
        10'b0101010110: data <= 19'h7f621; 
        10'b0101010111: data <= 19'h7f3a7; 
        10'b0101011000: data <= 19'h7f4d6; 
        10'b0101011001: data <= 19'h7fa0e; 
        10'b0101011010: data <= 19'h0001e; 
        10'b0101011011: data <= 19'h000fe; 
        10'b0101011100: data <= 19'h00192; 
        10'b0101011101: data <= 19'h00391; 
        10'b0101011110: data <= 19'h008d6; 
        10'b0101011111: data <= 19'h00491; 
        10'b0101100000: data <= 19'h0031e; 
        10'b0101100001: data <= 19'h0046a; 
        10'b0101100010: data <= 19'h00389; 
        10'b0101100011: data <= 19'h7ffb1; 
        10'b0101100100: data <= 19'h7fb6d; 
        10'b0101100101: data <= 19'h7f9b8; 
        10'b0101100110: data <= 19'h7f96c; 
        10'b0101100111: data <= 19'h7fbd1; 
        10'b0101101000: data <= 19'h7ff44; 
        10'b0101101001: data <= 19'h7febc; 
        10'b0101101010: data <= 19'h7ff51; 
        10'b0101101011: data <= 19'h7ff85; 
        10'b0101101100: data <= 19'h7ff1c; 
        10'b0101101101: data <= 19'h7fea6; 
        10'b0101101110: data <= 19'h7ff2b; 
        10'b0101101111: data <= 19'h7ff72; 
        10'b0101110000: data <= 19'h7fd63; 
        10'b0101110001: data <= 19'h7fc25; 
        10'b0101110010: data <= 19'h7f7f9; 
        10'b0101110011: data <= 19'h7f6bc; 
        10'b0101110100: data <= 19'h7f9b7; 
        10'b0101110101: data <= 19'h7fec3; 
        10'b0101110110: data <= 19'h7fdf5; 
        10'b0101110111: data <= 19'h7faac; 
        10'b0101111000: data <= 19'h0006d; 
        10'b0101111001: data <= 19'h0079b; 
        10'b0101111010: data <= 19'h007af; 
        10'b0101111011: data <= 19'h00167; 
        10'b0101111100: data <= 19'h0037d; 
        10'b0101111101: data <= 19'h003b8; 
        10'b0101111110: data <= 19'h001f9; 
        10'b0101111111: data <= 19'h7fd62; 
        10'b0110000000: data <= 19'h7f8fd; 
        10'b0110000001: data <= 19'h7f8f4; 
        10'b0110000010: data <= 19'h7fa6f; 
        10'b0110000011: data <= 19'h7fc17; 
        10'b0110000100: data <= 19'h7fdc1; 
        10'b0110000101: data <= 19'h7fff4; 
        10'b0110000110: data <= 19'h7ff97; 
        10'b0110000111: data <= 19'h7fece; 
        10'b0110001000: data <= 19'h0002f; 
        10'b0110001001: data <= 19'h7fe79; 
        10'b0110001010: data <= 19'h7ff06; 
        10'b0110001011: data <= 19'h7ff5d; 
        10'b0110001100: data <= 19'h7ff84; 
        10'b0110001101: data <= 19'h7fcc7; 
        10'b0110001110: data <= 19'h7f8c2; 
        10'b0110001111: data <= 19'h7f974; 
        10'b0110010000: data <= 19'h7fb8e; 
        10'b0110010001: data <= 19'h7ff62; 
        10'b0110010010: data <= 19'h7fb56; 
        10'b0110010011: data <= 19'h7fb07; 
        10'b0110010100: data <= 19'h00169; 
        10'b0110010101: data <= 19'h003ae; 
        10'b0110010110: data <= 19'h003ee; 
        10'b0110010111: data <= 19'h7ff6a; 
        10'b0110011000: data <= 19'h7fe67; 
        10'b0110011001: data <= 19'h7fed0; 
        10'b0110011010: data <= 19'h00089; 
        10'b0110011011: data <= 19'h7fcf3; 
        10'b0110011100: data <= 19'h7fbdf; 
        10'b0110011101: data <= 19'h7fe00; 
        10'b0110011110: data <= 19'h7fd29; 
        10'b0110011111: data <= 19'h7fe15; 
        10'b0110100000: data <= 19'h7fd7a; 
        10'b0110100001: data <= 19'h7fdbb; 
        10'b0110100010: data <= 19'h0000f; 
        10'b0110100011: data <= 19'h0001d; 
        10'b0110100100: data <= 19'h0002b; 
        10'b0110100101: data <= 19'h7fe7f; 
        10'b0110100110: data <= 19'h0003a; 
        10'b0110100111: data <= 19'h0008e; 
        10'b0110101000: data <= 19'h7ff5a; 
        10'b0110101001: data <= 19'h7fc61; 
        10'b0110101010: data <= 19'h7f948; 
        10'b0110101011: data <= 19'h7f8cf; 
        10'b0110101100: data <= 19'h7fa9f; 
        10'b0110101101: data <= 19'h7fcd9; 
        10'b0110101110: data <= 19'h7fc82; 
        10'b0110101111: data <= 19'h7fed2; 
        10'b0110110000: data <= 19'h00174; 
        10'b0110110001: data <= 19'h005fc; 
        10'b0110110010: data <= 19'h0036f; 
        10'b0110110011: data <= 19'h7ffa9; 
        10'b0110110100: data <= 19'h7fb01; 
        10'b0110110101: data <= 19'h7fe8d; 
        10'b0110110110: data <= 19'h7ff82; 
        10'b0110110111: data <= 19'h00150; 
        10'b0110111000: data <= 19'h0031a; 
        10'b0110111001: data <= 19'h00307; 
        10'b0110111010: data <= 19'h0010c; 
        10'b0110111011: data <= 19'h00066; 
        10'b0110111100: data <= 19'h7fe1b; 
        10'b0110111101: data <= 19'h7ff93; 
        10'b0110111110: data <= 19'h7ff66; 
        10'b0110111111: data <= 19'h7fe7e; 
        10'b0111000000: data <= 19'h7ff6f; 
        10'b0111000001: data <= 19'h7ffae; 
        10'b0111000010: data <= 19'h00161; 
        10'b0111000011: data <= 19'h0003f; 
        10'b0111000100: data <= 19'h00103; 
        10'b0111000101: data <= 19'h7fe54; 
        10'b0111000110: data <= 19'h7fd41; 
        10'b0111000111: data <= 19'h7fb3f; 
        10'b0111001000: data <= 19'h7f5a8; 
        10'b0111001001: data <= 19'h7f519; 
        10'b0111001010: data <= 19'h7f657; 
        10'b0111001011: data <= 19'h7fd8e; 
        10'b0111001100: data <= 19'h002e2; 
        10'b0111001101: data <= 19'h00776; 
        10'b0111001110: data <= 19'h7ff31; 
        10'b0111001111: data <= 19'h7fa8e; 
        10'b0111010000: data <= 19'h7fa3d; 
        10'b0111010001: data <= 19'h7fe20; 
        10'b0111010010: data <= 19'h0026e; 
        10'b0111010011: data <= 19'h0065d; 
        10'b0111010100: data <= 19'h0047b; 
        10'b0111010101: data <= 19'h005a3; 
        10'b0111010110: data <= 19'h0057a; 
        10'b0111010111: data <= 19'h0026d; 
        10'b0111011000: data <= 19'h7ff48; 
        10'b0111011001: data <= 19'h7ff84; 
        10'b0111011010: data <= 19'h7ffef; 
        10'b0111011011: data <= 19'h7ffd2; 
        10'b0111011100: data <= 19'h7ffc7; 
        10'b0111011101: data <= 19'h0003c; 
        10'b0111011110: data <= 19'h00008; 
        10'b0111011111: data <= 19'h0037d; 
        10'b0111100000: data <= 19'h001ed; 
        10'b0111100001: data <= 19'h0009a; 
        10'b0111100010: data <= 19'h7fe27; 
        10'b0111100011: data <= 19'h7f9b9; 
        10'b0111100100: data <= 19'h7f4d3; 
        10'b0111100101: data <= 19'h7ee47; 
        10'b0111100110: data <= 19'h7e9f1; 
        10'b0111100111: data <= 19'h7ebde; 
        10'b0111101000: data <= 19'h7f0b7; 
        10'b0111101001: data <= 19'h7f74b; 
        10'b0111101010: data <= 19'h7f7eb; 
        10'b0111101011: data <= 19'h7f8c9; 
        10'b0111101100: data <= 19'h7ffb7; 
        10'b0111101101: data <= 19'h0023a; 
        10'b0111101110: data <= 19'h00414; 
        10'b0111101111: data <= 19'h00675; 
        10'b0111110000: data <= 19'h00156; 
        10'b0111110001: data <= 19'h007d0; 
        10'b0111110010: data <= 19'h007cc; 
        10'b0111110011: data <= 19'h00259; 
        10'b0111110100: data <= 19'h7fed9; 
        10'b0111110101: data <= 19'h7fe57; 
        10'b0111110110: data <= 19'h7fe7c; 
        10'b0111110111: data <= 19'h7fe9e; 
        10'b0111111000: data <= 19'h7ff25; 
        10'b0111111001: data <= 19'h7ff33; 
        10'b0111111010: data <= 19'h000ad; 
        10'b0111111011: data <= 19'h00529; 
        10'b0111111100: data <= 19'h003b7; 
        10'b0111111101: data <= 19'h0023e; 
        10'b0111111110: data <= 19'h0012d; 
        10'b0111111111: data <= 19'h7fea3; 
        10'b1000000000: data <= 19'h7fc07; 
        10'b1000000001: data <= 19'h7f306; 
        10'b1000000010: data <= 19'h7ece4; 
        10'b1000000011: data <= 19'h7edeb; 
        10'b1000000100: data <= 19'h7ea2b; 
        10'b1000000101: data <= 19'h7ee2e; 
        10'b1000000110: data <= 19'h7f4ba; 
        10'b1000000111: data <= 19'h7fd70; 
        10'b1000001000: data <= 19'h0048d; 
        10'b1000001001: data <= 19'h00622; 
        10'b1000001010: data <= 19'h0069c; 
        10'b1000001011: data <= 19'h00689; 
        10'b1000001100: data <= 19'h00494; 
        10'b1000001101: data <= 19'h0091f; 
        10'b1000001110: data <= 19'h00883; 
        10'b1000001111: data <= 19'h00341; 
        10'b1000010000: data <= 19'h7fd01; 
        10'b1000010001: data <= 19'h7fdf9; 
        10'b1000010010: data <= 19'h7fe86; 
        10'b1000010011: data <= 19'h7ffc4; 
        10'b1000010100: data <= 19'h7ffc4; 
        10'b1000010101: data <= 19'h7fe82; 
        10'b1000010110: data <= 19'h7ff0b; 
        10'b1000010111: data <= 19'h00678; 
        10'b1000011000: data <= 19'h00699; 
        10'b1000011001: data <= 19'h007c0; 
        10'b1000011010: data <= 19'h006ae; 
        10'b1000011011: data <= 19'h00274; 
        10'b1000011100: data <= 19'h000bc; 
        10'b1000011101: data <= 19'h7fd47; 
        10'b1000011110: data <= 19'h7fe09; 
        10'b1000011111: data <= 19'h7f9d7; 
        10'b1000100000: data <= 19'h7f700; 
        10'b1000100001: data <= 19'h7f66e; 
        10'b1000100010: data <= 19'h7f97a; 
        10'b1000100011: data <= 19'h0024c; 
        10'b1000100100: data <= 19'h00629; 
        10'b1000100101: data <= 19'h007b3; 
        10'b1000100110: data <= 19'h008a1; 
        10'b1000100111: data <= 19'h007b8; 
        10'b1000101000: data <= 19'h006d5; 
        10'b1000101001: data <= 19'h007f8; 
        10'b1000101010: data <= 19'h0030e; 
        10'b1000101011: data <= 19'h0005b; 
        10'b1000101100: data <= 19'h7fd77; 
        10'b1000101101: data <= 19'h7ff88; 
        10'b1000101110: data <= 19'h7ffbf; 
        10'b1000101111: data <= 19'h7ff75; 
        10'b1000110000: data <= 19'h7ffac; 
        10'b1000110001: data <= 19'h7fe08; 
        10'b1000110010: data <= 19'h0012a; 
        10'b1000110011: data <= 19'h006f1; 
        10'b1000110100: data <= 19'h00888; 
        10'b1000110101: data <= 19'h0093c; 
        10'b1000110110: data <= 19'h009c8; 
        10'b1000110111: data <= 19'h004ef; 
        10'b1000111000: data <= 19'h005cf; 
        10'b1000111001: data <= 19'h00692; 
        10'b1000111010: data <= 19'h0026d; 
        10'b1000111011: data <= 19'h7ff57; 
        10'b1000111100: data <= 19'h7fdcb; 
        10'b1000111101: data <= 19'h7fc9f; 
        10'b1000111110: data <= 19'h00106; 
        10'b1000111111: data <= 19'h001d2; 
        10'b1001000000: data <= 19'h00379; 
        10'b1001000001: data <= 19'h00631; 
        10'b1001000010: data <= 19'h0067c; 
        10'b1001000011: data <= 19'h0046a; 
        10'b1001000100: data <= 19'h007af; 
        10'b1001000101: data <= 19'h0045e; 
        10'b1001000110: data <= 19'h7ff30; 
        10'b1001000111: data <= 19'h7fe40; 
        10'b1001001000: data <= 19'h7fdf8; 
        10'b1001001001: data <= 19'h7ff67; 
        10'b1001001010: data <= 19'h7ff60; 
        10'b1001001011: data <= 19'h7ff4d; 
        10'b1001001100: data <= 19'h7fead; 
        10'b1001001101: data <= 19'h7ffe9; 
        10'b1001001110: data <= 19'h7ff85; 
        10'b1001001111: data <= 19'h00374; 
        10'b1001010000: data <= 19'h0083d; 
        10'b1001010001: data <= 19'h0083a; 
        10'b1001010010: data <= 19'h00730; 
        10'b1001010011: data <= 19'h0040e; 
        10'b1001010100: data <= 19'h00453; 
        10'b1001010101: data <= 19'h0016e; 
        10'b1001010110: data <= 19'h7ff6e; 
        10'b1001010111: data <= 19'h7fe0e; 
        10'b1001011000: data <= 19'h000a0; 
        10'b1001011001: data <= 19'h7ffa6; 
        10'b1001011010: data <= 19'h7ff7e; 
        10'b1001011011: data <= 19'h7ff0d; 
        10'b1001011100: data <= 19'h00204; 
        10'b1001011101: data <= 19'h000bd; 
        10'b1001011110: data <= 19'h003f5; 
        10'b1001011111: data <= 19'h0065d; 
        10'b1001100000: data <= 19'h003b3; 
        10'b1001100001: data <= 19'h0016a; 
        10'b1001100010: data <= 19'h7fe91; 
        10'b1001100011: data <= 19'h7fc4e; 
        10'b1001100100: data <= 19'h7fecc; 
        10'b1001100101: data <= 19'h7fe7a; 
        10'b1001100110: data <= 19'h7fdfe; 
        10'b1001100111: data <= 19'h7fe1e; 
        10'b1001101000: data <= 19'h7ff2c; 
        10'b1001101001: data <= 19'h7ff6c; 
        10'b1001101010: data <= 19'h7ff9e; 
        10'b1001101011: data <= 19'h00225; 
        10'b1001101100: data <= 19'h00423; 
        10'b1001101101: data <= 19'h005a2; 
        10'b1001101110: data <= 19'h00506; 
        10'b1001101111: data <= 19'h002dc; 
        10'b1001110000: data <= 19'h00039; 
        10'b1001110001: data <= 19'h00212; 
        10'b1001110010: data <= 19'h00280; 
        10'b1001110011: data <= 19'h0030a; 
        10'b1001110100: data <= 19'h000d7; 
        10'b1001110101: data <= 19'h7fee5; 
        10'b1001110110: data <= 19'h7fed2; 
        10'b1001110111: data <= 19'h7fe53; 
        10'b1001111000: data <= 19'h0014f; 
        10'b1001111001: data <= 19'h00100; 
        10'b1001111010: data <= 19'h000fc; 
        10'b1001111011: data <= 19'h00466; 
        10'b1001111100: data <= 19'h00222; 
        10'b1001111101: data <= 19'h7ff3e; 
        10'b1001111110: data <= 19'h7ff04; 
        10'b1001111111: data <= 19'h7feb7; 
        10'b1010000000: data <= 19'h7fd2c; 
        10'b1010000001: data <= 19'h7fde2; 
        10'b1010000010: data <= 19'h7ff9e; 
        10'b1010000011: data <= 19'h7fff1; 
        10'b1010000100: data <= 19'h7ff69; 
        10'b1010000101: data <= 19'h7fe6a; 
        10'b1010000110: data <= 19'h7feaf; 
        10'b1010000111: data <= 19'h0016a; 
        10'b1010001000: data <= 19'h00485; 
        10'b1010001001: data <= 19'h006d3; 
        10'b1010001010: data <= 19'h00516; 
        10'b1010001011: data <= 19'h0055f; 
        10'b1010001100: data <= 19'h0014d; 
        10'b1010001101: data <= 19'h00370; 
        10'b1010001110: data <= 19'h0022f; 
        10'b1010001111: data <= 19'h7fff7; 
        10'b1010010000: data <= 19'h7fe47; 
        10'b1010010001: data <= 19'h00047; 
        10'b1010010010: data <= 19'h000b3; 
        10'b1010010011: data <= 19'h001b8; 
        10'b1010010100: data <= 19'h00148; 
        10'b1010010101: data <= 19'h002a9; 
        10'b1010010110: data <= 19'h0043b; 
        10'b1010010111: data <= 19'h7ff49; 
        10'b1010011000: data <= 19'h7fd2b; 
        10'b1010011001: data <= 19'h7fd33; 
        10'b1010011010: data <= 19'h7fe86; 
        10'b1010011011: data <= 19'h7fe27; 
        10'b1010011100: data <= 19'h7ffd6; 
        10'b1010011101: data <= 19'h7ff86; 
        10'b1010011110: data <= 19'h7fe3e; 
        10'b1010011111: data <= 19'h7fe65; 
        10'b1010100000: data <= 19'h7febc; 
        10'b1010100001: data <= 19'h00033; 
        10'b1010100010: data <= 19'h00036; 
        10'b1010100011: data <= 19'h00007; 
        10'b1010100100: data <= 19'h002e8; 
        10'b1010100101: data <= 19'h004ae; 
        10'b1010100110: data <= 19'h00583; 
        10'b1010100111: data <= 19'h00681; 
        10'b1010101000: data <= 19'h0069b; 
        10'b1010101001: data <= 19'h0056b; 
        10'b1010101010: data <= 19'h007e6; 
        10'b1010101011: data <= 19'h00857; 
        10'b1010101100: data <= 19'h0088b; 
        10'b1010101101: data <= 19'h006ba; 
        10'b1010101110: data <= 19'h005ef; 
        10'b1010101111: data <= 19'h00463; 
        10'b1010110000: data <= 19'h00430; 
        10'b1010110001: data <= 19'h7ffa3; 
        10'b1010110010: data <= 19'h7fc98; 
        10'b1010110011: data <= 19'h7fb4a; 
        10'b1010110100: data <= 19'h7fbc4; 
        10'b1010110101: data <= 19'h7fd6b; 
        10'b1010110110: data <= 19'h7fd96; 
        10'b1010110111: data <= 19'h7ff49; 
        10'b1010111000: data <= 19'h7fecd; 
        10'b1010111001: data <= 19'h7fff8; 
        10'b1010111010: data <= 19'h7fec6; 
        10'b1010111011: data <= 19'h00039; 
        10'b1010111100: data <= 19'h7ffd0; 
        10'b1010111101: data <= 19'h7fdf9; 
        10'b1010111110: data <= 19'h00028; 
        10'b1010111111: data <= 19'h00054; 
        10'b1011000000: data <= 19'h7ff80; 
        10'b1011000001: data <= 19'h001d3; 
        10'b1011000010: data <= 19'h002bf; 
        10'b1011000011: data <= 19'h00189; 
        10'b1011000100: data <= 19'h003b4; 
        10'b1011000101: data <= 19'h003be; 
        10'b1011000110: data <= 19'h00700; 
        10'b1011000111: data <= 19'h00800; 
        10'b1011001000: data <= 19'h00897; 
        10'b1011001001: data <= 19'h006b9; 
        10'b1011001010: data <= 19'h004c8; 
        10'b1011001011: data <= 19'h001ec; 
        10'b1011001100: data <= 19'h7ff3a; 
        10'b1011001101: data <= 19'h7fcf8; 
        10'b1011001110: data <= 19'h7fcf4; 
        10'b1011001111: data <= 19'h7fd81; 
        10'b1011010000: data <= 19'h7fd86; 
        10'b1011010001: data <= 19'h7fec1; 
        10'b1011010010: data <= 19'h7fec1; 
        10'b1011010011: data <= 19'h7ffdd; 
        10'b1011010100: data <= 19'h7fe7c; 
        10'b1011010101: data <= 19'h00031; 
        10'b1011010110: data <= 19'h7fe04; 
        10'b1011010111: data <= 19'h7ffb9; 
        10'b1011011000: data <= 19'h7fe90; 
        10'b1011011001: data <= 19'h7fdf4; 
        10'b1011011010: data <= 19'h7fe0c; 
        10'b1011011011: data <= 19'h7ff80; 
        10'b1011011100: data <= 19'h7ff87; 
        10'b1011011101: data <= 19'h7fea7; 
        10'b1011011110: data <= 19'h7fe6e; 
        10'b1011011111: data <= 19'h7ff75; 
        10'b1011100000: data <= 19'h7ff80; 
        10'b1011100001: data <= 19'h7ff58; 
        10'b1011100010: data <= 19'h7ff15; 
        10'b1011100011: data <= 19'h7ff3c; 
        10'b1011100100: data <= 19'h7fedd; 
        10'b1011100101: data <= 19'h7ff63; 
        10'b1011100110: data <= 19'h7fedb; 
        10'b1011100111: data <= 19'h7fdca; 
        10'b1011101000: data <= 19'h7fea5; 
        10'b1011101001: data <= 19'h7ff5b; 
        10'b1011101010: data <= 19'h7ff1c; 
        10'b1011101011: data <= 19'h7ff6c; 
        10'b1011101100: data <= 19'h7fe17; 
        10'b1011101101: data <= 19'h7fe1f; 
        10'b1011101110: data <= 19'h7ffb7; 
        10'b1011101111: data <= 19'h7fee8; 
        10'b1011110000: data <= 19'h0000d; 
        10'b1011110001: data <= 19'h7fe88; 
        10'b1011110010: data <= 19'h7ffd7; 
        10'b1011110011: data <= 19'h0003a; 
        10'b1011110100: data <= 19'h7ff06; 
        10'b1011110101: data <= 19'h7fe79; 
        10'b1011110110: data <= 19'h7ff53; 
        10'b1011110111: data <= 19'h7fe15; 
        10'b1011111000: data <= 19'h00019; 
        10'b1011111001: data <= 19'h7ff7a; 
        10'b1011111010: data <= 19'h7ffe7; 
        10'b1011111011: data <= 19'h7ff64; 
        10'b1011111100: data <= 19'h7ffb0; 
        10'b1011111101: data <= 19'h7fe0f; 
        10'b1011111110: data <= 19'h7fe69; 
        10'b1011111111: data <= 19'h7ff95; 
        10'b1100000000: data <= 19'h7fe66; 
        10'b1100000001: data <= 19'h7ffb3; 
        10'b1100000010: data <= 19'h7fece; 
        10'b1100000011: data <= 19'h7ff4c; 
        10'b1100000100: data <= 19'h7fedc; 
        10'b1100000101: data <= 19'h7fff6; 
        10'b1100000110: data <= 19'h7fe2a; 
        10'b1100000111: data <= 19'h7fe7c; 
        10'b1100001000: data <= 19'h7ffdf; 
        10'b1100001001: data <= 19'h7ff56; 
        10'b1100001010: data <= 19'h7fe78; 
        10'b1100001011: data <= 19'h7ff86; 
        10'b1100001100: data <= 19'h7fe31; 
        10'b1100001101: data <= 19'h7fe0a; 
        10'b1100001110: data <= 19'h7ffe3; 
        10'b1100001111: data <= 19'h7ff16; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 14) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 20'hffebd; 
        10'b0000000001: data <= 20'hffce3; 
        10'b0000000010: data <= 20'hfffd9; 
        10'b0000000011: data <= 20'h00024; 
        10'b0000000100: data <= 20'h00050; 
        10'b0000000101: data <= 20'hfffba; 
        10'b0000000110: data <= 20'hffed1; 
        10'b0000000111: data <= 20'h00053; 
        10'b0000001000: data <= 20'hffd7c; 
        10'b0000001001: data <= 20'h00033; 
        10'b0000001010: data <= 20'h00036; 
        10'b0000001011: data <= 20'hffddb; 
        10'b0000001100: data <= 20'hffdce; 
        10'b0000001101: data <= 20'hffdc0; 
        10'b0000001110: data <= 20'hffdeb; 
        10'b0000001111: data <= 20'hffe31; 
        10'b0000010000: data <= 20'h0000b; 
        10'b0000010001: data <= 20'h00023; 
        10'b0000010010: data <= 20'hffce4; 
        10'b0000010011: data <= 20'h00051; 
        10'b0000010100: data <= 20'hffefd; 
        10'b0000010101: data <= 20'hfff20; 
        10'b0000010110: data <= 20'hffbeb; 
        10'b0000010111: data <= 20'hfffc6; 
        10'b0000011000: data <= 20'hfffd9; 
        10'b0000011001: data <= 20'hffc29; 
        10'b0000011010: data <= 20'hffe1c; 
        10'b0000011011: data <= 20'h0001d; 
        10'b0000011100: data <= 20'hffcca; 
        10'b0000011101: data <= 20'hffdfd; 
        10'b0000011110: data <= 20'hffcd7; 
        10'b0000011111: data <= 20'hffee7; 
        10'b0000100000: data <= 20'hffc60; 
        10'b0000100001: data <= 20'hffe44; 
        10'b0000100010: data <= 20'h0006a; 
        10'b0000100011: data <= 20'h0003b; 
        10'b0000100100: data <= 20'hffc24; 
        10'b0000100101: data <= 20'hffbf6; 
        10'b0000100110: data <= 20'hffc5f; 
        10'b0000100111: data <= 20'hffecf; 
        10'b0000101000: data <= 20'hfff24; 
        10'b0000101001: data <= 20'hffe27; 
        10'b0000101010: data <= 20'hffdd8; 
        10'b0000101011: data <= 20'hffd19; 
        10'b0000101100: data <= 20'h00066; 
        10'b0000101101: data <= 20'hffce6; 
        10'b0000101110: data <= 20'hfff50; 
        10'b0000101111: data <= 20'hffda3; 
        10'b0000110000: data <= 20'hffdaf; 
        10'b0000110001: data <= 20'hffc3f; 
        10'b0000110010: data <= 20'hffe6f; 
        10'b0000110011: data <= 20'hfffa1; 
        10'b0000110100: data <= 20'hffc9c; 
        10'b0000110101: data <= 20'hfffce; 
        10'b0000110110: data <= 20'hffea9; 
        10'b0000110111: data <= 20'hffca4; 
        10'b0000111000: data <= 20'hffd2d; 
        10'b0000111001: data <= 20'hffe6a; 
        10'b0000111010: data <= 20'hffe4f; 
        10'b0000111011: data <= 20'hffce7; 
        10'b0000111100: data <= 20'hfff03; 
        10'b0000111101: data <= 20'hfff56; 
        10'b0000111110: data <= 20'hffd5c; 
        10'b0000111111: data <= 20'hfff48; 
        10'b0001000000: data <= 20'hfffa7; 
        10'b0001000001: data <= 20'hffe27; 
        10'b0001000010: data <= 20'hffc8c; 
        10'b0001000011: data <= 20'hffca4; 
        10'b0001000100: data <= 20'hffc38; 
        10'b0001000101: data <= 20'hffcb8; 
        10'b0001000110: data <= 20'hffded; 
        10'b0001000111: data <= 20'hffda0; 
        10'b0001001000: data <= 20'hffd50; 
        10'b0001001001: data <= 20'hffd37; 
        10'b0001001010: data <= 20'hfff49; 
        10'b0001001011: data <= 20'hfffeb; 
        10'b0001001100: data <= 20'hffe12; 
        10'b0001001101: data <= 20'hffcd2; 
        10'b0001001110: data <= 20'h0005a; 
        10'b0001001111: data <= 20'hfffbd; 
        10'b0001010000: data <= 20'h00003; 
        10'b0001010001: data <= 20'hffd85; 
        10'b0001010010: data <= 20'hffc14; 
        10'b0001010011: data <= 20'hffe2d; 
        10'b0001010100: data <= 20'h0006f; 
        10'b0001010101: data <= 20'hfff40; 
        10'b0001010110: data <= 20'hffe3a; 
        10'b0001010111: data <= 20'hfff86; 
        10'b0001011000: data <= 20'hfff35; 
        10'b0001011001: data <= 20'h00004; 
        10'b0001011010: data <= 20'hffed4; 
        10'b0001011011: data <= 20'hfffc7; 
        10'b0001011100: data <= 20'hfff8c; 
        10'b0001011101: data <= 20'hffe81; 
        10'b0001011110: data <= 20'h00164; 
        10'b0001011111: data <= 20'h004a2; 
        10'b0001100000: data <= 20'h009c7; 
        10'b0001100001: data <= 20'h0081f; 
        10'b0001100010: data <= 20'h00848; 
        10'b0001100011: data <= 20'h00924; 
        10'b0001100100: data <= 20'h00656; 
        10'b0001100101: data <= 20'h00725; 
        10'b0001100110: data <= 20'h00595; 
        10'b0001100111: data <= 20'h0006b; 
        10'b0001101000: data <= 20'hfff72; 
        10'b0001101001: data <= 20'hff92e; 
        10'b0001101010: data <= 20'hffc0f; 
        10'b0001101011: data <= 20'hfffa9; 
        10'b0001101100: data <= 20'h00031; 
        10'b0001101101: data <= 20'hffd02; 
        10'b0001101110: data <= 20'hffea3; 
        10'b0001101111: data <= 20'hffd60; 
        10'b0001110000: data <= 20'hffe98; 
        10'b0001110001: data <= 20'hfffc6; 
        10'b0001110010: data <= 20'hffef0; 
        10'b0001110011: data <= 20'h0001e; 
        10'b0001110100: data <= 20'h0017c; 
        10'b0001110101: data <= 20'hffffd; 
        10'b0001110110: data <= 20'h005bf; 
        10'b0001110111: data <= 20'h004d9; 
        10'b0001111000: data <= 20'h00d39; 
        10'b0001111001: data <= 20'h00b5c; 
        10'b0001111010: data <= 20'h00e15; 
        10'b0001111011: data <= 20'h010f1; 
        10'b0001111100: data <= 20'h013a8; 
        10'b0001111101: data <= 20'h01511; 
        10'b0001111110: data <= 20'h012f1; 
        10'b0001111111: data <= 20'h00de3; 
        10'b0010000000: data <= 20'h007d5; 
        10'b0010000001: data <= 20'h00644; 
        10'b0010000010: data <= 20'h00a3d; 
        10'b0010000011: data <= 20'h00142; 
        10'b0010000100: data <= 20'hff8fd; 
        10'b0010000101: data <= 20'hff511; 
        10'b0010000110: data <= 20'hff6a8; 
        10'b0010000111: data <= 20'hff6db; 
        10'b0010001000: data <= 20'hffee3; 
        10'b0010001001: data <= 20'hffe56; 
        10'b0010001010: data <= 20'hffd9e; 
        10'b0010001011: data <= 20'hfff60; 
        10'b0010001100: data <= 20'hffc8d; 
        10'b0010001101: data <= 20'hffc0e; 
        10'b0010001110: data <= 20'hffd0d; 
        10'b0010001111: data <= 20'hffd0e; 
        10'b0010010000: data <= 20'h000bd; 
        10'b0010010001: data <= 20'h005f9; 
        10'b0010010010: data <= 20'h00aeb; 
        10'b0010010011: data <= 20'h008b9; 
        10'b0010010100: data <= 20'h009fc; 
        10'b0010010101: data <= 20'h008d0; 
        10'b0010010110: data <= 20'h007fa; 
        10'b0010010111: data <= 20'h00a62; 
        10'b0010011000: data <= 20'h00a8b; 
        10'b0010011001: data <= 20'h00ca5; 
        10'b0010011010: data <= 20'h00229; 
        10'b0010011011: data <= 20'h0086c; 
        10'b0010011100: data <= 20'h009ba; 
        10'b0010011101: data <= 20'hfff40; 
        10'b0010011110: data <= 20'hfff7b; 
        10'b0010011111: data <= 20'hffb97; 
        10'b0010100000: data <= 20'hff9df; 
        10'b0010100001: data <= 20'hff2fd; 
        10'b0010100010: data <= 20'hfef5c; 
        10'b0010100011: data <= 20'hff1ea; 
        10'b0010100100: data <= 20'hffbeb; 
        10'b0010100101: data <= 20'h00004; 
        10'b0010100110: data <= 20'hffd31; 
        10'b0010100111: data <= 20'hffe47; 
        10'b0010101000: data <= 20'hffce8; 
        10'b0010101001: data <= 20'hffd92; 
        10'b0010101010: data <= 20'hffd4e; 
        10'b0010101011: data <= 20'h00142; 
        10'b0010101100: data <= 20'h00765; 
        10'b0010101101: data <= 20'h00dc0; 
        10'b0010101110: data <= 20'h00a84; 
        10'b0010101111: data <= 20'h0080f; 
        10'b0010110000: data <= 20'h00c34; 
        10'b0010110001: data <= 20'h009f5; 
        10'b0010110010: data <= 20'h008d9; 
        10'b0010110011: data <= 20'h00877; 
        10'b0010110100: data <= 20'h00b52; 
        10'b0010110101: data <= 20'h0103e; 
        10'b0010110110: data <= 20'h00b4b; 
        10'b0010110111: data <= 20'h00414; 
        10'b0010111000: data <= 20'h00abf; 
        10'b0010111001: data <= 20'h009da; 
        10'b0010111010: data <= 20'h00960; 
        10'b0010111011: data <= 20'hffbce; 
        10'b0010111100: data <= 20'h00400; 
        10'b0010111101: data <= 20'hffc09; 
        10'b0010111110: data <= 20'hff1b8; 
        10'b0010111111: data <= 20'hff1b7; 
        10'b0011000000: data <= 20'hff741; 
        10'b0011000001: data <= 20'hffe3e; 
        10'b0011000010: data <= 20'hfff9c; 
        10'b0011000011: data <= 20'hffea0; 
        10'b0011000100: data <= 20'h0002b; 
        10'b0011000101: data <= 20'hfff84; 
        10'b0011000110: data <= 20'h000d7; 
        10'b0011000111: data <= 20'h0062c; 
        10'b0011001000: data <= 20'h0103c; 
        10'b0011001001: data <= 20'h01026; 
        10'b0011001010: data <= 20'h00b61; 
        10'b0011001011: data <= 20'h00333; 
        10'b0011001100: data <= 20'h0036e; 
        10'b0011001101: data <= 20'h0073c; 
        10'b0011001110: data <= 20'h00238; 
        10'b0011001111: data <= 20'h0034c; 
        10'b0011010000: data <= 20'h00986; 
        10'b0011010001: data <= 20'h00905; 
        10'b0011010010: data <= 20'h00ef2; 
        10'b0011010011: data <= 20'h008c8; 
        10'b0011010100: data <= 20'h002b1; 
        10'b0011010101: data <= 20'h00780; 
        10'b0011010110: data <= 20'h00638; 
        10'b0011010111: data <= 20'h006c1; 
        10'b0011011000: data <= 20'h006d9; 
        10'b0011011001: data <= 20'h000f8; 
        10'b0011011010: data <= 20'hff91b; 
        10'b0011011011: data <= 20'hfeff9; 
        10'b0011011100: data <= 20'hff482; 
        10'b0011011101: data <= 20'hffcfb; 
        10'b0011011110: data <= 20'hffc12; 
        10'b0011011111: data <= 20'hffde7; 
        10'b0011100000: data <= 20'hffe7a; 
        10'b0011100001: data <= 20'hffda5; 
        10'b0011100010: data <= 20'h000ae; 
        10'b0011100011: data <= 20'h005c4; 
        10'b0011100100: data <= 20'h00d62; 
        10'b0011100101: data <= 20'h00cb7; 
        10'b0011100110: data <= 20'h0098f; 
        10'b0011100111: data <= 20'h003e7; 
        10'b0011101000: data <= 20'h00679; 
        10'b0011101001: data <= 20'h00316; 
        10'b0011101010: data <= 20'h0082d; 
        10'b0011101011: data <= 20'h002a0; 
        10'b0011101100: data <= 20'h0023c; 
        10'b0011101101: data <= 20'h003ff; 
        10'b0011101110: data <= 20'h01040; 
        10'b0011101111: data <= 20'h00d7b; 
        10'b0011110000: data <= 20'h0031c; 
        10'b0011110001: data <= 20'h0077e; 
        10'b0011110010: data <= 20'h00ac4; 
        10'b0011110011: data <= 20'h00704; 
        10'b0011110100: data <= 20'h00a45; 
        10'b0011110101: data <= 20'h00549; 
        10'b0011110110: data <= 20'hffd40; 
        10'b0011110111: data <= 20'hff125; 
        10'b0011111000: data <= 20'hff4e1; 
        10'b0011111001: data <= 20'hffbf1; 
        10'b0011111010: data <= 20'hffc8c; 
        10'b0011111011: data <= 20'hffd85; 
        10'b0011111100: data <= 20'hffe0d; 
        10'b0011111101: data <= 20'hffc2f; 
        10'b0011111110: data <= 20'hffec8; 
        10'b0011111111: data <= 20'h0027c; 
        10'b0100000000: data <= 20'h006ea; 
        10'b0100000001: data <= 20'h0092d; 
        10'b0100000010: data <= 20'h00799; 
        10'b0100000011: data <= 20'h001d9; 
        10'b0100000100: data <= 20'hfff09; 
        10'b0100000101: data <= 20'hff8ea; 
        10'b0100000110: data <= 20'hff27d; 
        10'b0100000111: data <= 20'hfe731; 
        10'b0100001000: data <= 20'hfebde; 
        10'b0100001001: data <= 20'hffd52; 
        10'b0100001010: data <= 20'h0135b; 
        10'b0100001011: data <= 20'h01dc0; 
        10'b0100001100: data <= 20'h0112f; 
        10'b0100001101: data <= 20'h00a0d; 
        10'b0100001110: data <= 20'h00aec; 
        10'b0100001111: data <= 20'h00a19; 
        10'b0100010000: data <= 20'h00f1f; 
        10'b0100010001: data <= 20'h009a7; 
        10'b0100010010: data <= 20'hffd13; 
        10'b0100010011: data <= 20'hff13f; 
        10'b0100010100: data <= 20'hff893; 
        10'b0100010101: data <= 20'hffbd0; 
        10'b0100010110: data <= 20'hffcda; 
        10'b0100010111: data <= 20'hffd5f; 
        10'b0100011000: data <= 20'hfff94; 
        10'b0100011001: data <= 20'hfff5f; 
        10'b0100011010: data <= 20'h00035; 
        10'b0100011011: data <= 20'h003ba; 
        10'b0100011100: data <= 20'h0035a; 
        10'b0100011101: data <= 20'h0016d; 
        10'b0100011110: data <= 20'hffbad; 
        10'b0100011111: data <= 20'hff50b; 
        10'b0100100000: data <= 20'hfebf6; 
        10'b0100100001: data <= 20'hfe35b; 
        10'b0100100010: data <= 20'hfdce6; 
        10'b0100100011: data <= 20'hfdbff; 
        10'b0100100100: data <= 20'hfe57b; 
        10'b0100100101: data <= 20'hff94e; 
        10'b0100100110: data <= 20'h00fde; 
        10'b0100100111: data <= 20'h01258; 
        10'b0100101000: data <= 20'h00f9e; 
        10'b0100101001: data <= 20'h00e90; 
        10'b0100101010: data <= 20'h008fd; 
        10'b0100101011: data <= 20'h00f97; 
        10'b0100101100: data <= 20'h00e79; 
        10'b0100101101: data <= 20'h005cc; 
        10'b0100101110: data <= 20'hffad0; 
        10'b0100101111: data <= 20'hff66e; 
        10'b0100110000: data <= 20'hffc6c; 
        10'b0100110001: data <= 20'hffbf3; 
        10'b0100110010: data <= 20'hffe49; 
        10'b0100110011: data <= 20'hfff90; 
        10'b0100110100: data <= 20'h00079; 
        10'b0100110101: data <= 20'hfff91; 
        10'b0100110110: data <= 20'hffcaf; 
        10'b0100110111: data <= 20'h003a2; 
        10'b0100111000: data <= 20'hffdda; 
        10'b0100111001: data <= 20'hff4c4; 
        10'b0100111010: data <= 20'hfef27; 
        10'b0100111011: data <= 20'hfe73b; 
        10'b0100111100: data <= 20'hfe109; 
        10'b0100111101: data <= 20'hfe53e; 
        10'b0100111110: data <= 20'hfeba1; 
        10'b0100111111: data <= 20'hff665; 
        10'b0101000000: data <= 20'hffacc; 
        10'b0101000001: data <= 20'h006ba; 
        10'b0101000010: data <= 20'h00a90; 
        10'b0101000011: data <= 20'h00a9e; 
        10'b0101000100: data <= 20'h004d9; 
        10'b0101000101: data <= 20'h00aff; 
        10'b0101000110: data <= 20'h00d9b; 
        10'b0101000111: data <= 20'h00d44; 
        10'b0101001000: data <= 20'h00b95; 
        10'b0101001001: data <= 20'h0000e; 
        10'b0101001010: data <= 20'hffae7; 
        10'b0101001011: data <= 20'hffbbc; 
        10'b0101001100: data <= 20'hffc3e; 
        10'b0101001101: data <= 20'hffdc7; 
        10'b0101001110: data <= 20'hffceb; 
        10'b0101001111: data <= 20'hffc8d; 
        10'b0101010000: data <= 20'h00022; 
        10'b0101010001: data <= 20'hffd66; 
        10'b0101010010: data <= 20'hfff56; 
        10'b0101010011: data <= 20'hfffcc; 
        10'b0101010100: data <= 20'hffbeb; 
        10'b0101010101: data <= 20'hff4ba; 
        10'b0101010110: data <= 20'hfec43; 
        10'b0101010111: data <= 20'hfe74e; 
        10'b0101011000: data <= 20'hfe9ab; 
        10'b0101011001: data <= 20'hff41b; 
        10'b0101011010: data <= 20'h0003c; 
        10'b0101011011: data <= 20'h001fc; 
        10'b0101011100: data <= 20'h00325; 
        10'b0101011101: data <= 20'h00722; 
        10'b0101011110: data <= 20'h011ad; 
        10'b0101011111: data <= 20'h00922; 
        10'b0101100000: data <= 20'h0063d; 
        10'b0101100001: data <= 20'h008d3; 
        10'b0101100010: data <= 20'h00712; 
        10'b0101100011: data <= 20'hfff62; 
        10'b0101100100: data <= 20'hff6d9; 
        10'b0101100101: data <= 20'hff36f; 
        10'b0101100110: data <= 20'hff2d8; 
        10'b0101100111: data <= 20'hff7a3; 
        10'b0101101000: data <= 20'hffe88; 
        10'b0101101001: data <= 20'hffd77; 
        10'b0101101010: data <= 20'hffea2; 
        10'b0101101011: data <= 20'hfff0a; 
        10'b0101101100: data <= 20'hffe38; 
        10'b0101101101: data <= 20'hffd4c; 
        10'b0101101110: data <= 20'hffe57; 
        10'b0101101111: data <= 20'hffee4; 
        10'b0101110000: data <= 20'hffac7; 
        10'b0101110001: data <= 20'hff84b; 
        10'b0101110010: data <= 20'hfeff2; 
        10'b0101110011: data <= 20'hfed77; 
        10'b0101110100: data <= 20'hff36e; 
        10'b0101110101: data <= 20'hffd87; 
        10'b0101110110: data <= 20'hffbea; 
        10'b0101110111: data <= 20'hff558; 
        10'b0101111000: data <= 20'h000d9; 
        10'b0101111001: data <= 20'h00f37; 
        10'b0101111010: data <= 20'h00f5e; 
        10'b0101111011: data <= 20'h002ce; 
        10'b0101111100: data <= 20'h006fa; 
        10'b0101111101: data <= 20'h00770; 
        10'b0101111110: data <= 20'h003f2; 
        10'b0101111111: data <= 20'hffac4; 
        10'b0110000000: data <= 20'hff1f9; 
        10'b0110000001: data <= 20'hff1e8; 
        10'b0110000010: data <= 20'hff4de; 
        10'b0110000011: data <= 20'hff82e; 
        10'b0110000100: data <= 20'hffb82; 
        10'b0110000101: data <= 20'hfffe7; 
        10'b0110000110: data <= 20'hfff2e; 
        10'b0110000111: data <= 20'hffd9c; 
        10'b0110001000: data <= 20'h0005f; 
        10'b0110001001: data <= 20'hffcf3; 
        10'b0110001010: data <= 20'hffe0c; 
        10'b0110001011: data <= 20'hffebb; 
        10'b0110001100: data <= 20'hfff09; 
        10'b0110001101: data <= 20'hff98e; 
        10'b0110001110: data <= 20'hff183; 
        10'b0110001111: data <= 20'hff2e8; 
        10'b0110010000: data <= 20'hff71b; 
        10'b0110010001: data <= 20'hffec4; 
        10'b0110010010: data <= 20'hff6ad; 
        10'b0110010011: data <= 20'hff60f; 
        10'b0110010100: data <= 20'h002d1; 
        10'b0110010101: data <= 20'h0075d; 
        10'b0110010110: data <= 20'h007dc; 
        10'b0110010111: data <= 20'hffed5; 
        10'b0110011000: data <= 20'hffcce; 
        10'b0110011001: data <= 20'hffd9f; 
        10'b0110011010: data <= 20'h00113; 
        10'b0110011011: data <= 20'hff9e6; 
        10'b0110011100: data <= 20'hff7be; 
        10'b0110011101: data <= 20'hffc00; 
        10'b0110011110: data <= 20'hffa51; 
        10'b0110011111: data <= 20'hffc2a; 
        10'b0110100000: data <= 20'hffaf3; 
        10'b0110100001: data <= 20'hffb76; 
        10'b0110100010: data <= 20'h0001d; 
        10'b0110100011: data <= 20'h0003a; 
        10'b0110100100: data <= 20'h00055; 
        10'b0110100101: data <= 20'hffcff; 
        10'b0110100110: data <= 20'h00074; 
        10'b0110100111: data <= 20'h0011d; 
        10'b0110101000: data <= 20'hffeb4; 
        10'b0110101001: data <= 20'hff8c2; 
        10'b0110101010: data <= 20'hff28f; 
        10'b0110101011: data <= 20'hff19e; 
        10'b0110101100: data <= 20'hff53e; 
        10'b0110101101: data <= 20'hff9b1; 
        10'b0110101110: data <= 20'hff903; 
        10'b0110101111: data <= 20'hffda4; 
        10'b0110110000: data <= 20'h002e7; 
        10'b0110110001: data <= 20'h00bf7; 
        10'b0110110010: data <= 20'h006df; 
        10'b0110110011: data <= 20'hfff52; 
        10'b0110110100: data <= 20'hff603; 
        10'b0110110101: data <= 20'hffd1a; 
        10'b0110110110: data <= 20'hfff04; 
        10'b0110110111: data <= 20'h002a1; 
        10'b0110111000: data <= 20'h00634; 
        10'b0110111001: data <= 20'h0060f; 
        10'b0110111010: data <= 20'h00218; 
        10'b0110111011: data <= 20'h000cb; 
        10'b0110111100: data <= 20'hffc36; 
        10'b0110111101: data <= 20'hfff26; 
        10'b0110111110: data <= 20'hffecd; 
        10'b0110111111: data <= 20'hffcfc; 
        10'b0111000000: data <= 20'hffedd; 
        10'b0111000001: data <= 20'hfff5c; 
        10'b0111000010: data <= 20'h002c1; 
        10'b0111000011: data <= 20'h0007d; 
        10'b0111000100: data <= 20'h00205; 
        10'b0111000101: data <= 20'hffca8; 
        10'b0111000110: data <= 20'hffa82; 
        10'b0111000111: data <= 20'hff67e; 
        10'b0111001000: data <= 20'hfeb50; 
        10'b0111001001: data <= 20'hfea33; 
        10'b0111001010: data <= 20'hfecad; 
        10'b0111001011: data <= 20'hffb1b; 
        10'b0111001100: data <= 20'h005c4; 
        10'b0111001101: data <= 20'h00eed; 
        10'b0111001110: data <= 20'hffe63; 
        10'b0111001111: data <= 20'hff51c; 
        10'b0111010000: data <= 20'hff47b; 
        10'b0111010001: data <= 20'hffc40; 
        10'b0111010010: data <= 20'h004dc; 
        10'b0111010011: data <= 20'h00cbb; 
        10'b0111010100: data <= 20'h008f5; 
        10'b0111010101: data <= 20'h00b47; 
        10'b0111010110: data <= 20'h00af4; 
        10'b0111010111: data <= 20'h004d9; 
        10'b0111011000: data <= 20'hffe91; 
        10'b0111011001: data <= 20'hfff08; 
        10'b0111011010: data <= 20'hfffde; 
        10'b0111011011: data <= 20'hfffa4; 
        10'b0111011100: data <= 20'hfff8f; 
        10'b0111011101: data <= 20'h00077; 
        10'b0111011110: data <= 20'h0000f; 
        10'b0111011111: data <= 20'h006fa; 
        10'b0111100000: data <= 20'h003db; 
        10'b0111100001: data <= 20'h00135; 
        10'b0111100010: data <= 20'hffc4f; 
        10'b0111100011: data <= 20'hff372; 
        10'b0111100100: data <= 20'hfe9a5; 
        10'b0111100101: data <= 20'hfdc8d; 
        10'b0111100110: data <= 20'hfd3e3; 
        10'b0111100111: data <= 20'hfd7bc; 
        10'b0111101000: data <= 20'hfe16e; 
        10'b0111101001: data <= 20'hfee95; 
        10'b0111101010: data <= 20'hfefd6; 
        10'b0111101011: data <= 20'hff193; 
        10'b0111101100: data <= 20'hfff6d; 
        10'b0111101101: data <= 20'h00474; 
        10'b0111101110: data <= 20'h00828; 
        10'b0111101111: data <= 20'h00ce9; 
        10'b0111110000: data <= 20'h002ad; 
        10'b0111110001: data <= 20'h00f9f; 
        10'b0111110010: data <= 20'h00f99; 
        10'b0111110011: data <= 20'h004b2; 
        10'b0111110100: data <= 20'hffdb1; 
        10'b0111110101: data <= 20'hffcae; 
        10'b0111110110: data <= 20'hffcf9; 
        10'b0111110111: data <= 20'hffd3b; 
        10'b0111111000: data <= 20'hffe4a; 
        10'b0111111001: data <= 20'hffe65; 
        10'b0111111010: data <= 20'h0015b; 
        10'b0111111011: data <= 20'h00a52; 
        10'b0111111100: data <= 20'h0076e; 
        10'b0111111101: data <= 20'h0047b; 
        10'b0111111110: data <= 20'h00259; 
        10'b0111111111: data <= 20'hffd47; 
        10'b1000000000: data <= 20'hff80d; 
        10'b1000000001: data <= 20'hfe60d; 
        10'b1000000010: data <= 20'hfd9c7; 
        10'b1000000011: data <= 20'hfdbd6; 
        10'b1000000100: data <= 20'hfd455; 
        10'b1000000101: data <= 20'hfdc5c; 
        10'b1000000110: data <= 20'hfe974; 
        10'b1000000111: data <= 20'hffadf; 
        10'b1000001000: data <= 20'h0091a; 
        10'b1000001001: data <= 20'h00c45; 
        10'b1000001010: data <= 20'h00d39; 
        10'b1000001011: data <= 20'h00d12; 
        10'b1000001100: data <= 20'h00927; 
        10'b1000001101: data <= 20'h0123e; 
        10'b1000001110: data <= 20'h01107; 
        10'b1000001111: data <= 20'h00681; 
        10'b1000010000: data <= 20'hffa02; 
        10'b1000010001: data <= 20'hffbf1; 
        10'b1000010010: data <= 20'hffd0c; 
        10'b1000010011: data <= 20'hfff88; 
        10'b1000010100: data <= 20'hfff88; 
        10'b1000010101: data <= 20'hffd04; 
        10'b1000010110: data <= 20'hffe17; 
        10'b1000010111: data <= 20'h00cf0; 
        10'b1000011000: data <= 20'h00d32; 
        10'b1000011001: data <= 20'h00f80; 
        10'b1000011010: data <= 20'h00d5c; 
        10'b1000011011: data <= 20'h004e7; 
        10'b1000011100: data <= 20'h00179; 
        10'b1000011101: data <= 20'hffa8d; 
        10'b1000011110: data <= 20'hffc12; 
        10'b1000011111: data <= 20'hff3af; 
        10'b1000100000: data <= 20'hfee01; 
        10'b1000100001: data <= 20'hfecdc; 
        10'b1000100010: data <= 20'hff2f5; 
        10'b1000100011: data <= 20'h00498; 
        10'b1000100100: data <= 20'h00c51; 
        10'b1000100101: data <= 20'h00f66; 
        10'b1000100110: data <= 20'h01142; 
        10'b1000100111: data <= 20'h00f6f; 
        10'b1000101000: data <= 20'h00daa; 
        10'b1000101001: data <= 20'h00ff0; 
        10'b1000101010: data <= 20'h0061c; 
        10'b1000101011: data <= 20'h000b6; 
        10'b1000101100: data <= 20'hffaef; 
        10'b1000101101: data <= 20'hfff10; 
        10'b1000101110: data <= 20'hfff7f; 
        10'b1000101111: data <= 20'hffeeb; 
        10'b1000110000: data <= 20'hfff58; 
        10'b1000110001: data <= 20'hffc10; 
        10'b1000110010: data <= 20'h00254; 
        10'b1000110011: data <= 20'h00de2; 
        10'b1000110100: data <= 20'h01110; 
        10'b1000110101: data <= 20'h01278; 
        10'b1000110110: data <= 20'h01390; 
        10'b1000110111: data <= 20'h009df; 
        10'b1000111000: data <= 20'h00b9d; 
        10'b1000111001: data <= 20'h00d24; 
        10'b1000111010: data <= 20'h004da; 
        10'b1000111011: data <= 20'hffead; 
        10'b1000111100: data <= 20'hffb97; 
        10'b1000111101: data <= 20'hff93f; 
        10'b1000111110: data <= 20'h0020b; 
        10'b1000111111: data <= 20'h003a4; 
        10'b1001000000: data <= 20'h006f2; 
        10'b1001000001: data <= 20'h00c61; 
        10'b1001000010: data <= 20'h00cf7; 
        10'b1001000011: data <= 20'h008d3; 
        10'b1001000100: data <= 20'h00f5e; 
        10'b1001000101: data <= 20'h008bb; 
        10'b1001000110: data <= 20'hffe5f; 
        10'b1001000111: data <= 20'hffc80; 
        10'b1001001000: data <= 20'hffbf0; 
        10'b1001001001: data <= 20'hffecd; 
        10'b1001001010: data <= 20'hffec0; 
        10'b1001001011: data <= 20'hffe9b; 
        10'b1001001100: data <= 20'hffd5a; 
        10'b1001001101: data <= 20'hfffd2; 
        10'b1001001110: data <= 20'hfff0a; 
        10'b1001001111: data <= 20'h006e7; 
        10'b1001010000: data <= 20'h0107a; 
        10'b1001010001: data <= 20'h01074; 
        10'b1001010010: data <= 20'h00e5f; 
        10'b1001010011: data <= 20'h0081c; 
        10'b1001010100: data <= 20'h008a7; 
        10'b1001010101: data <= 20'h002dc; 
        10'b1001010110: data <= 20'hffedd; 
        10'b1001010111: data <= 20'hffc1c; 
        10'b1001011000: data <= 20'h0013f; 
        10'b1001011001: data <= 20'hfff4d; 
        10'b1001011010: data <= 20'hffefb; 
        10'b1001011011: data <= 20'hffe1a; 
        10'b1001011100: data <= 20'h00409; 
        10'b1001011101: data <= 20'h00179; 
        10'b1001011110: data <= 20'h007ea; 
        10'b1001011111: data <= 20'h00cba; 
        10'b1001100000: data <= 20'h00767; 
        10'b1001100001: data <= 20'h002d4; 
        10'b1001100010: data <= 20'hffd22; 
        10'b1001100011: data <= 20'hff89c; 
        10'b1001100100: data <= 20'hffd99; 
        10'b1001100101: data <= 20'hffcf4; 
        10'b1001100110: data <= 20'hffbfc; 
        10'b1001100111: data <= 20'hffc3c; 
        10'b1001101000: data <= 20'hffe58; 
        10'b1001101001: data <= 20'hffed9; 
        10'b1001101010: data <= 20'hfff3b; 
        10'b1001101011: data <= 20'h0044b; 
        10'b1001101100: data <= 20'h00846; 
        10'b1001101101: data <= 20'h00b43; 
        10'b1001101110: data <= 20'h00a0c; 
        10'b1001101111: data <= 20'h005b9; 
        10'b1001110000: data <= 20'h00072; 
        10'b1001110001: data <= 20'h00424; 
        10'b1001110010: data <= 20'h00500; 
        10'b1001110011: data <= 20'h00614; 
        10'b1001110100: data <= 20'h001af; 
        10'b1001110101: data <= 20'hffdca; 
        10'b1001110110: data <= 20'hffda5; 
        10'b1001110111: data <= 20'hffca7; 
        10'b1001111000: data <= 20'h0029f; 
        10'b1001111001: data <= 20'h00200; 
        10'b1001111010: data <= 20'h001f7; 
        10'b1001111011: data <= 20'h008cb; 
        10'b1001111100: data <= 20'h00444; 
        10'b1001111101: data <= 20'hffe7c; 
        10'b1001111110: data <= 20'hffe08; 
        10'b1001111111: data <= 20'hffd6d; 
        10'b1010000000: data <= 20'hffa59; 
        10'b1010000001: data <= 20'hffbc4; 
        10'b1010000010: data <= 20'hfff3b; 
        10'b1010000011: data <= 20'hfffe2; 
        10'b1010000100: data <= 20'hffed3; 
        10'b1010000101: data <= 20'hffcd3; 
        10'b1010000110: data <= 20'hffd5d; 
        10'b1010000111: data <= 20'h002d4; 
        10'b1010001000: data <= 20'h0090a; 
        10'b1010001001: data <= 20'h00da6; 
        10'b1010001010: data <= 20'h00a2b; 
        10'b1010001011: data <= 20'h00abd; 
        10'b1010001100: data <= 20'h00299; 
        10'b1010001101: data <= 20'h006e1; 
        10'b1010001110: data <= 20'h0045f; 
        10'b1010001111: data <= 20'hfffee; 
        10'b1010010000: data <= 20'hffc8e; 
        10'b1010010001: data <= 20'h0008d; 
        10'b1010010010: data <= 20'h00166; 
        10'b1010010011: data <= 20'h00371; 
        10'b1010010100: data <= 20'h00290; 
        10'b1010010101: data <= 20'h00551; 
        10'b1010010110: data <= 20'h00877; 
        10'b1010010111: data <= 20'hffe92; 
        10'b1010011000: data <= 20'hffa57; 
        10'b1010011001: data <= 20'hffa65; 
        10'b1010011010: data <= 20'hffd0c; 
        10'b1010011011: data <= 20'hffc4d; 
        10'b1010011100: data <= 20'hfffac; 
        10'b1010011101: data <= 20'hfff0b; 
        10'b1010011110: data <= 20'hffc7c; 
        10'b1010011111: data <= 20'hffcca; 
        10'b1010100000: data <= 20'hffd78; 
        10'b1010100001: data <= 20'h00067; 
        10'b1010100010: data <= 20'h0006d; 
        10'b1010100011: data <= 20'h0000e; 
        10'b1010100100: data <= 20'h005cf; 
        10'b1010100101: data <= 20'h0095b; 
        10'b1010100110: data <= 20'h00b06; 
        10'b1010100111: data <= 20'h00d02; 
        10'b1010101000: data <= 20'h00d37; 
        10'b1010101001: data <= 20'h00ad6; 
        10'b1010101010: data <= 20'h00fcb; 
        10'b1010101011: data <= 20'h010ad; 
        10'b1010101100: data <= 20'h01115; 
        10'b1010101101: data <= 20'h00d75; 
        10'b1010101110: data <= 20'h00bde; 
        10'b1010101111: data <= 20'h008c7; 
        10'b1010110000: data <= 20'h00861; 
        10'b1010110001: data <= 20'hfff46; 
        10'b1010110010: data <= 20'hff931; 
        10'b1010110011: data <= 20'hff694; 
        10'b1010110100: data <= 20'hff789; 
        10'b1010110101: data <= 20'hffad5; 
        10'b1010110110: data <= 20'hffb2d; 
        10'b1010110111: data <= 20'hffe93; 
        10'b1010111000: data <= 20'hffd9a; 
        10'b1010111001: data <= 20'hffff0; 
        10'b1010111010: data <= 20'hffd8c; 
        10'b1010111011: data <= 20'h00071; 
        10'b1010111100: data <= 20'hfffa0; 
        10'b1010111101: data <= 20'hffbf2; 
        10'b1010111110: data <= 20'h00050; 
        10'b1010111111: data <= 20'h000a8; 
        10'b1011000000: data <= 20'hffeff; 
        10'b1011000001: data <= 20'h003a7; 
        10'b1011000010: data <= 20'h0057f; 
        10'b1011000011: data <= 20'h00313; 
        10'b1011000100: data <= 20'h00768; 
        10'b1011000101: data <= 20'h0077d; 
        10'b1011000110: data <= 20'h00dff; 
        10'b1011000111: data <= 20'h01000; 
        10'b1011001000: data <= 20'h0112d; 
        10'b1011001001: data <= 20'h00d73; 
        10'b1011001010: data <= 20'h0098f; 
        10'b1011001011: data <= 20'h003d7; 
        10'b1011001100: data <= 20'hffe75; 
        10'b1011001101: data <= 20'hff9f1; 
        10'b1011001110: data <= 20'hff9e9; 
        10'b1011001111: data <= 20'hffb02; 
        10'b1011010000: data <= 20'hffb0c; 
        10'b1011010001: data <= 20'hffd81; 
        10'b1011010010: data <= 20'hffd81; 
        10'b1011010011: data <= 20'hfffbb; 
        10'b1011010100: data <= 20'hffcf9; 
        10'b1011010101: data <= 20'h00062; 
        10'b1011010110: data <= 20'hffc07; 
        10'b1011010111: data <= 20'hfff71; 
        10'b1011011000: data <= 20'hffd20; 
        10'b1011011001: data <= 20'hffbe9; 
        10'b1011011010: data <= 20'hffc19; 
        10'b1011011011: data <= 20'hfff00; 
        10'b1011011100: data <= 20'hfff0e; 
        10'b1011011101: data <= 20'hffd4e; 
        10'b1011011110: data <= 20'hffcdc; 
        10'b1011011111: data <= 20'hffee9; 
        10'b1011100000: data <= 20'hfff01; 
        10'b1011100001: data <= 20'hffeb1; 
        10'b1011100010: data <= 20'hffe2a; 
        10'b1011100011: data <= 20'hffe78; 
        10'b1011100100: data <= 20'hffdbb; 
        10'b1011100101: data <= 20'hffec7; 
        10'b1011100110: data <= 20'hffdb5; 
        10'b1011100111: data <= 20'hffb93; 
        10'b1011101000: data <= 20'hffd49; 
        10'b1011101001: data <= 20'hffeb6; 
        10'b1011101010: data <= 20'hffe38; 
        10'b1011101011: data <= 20'hffed7; 
        10'b1011101100: data <= 20'hffc2e; 
        10'b1011101101: data <= 20'hffc3f; 
        10'b1011101110: data <= 20'hfff6d; 
        10'b1011101111: data <= 20'hffdd1; 
        10'b1011110000: data <= 20'h0001a; 
        10'b1011110001: data <= 20'hffd0f; 
        10'b1011110010: data <= 20'hfffad; 
        10'b1011110011: data <= 20'h00074; 
        10'b1011110100: data <= 20'hffe0c; 
        10'b1011110101: data <= 20'hffcf2; 
        10'b1011110110: data <= 20'hffea6; 
        10'b1011110111: data <= 20'hffc2b; 
        10'b1011111000: data <= 20'h00033; 
        10'b1011111001: data <= 20'hffef5; 
        10'b1011111010: data <= 20'hfffce; 
        10'b1011111011: data <= 20'hffec8; 
        10'b1011111100: data <= 20'hfff60; 
        10'b1011111101: data <= 20'hffc1e; 
        10'b1011111110: data <= 20'hffcd1; 
        10'b1011111111: data <= 20'hfff29; 
        10'b1100000000: data <= 20'hffccd; 
        10'b1100000001: data <= 20'hfff66; 
        10'b1100000010: data <= 20'hffd9d; 
        10'b1100000011: data <= 20'hffe99; 
        10'b1100000100: data <= 20'hffdb9; 
        10'b1100000101: data <= 20'hfffed; 
        10'b1100000110: data <= 20'hffc54; 
        10'b1100000111: data <= 20'hffcf7; 
        10'b1100001000: data <= 20'hfffbe; 
        10'b1100001001: data <= 20'hffeac; 
        10'b1100001010: data <= 20'hffcf0; 
        10'b1100001011: data <= 20'hfff0c; 
        10'b1100001100: data <= 20'hffc61; 
        10'b1100001101: data <= 20'hffc13; 
        10'b1100001110: data <= 20'hfffc7; 
        10'b1100001111: data <= 20'hffe2d; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 15) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 21'h1ffd7b; 
        10'b0000000001: data <= 21'h1ff9c5; 
        10'b0000000010: data <= 21'h1fffb1; 
        10'b0000000011: data <= 21'h000048; 
        10'b0000000100: data <= 21'h0000a1; 
        10'b0000000101: data <= 21'h1fff74; 
        10'b0000000110: data <= 21'h1ffda2; 
        10'b0000000111: data <= 21'h0000a6; 
        10'b0000001000: data <= 21'h1ffaf8; 
        10'b0000001001: data <= 21'h000065; 
        10'b0000001010: data <= 21'h00006d; 
        10'b0000001011: data <= 21'h1ffbb6; 
        10'b0000001100: data <= 21'h1ffb9c; 
        10'b0000001101: data <= 21'h1ffb80; 
        10'b0000001110: data <= 21'h1ffbd7; 
        10'b0000001111: data <= 21'h1ffc62; 
        10'b0000010000: data <= 21'h000016; 
        10'b0000010001: data <= 21'h000047; 
        10'b0000010010: data <= 21'h1ff9c9; 
        10'b0000010011: data <= 21'h0000a2; 
        10'b0000010100: data <= 21'h1ffdfb; 
        10'b0000010101: data <= 21'h1ffe40; 
        10'b0000010110: data <= 21'h1ff7d6; 
        10'b0000010111: data <= 21'h1fff8d; 
        10'b0000011000: data <= 21'h1fffb2; 
        10'b0000011001: data <= 21'h1ff853; 
        10'b0000011010: data <= 21'h1ffc39; 
        10'b0000011011: data <= 21'h000039; 
        10'b0000011100: data <= 21'h1ff994; 
        10'b0000011101: data <= 21'h1ffbf9; 
        10'b0000011110: data <= 21'h1ff9ae; 
        10'b0000011111: data <= 21'h1ffdcd; 
        10'b0000100000: data <= 21'h1ff8c1; 
        10'b0000100001: data <= 21'h1ffc88; 
        10'b0000100010: data <= 21'h0000d5; 
        10'b0000100011: data <= 21'h000076; 
        10'b0000100100: data <= 21'h1ff847; 
        10'b0000100101: data <= 21'h1ff7ed; 
        10'b0000100110: data <= 21'h1ff8be; 
        10'b0000100111: data <= 21'h1ffd9e; 
        10'b0000101000: data <= 21'h1ffe47; 
        10'b0000101001: data <= 21'h1ffc4f; 
        10'b0000101010: data <= 21'h1ffbb0; 
        10'b0000101011: data <= 21'h1ffa31; 
        10'b0000101100: data <= 21'h0000cc; 
        10'b0000101101: data <= 21'h1ff9cc; 
        10'b0000101110: data <= 21'h1ffea0; 
        10'b0000101111: data <= 21'h1ffb45; 
        10'b0000110000: data <= 21'h1ffb5e; 
        10'b0000110001: data <= 21'h1ff87e; 
        10'b0000110010: data <= 21'h1ffcdf; 
        10'b0000110011: data <= 21'h1fff41; 
        10'b0000110100: data <= 21'h1ff939; 
        10'b0000110101: data <= 21'h1fff9b; 
        10'b0000110110: data <= 21'h1ffd52; 
        10'b0000110111: data <= 21'h1ff948; 
        10'b0000111000: data <= 21'h1ffa59; 
        10'b0000111001: data <= 21'h1ffcd5; 
        10'b0000111010: data <= 21'h1ffc9d; 
        10'b0000111011: data <= 21'h1ff9ce; 
        10'b0000111100: data <= 21'h1ffe06; 
        10'b0000111101: data <= 21'h1ffeac; 
        10'b0000111110: data <= 21'h1ffab8; 
        10'b0000111111: data <= 21'h1ffe91; 
        10'b0001000000: data <= 21'h1fff4d; 
        10'b0001000001: data <= 21'h1ffc4f; 
        10'b0001000010: data <= 21'h1ff919; 
        10'b0001000011: data <= 21'h1ff948; 
        10'b0001000100: data <= 21'h1ff870; 
        10'b0001000101: data <= 21'h1ff971; 
        10'b0001000110: data <= 21'h1ffbd9; 
        10'b0001000111: data <= 21'h1ffb40; 
        10'b0001001000: data <= 21'h1ffaa1; 
        10'b0001001001: data <= 21'h1ffa6f; 
        10'b0001001010: data <= 21'h1ffe92; 
        10'b0001001011: data <= 21'h1fffd6; 
        10'b0001001100: data <= 21'h1ffc25; 
        10'b0001001101: data <= 21'h1ff9a4; 
        10'b0001001110: data <= 21'h0000b3; 
        10'b0001001111: data <= 21'h1fff7b; 
        10'b0001010000: data <= 21'h000005; 
        10'b0001010001: data <= 21'h1ffb0a; 
        10'b0001010010: data <= 21'h1ff828; 
        10'b0001010011: data <= 21'h1ffc5a; 
        10'b0001010100: data <= 21'h0000de; 
        10'b0001010101: data <= 21'h1ffe81; 
        10'b0001010110: data <= 21'h1ffc73; 
        10'b0001010111: data <= 21'h1fff0c; 
        10'b0001011000: data <= 21'h1ffe69; 
        10'b0001011001: data <= 21'h000008; 
        10'b0001011010: data <= 21'h1ffda8; 
        10'b0001011011: data <= 21'h1fff8f; 
        10'b0001011100: data <= 21'h1fff18; 
        10'b0001011101: data <= 21'h1ffd02; 
        10'b0001011110: data <= 21'h0002c7; 
        10'b0001011111: data <= 21'h000943; 
        10'b0001100000: data <= 21'h00138e; 
        10'b0001100001: data <= 21'h00103f; 
        10'b0001100010: data <= 21'h00108f; 
        10'b0001100011: data <= 21'h001248; 
        10'b0001100100: data <= 21'h000cad; 
        10'b0001100101: data <= 21'h000e4b; 
        10'b0001100110: data <= 21'h000b2a; 
        10'b0001100111: data <= 21'h0000d6; 
        10'b0001101000: data <= 21'h1ffee3; 
        10'b0001101001: data <= 21'h1ff25c; 
        10'b0001101010: data <= 21'h1ff81d; 
        10'b0001101011: data <= 21'h1fff52; 
        10'b0001101100: data <= 21'h000062; 
        10'b0001101101: data <= 21'h1ffa03; 
        10'b0001101110: data <= 21'h1ffd47; 
        10'b0001101111: data <= 21'h1ffac0; 
        10'b0001110000: data <= 21'h1ffd31; 
        10'b0001110001: data <= 21'h1fff8b; 
        10'b0001110010: data <= 21'h1ffde0; 
        10'b0001110011: data <= 21'h00003d; 
        10'b0001110100: data <= 21'h0002f9; 
        10'b0001110101: data <= 21'h1ffff9; 
        10'b0001110110: data <= 21'h000b7d; 
        10'b0001110111: data <= 21'h0009b2; 
        10'b0001111000: data <= 21'h001a71; 
        10'b0001111001: data <= 21'h0016b8; 
        10'b0001111010: data <= 21'h001c2b; 
        10'b0001111011: data <= 21'h0021e3; 
        10'b0001111100: data <= 21'h002750; 
        10'b0001111101: data <= 21'h002a22; 
        10'b0001111110: data <= 21'h0025e1; 
        10'b0001111111: data <= 21'h001bc6; 
        10'b0010000000: data <= 21'h000fa9; 
        10'b0010000001: data <= 21'h000c88; 
        10'b0010000010: data <= 21'h00147b; 
        10'b0010000011: data <= 21'h000284; 
        10'b0010000100: data <= 21'h1ff1fa; 
        10'b0010000101: data <= 21'h1fea21; 
        10'b0010000110: data <= 21'h1fed4f; 
        10'b0010000111: data <= 21'h1fedb6; 
        10'b0010001000: data <= 21'h1ffdc7; 
        10'b0010001001: data <= 21'h1ffcac; 
        10'b0010001010: data <= 21'h1ffb3b; 
        10'b0010001011: data <= 21'h1ffec0; 
        10'b0010001100: data <= 21'h1ff91b; 
        10'b0010001101: data <= 21'h1ff81b; 
        10'b0010001110: data <= 21'h1ffa1a; 
        10'b0010001111: data <= 21'h1ffa1c; 
        10'b0010010000: data <= 21'h00017a; 
        10'b0010010001: data <= 21'h000bf2; 
        10'b0010010010: data <= 21'h0015d6; 
        10'b0010010011: data <= 21'h001172; 
        10'b0010010100: data <= 21'h0013f9; 
        10'b0010010101: data <= 21'h00119f; 
        10'b0010010110: data <= 21'h000ff3; 
        10'b0010010111: data <= 21'h0014c4; 
        10'b0010011000: data <= 21'h001515; 
        10'b0010011001: data <= 21'h00194b; 
        10'b0010011010: data <= 21'h000453; 
        10'b0010011011: data <= 21'h0010d9; 
        10'b0010011100: data <= 21'h001374; 
        10'b0010011101: data <= 21'h1ffe81; 
        10'b0010011110: data <= 21'h1ffef6; 
        10'b0010011111: data <= 21'h1ff72e; 
        10'b0010100000: data <= 21'h1ff3bd; 
        10'b0010100001: data <= 21'h1fe5f9; 
        10'b0010100010: data <= 21'h1fdeb7; 
        10'b0010100011: data <= 21'h1fe3d4; 
        10'b0010100100: data <= 21'h1ff7d6; 
        10'b0010100101: data <= 21'h000009; 
        10'b0010100110: data <= 21'h1ffa62; 
        10'b0010100111: data <= 21'h1ffc8d; 
        10'b0010101000: data <= 21'h1ff9d0; 
        10'b0010101001: data <= 21'h1ffb24; 
        10'b0010101010: data <= 21'h1ffa9c; 
        10'b0010101011: data <= 21'h000284; 
        10'b0010101100: data <= 21'h000ecb; 
        10'b0010101101: data <= 21'h001b80; 
        10'b0010101110: data <= 21'h001508; 
        10'b0010101111: data <= 21'h00101e; 
        10'b0010110000: data <= 21'h001868; 
        10'b0010110001: data <= 21'h0013e9; 
        10'b0010110010: data <= 21'h0011b2; 
        10'b0010110011: data <= 21'h0010ee; 
        10'b0010110100: data <= 21'h0016a5; 
        10'b0010110101: data <= 21'h00207c; 
        10'b0010110110: data <= 21'h001695; 
        10'b0010110111: data <= 21'h000828; 
        10'b0010111000: data <= 21'h00157d; 
        10'b0010111001: data <= 21'h0013b3; 
        10'b0010111010: data <= 21'h0012c1; 
        10'b0010111011: data <= 21'h1ff79d; 
        10'b0010111100: data <= 21'h000800; 
        10'b0010111101: data <= 21'h1ff812; 
        10'b0010111110: data <= 21'h1fe36f; 
        10'b0010111111: data <= 21'h1fe36f; 
        10'b0011000000: data <= 21'h1fee81; 
        10'b0011000001: data <= 21'h1ffc7b; 
        10'b0011000010: data <= 21'h1fff39; 
        10'b0011000011: data <= 21'h1ffd40; 
        10'b0011000100: data <= 21'h000056; 
        10'b0011000101: data <= 21'h1fff09; 
        10'b0011000110: data <= 21'h0001ae; 
        10'b0011000111: data <= 21'h000c58; 
        10'b0011001000: data <= 21'h002078; 
        10'b0011001001: data <= 21'h00204d; 
        10'b0011001010: data <= 21'h0016c2; 
        10'b0011001011: data <= 21'h000666; 
        10'b0011001100: data <= 21'h0006dc; 
        10'b0011001101: data <= 21'h000e78; 
        10'b0011001110: data <= 21'h000470; 
        10'b0011001111: data <= 21'h000698; 
        10'b0011010000: data <= 21'h00130c; 
        10'b0011010001: data <= 21'h001209; 
        10'b0011010010: data <= 21'h001de4; 
        10'b0011010011: data <= 21'h001190; 
        10'b0011010100: data <= 21'h000562; 
        10'b0011010101: data <= 21'h000f00; 
        10'b0011010110: data <= 21'h000c6f; 
        10'b0011010111: data <= 21'h000d83; 
        10'b0011011000: data <= 21'h000db1; 
        10'b0011011001: data <= 21'h0001f0; 
        10'b0011011010: data <= 21'h1ff235; 
        10'b0011011011: data <= 21'h1fdff2; 
        10'b0011011100: data <= 21'h1fe903; 
        10'b0011011101: data <= 21'h1ff9f7; 
        10'b0011011110: data <= 21'h1ff824; 
        10'b0011011111: data <= 21'h1ffbce; 
        10'b0011100000: data <= 21'h1ffcf4; 
        10'b0011100001: data <= 21'h1ffb4b; 
        10'b0011100010: data <= 21'h00015d; 
        10'b0011100011: data <= 21'h000b87; 
        10'b0011100100: data <= 21'h001ac4; 
        10'b0011100101: data <= 21'h00196e; 
        10'b0011100110: data <= 21'h00131d; 
        10'b0011100111: data <= 21'h0007ce; 
        10'b0011101000: data <= 21'h000cf2; 
        10'b0011101001: data <= 21'h00062c; 
        10'b0011101010: data <= 21'h00105a; 
        10'b0011101011: data <= 21'h00053f; 
        10'b0011101100: data <= 21'h000477; 
        10'b0011101101: data <= 21'h0007ff; 
        10'b0011101110: data <= 21'h002080; 
        10'b0011101111: data <= 21'h001af6; 
        10'b0011110000: data <= 21'h000638; 
        10'b0011110001: data <= 21'h000efc; 
        10'b0011110010: data <= 21'h001589; 
        10'b0011110011: data <= 21'h000e09; 
        10'b0011110100: data <= 21'h001489; 
        10'b0011110101: data <= 21'h000a93; 
        10'b0011110110: data <= 21'h1ffa81; 
        10'b0011110111: data <= 21'h1fe24b; 
        10'b0011111000: data <= 21'h1fe9c1; 
        10'b0011111001: data <= 21'h1ff7e2; 
        10'b0011111010: data <= 21'h1ff919; 
        10'b0011111011: data <= 21'h1ffb09; 
        10'b0011111100: data <= 21'h1ffc1a; 
        10'b0011111101: data <= 21'h1ff85e; 
        10'b0011111110: data <= 21'h1ffd90; 
        10'b0011111111: data <= 21'h0004f8; 
        10'b0100000000: data <= 21'h000dd5; 
        10'b0100000001: data <= 21'h00125a; 
        10'b0100000010: data <= 21'h000f32; 
        10'b0100000011: data <= 21'h0003b1; 
        10'b0100000100: data <= 21'h1ffe13; 
        10'b0100000101: data <= 21'h1ff1d3; 
        10'b0100000110: data <= 21'h1fe4fa; 
        10'b0100000111: data <= 21'h1fce61; 
        10'b0100001000: data <= 21'h1fd7bd; 
        10'b0100001001: data <= 21'h1ffaa3; 
        10'b0100001010: data <= 21'h0026b5; 
        10'b0100001011: data <= 21'h003b80; 
        10'b0100001100: data <= 21'h00225f; 
        10'b0100001101: data <= 21'h00141a; 
        10'b0100001110: data <= 21'h0015d9; 
        10'b0100001111: data <= 21'h001431; 
        10'b0100010000: data <= 21'h001e3f; 
        10'b0100010001: data <= 21'h00134d; 
        10'b0100010010: data <= 21'h1ffa27; 
        10'b0100010011: data <= 21'h1fe27e; 
        10'b0100010100: data <= 21'h1ff127; 
        10'b0100010101: data <= 21'h1ff7a0; 
        10'b0100010110: data <= 21'h1ff9b4; 
        10'b0100010111: data <= 21'h1ffabf; 
        10'b0100011000: data <= 21'h1fff28; 
        10'b0100011001: data <= 21'h1ffebe; 
        10'b0100011010: data <= 21'h00006a; 
        10'b0100011011: data <= 21'h000775; 
        10'b0100011100: data <= 21'h0006b4; 
        10'b0100011101: data <= 21'h0002db; 
        10'b0100011110: data <= 21'h1ff75a; 
        10'b0100011111: data <= 21'h1fea17; 
        10'b0100100000: data <= 21'h1fd7ec; 
        10'b0100100001: data <= 21'h1fc6b5; 
        10'b0100100010: data <= 21'h1fb9cb; 
        10'b0100100011: data <= 21'h1fb7ff; 
        10'b0100100100: data <= 21'h1fcaf5; 
        10'b0100100101: data <= 21'h1ff29d; 
        10'b0100100110: data <= 21'h001fbd; 
        10'b0100100111: data <= 21'h0024b1; 
        10'b0100101000: data <= 21'h001f3c; 
        10'b0100101001: data <= 21'h001d20; 
        10'b0100101010: data <= 21'h0011fa; 
        10'b0100101011: data <= 21'h001f2f; 
        10'b0100101100: data <= 21'h001cf2; 
        10'b0100101101: data <= 21'h000b98; 
        10'b0100101110: data <= 21'h1ff5a0; 
        10'b0100101111: data <= 21'h1fecdc; 
        10'b0100110000: data <= 21'h1ff8d8; 
        10'b0100110001: data <= 21'h1ff7e6; 
        10'b0100110010: data <= 21'h1ffc92; 
        10'b0100110011: data <= 21'h1fff21; 
        10'b0100110100: data <= 21'h0000f1; 
        10'b0100110101: data <= 21'h1fff21; 
        10'b0100110110: data <= 21'h1ff95f; 
        10'b0100110111: data <= 21'h000744; 
        10'b0100111000: data <= 21'h1ffbb4; 
        10'b0100111001: data <= 21'h1fe989; 
        10'b0100111010: data <= 21'h1fde4d; 
        10'b0100111011: data <= 21'h1fce76; 
        10'b0100111100: data <= 21'h1fc213; 
        10'b0100111101: data <= 21'h1fca7c; 
        10'b0100111110: data <= 21'h1fd741; 
        10'b0100111111: data <= 21'h1feccb; 
        10'b0101000000: data <= 21'h1ff599; 
        10'b0101000001: data <= 21'h000d73; 
        10'b0101000010: data <= 21'h00151f; 
        10'b0101000011: data <= 21'h00153c; 
        10'b0101000100: data <= 21'h0009b1; 
        10'b0101000101: data <= 21'h0015fd; 
        10'b0101000110: data <= 21'h001b36; 
        10'b0101000111: data <= 21'h001a88; 
        10'b0101001000: data <= 21'h001729; 
        10'b0101001001: data <= 21'h00001c; 
        10'b0101001010: data <= 21'h1ff5cd; 
        10'b0101001011: data <= 21'h1ff777; 
        10'b0101001100: data <= 21'h1ff87d; 
        10'b0101001101: data <= 21'h1ffb8d; 
        10'b0101001110: data <= 21'h1ff9d7; 
        10'b0101001111: data <= 21'h1ff91a; 
        10'b0101010000: data <= 21'h000044; 
        10'b0101010001: data <= 21'h1ffacc; 
        10'b0101010010: data <= 21'h1ffead; 
        10'b0101010011: data <= 21'h1fff99; 
        10'b0101010100: data <= 21'h1ff7d5; 
        10'b0101010101: data <= 21'h1fe973; 
        10'b0101010110: data <= 21'h1fd886; 
        10'b0101010111: data <= 21'h1fce9c; 
        10'b0101011000: data <= 21'h1fd356; 
        10'b0101011001: data <= 21'h1fe837; 
        10'b0101011010: data <= 21'h000078; 
        10'b0101011011: data <= 21'h0003f7; 
        10'b0101011100: data <= 21'h000649; 
        10'b0101011101: data <= 21'h000e45; 
        10'b0101011110: data <= 21'h002359; 
        10'b0101011111: data <= 21'h001244; 
        10'b0101100000: data <= 21'h000c7a; 
        10'b0101100001: data <= 21'h0011a6; 
        10'b0101100010: data <= 21'h000e24; 
        10'b0101100011: data <= 21'h1ffec4; 
        10'b0101100100: data <= 21'h1fedb3; 
        10'b0101100101: data <= 21'h1fe6de; 
        10'b0101100110: data <= 21'h1fe5b1; 
        10'b0101100111: data <= 21'h1fef46; 
        10'b0101101000: data <= 21'h1ffd10; 
        10'b0101101001: data <= 21'h1ffaee; 
        10'b0101101010: data <= 21'h1ffd44; 
        10'b0101101011: data <= 21'h1ffe13; 
        10'b0101101100: data <= 21'h1ffc6f; 
        10'b0101101101: data <= 21'h1ffa98; 
        10'b0101101110: data <= 21'h1ffcae; 
        10'b0101101111: data <= 21'h1ffdc7; 
        10'b0101110000: data <= 21'h1ff58e; 
        10'b0101110001: data <= 21'h1ff096; 
        10'b0101110010: data <= 21'h1fdfe4; 
        10'b0101110011: data <= 21'h1fdaee; 
        10'b0101110100: data <= 21'h1fe6db; 
        10'b0101110101: data <= 21'h1ffb0d; 
        10'b0101110110: data <= 21'h1ff7d4; 
        10'b0101110111: data <= 21'h1feab0; 
        10'b0101111000: data <= 21'h0001b2; 
        10'b0101111001: data <= 21'h001e6e; 
        10'b0101111010: data <= 21'h001ebc; 
        10'b0101111011: data <= 21'h00059c; 
        10'b0101111100: data <= 21'h000df4; 
        10'b0101111101: data <= 21'h000ee0; 
        10'b0101111110: data <= 21'h0007e5; 
        10'b0101111111: data <= 21'h1ff587; 
        10'b0110000000: data <= 21'h1fe3f2; 
        10'b0110000001: data <= 21'h1fe3cf; 
        10'b0110000010: data <= 21'h1fe9bc; 
        10'b0110000011: data <= 21'h1ff05c; 
        10'b0110000100: data <= 21'h1ff705; 
        10'b0110000101: data <= 21'h1fffcf; 
        10'b0110000110: data <= 21'h1ffe5d; 
        10'b0110000111: data <= 21'h1ffb38; 
        10'b0110001000: data <= 21'h0000be; 
        10'b0110001001: data <= 21'h1ff9e5; 
        10'b0110001010: data <= 21'h1ffc18; 
        10'b0110001011: data <= 21'h1ffd75; 
        10'b0110001100: data <= 21'h1ffe11; 
        10'b0110001101: data <= 21'h1ff31b; 
        10'b0110001110: data <= 21'h1fe307; 
        10'b0110001111: data <= 21'h1fe5d0; 
        10'b0110010000: data <= 21'h1fee37; 
        10'b0110010001: data <= 21'h1ffd88; 
        10'b0110010010: data <= 21'h1fed59; 
        10'b0110010011: data <= 21'h1fec1e; 
        10'b0110010100: data <= 21'h0005a3; 
        10'b0110010101: data <= 21'h000eb9; 
        10'b0110010110: data <= 21'h000fb8; 
        10'b0110010111: data <= 21'h1ffdaa; 
        10'b0110011000: data <= 21'h1ff99d; 
        10'b0110011001: data <= 21'h1ffb3e; 
        10'b0110011010: data <= 21'h000225; 
        10'b0110011011: data <= 21'h1ff3cd; 
        10'b0110011100: data <= 21'h1fef7d; 
        10'b0110011101: data <= 21'h1ff800; 
        10'b0110011110: data <= 21'h1ff4a3; 
        10'b0110011111: data <= 21'h1ff854; 
        10'b0110100000: data <= 21'h1ff5e7; 
        10'b0110100001: data <= 21'h1ff6ec; 
        10'b0110100010: data <= 21'h00003a; 
        10'b0110100011: data <= 21'h000074; 
        10'b0110100100: data <= 21'h0000aa; 
        10'b0110100101: data <= 21'h1ff9fe; 
        10'b0110100110: data <= 21'h0000e8; 
        10'b0110100111: data <= 21'h000239; 
        10'b0110101000: data <= 21'h1ffd69; 
        10'b0110101001: data <= 21'h1ff184; 
        10'b0110101010: data <= 21'h1fe51f; 
        10'b0110101011: data <= 21'h1fe33c; 
        10'b0110101100: data <= 21'h1fea7b; 
        10'b0110101101: data <= 21'h1ff362; 
        10'b0110101110: data <= 21'h1ff206; 
        10'b0110101111: data <= 21'h1ffb47; 
        10'b0110110000: data <= 21'h0005cf; 
        10'b0110110001: data <= 21'h0017ef; 
        10'b0110110010: data <= 21'h000dbd; 
        10'b0110110011: data <= 21'h1ffea5; 
        10'b0110110100: data <= 21'h1fec06; 
        10'b0110110101: data <= 21'h1ffa33; 
        10'b0110110110: data <= 21'h1ffe08; 
        10'b0110110111: data <= 21'h000541; 
        10'b0110111000: data <= 21'h000c68; 
        10'b0110111001: data <= 21'h000c1d; 
        10'b0110111010: data <= 21'h00042f; 
        10'b0110111011: data <= 21'h000197; 
        10'b0110111100: data <= 21'h1ff86b; 
        10'b0110111101: data <= 21'h1ffe4d; 
        10'b0110111110: data <= 21'h1ffd9a; 
        10'b0110111111: data <= 21'h1ff9f7; 
        10'b0111000000: data <= 21'h1ffdbb; 
        10'b0111000001: data <= 21'h1ffeb7; 
        10'b0111000010: data <= 21'h000583; 
        10'b0111000011: data <= 21'h0000fa; 
        10'b0111000100: data <= 21'h00040a; 
        10'b0111000101: data <= 21'h1ff950; 
        10'b0111000110: data <= 21'h1ff504; 
        10'b0111000111: data <= 21'h1fecfd; 
        10'b0111001000: data <= 21'h1fd69f; 
        10'b0111001001: data <= 21'h1fd465; 
        10'b0111001010: data <= 21'h1fd95b; 
        10'b0111001011: data <= 21'h1ff636; 
        10'b0111001100: data <= 21'h000b87; 
        10'b0111001101: data <= 21'h001dda; 
        10'b0111001110: data <= 21'h1ffcc6; 
        10'b0111001111: data <= 21'h1fea37; 
        10'b0111010000: data <= 21'h1fe8f6; 
        10'b0111010001: data <= 21'h1ff880; 
        10'b0111010010: data <= 21'h0009b8; 
        10'b0111010011: data <= 21'h001976; 
        10'b0111010100: data <= 21'h0011eb; 
        10'b0111010101: data <= 21'h00168d; 
        10'b0111010110: data <= 21'h0015e7; 
        10'b0111010111: data <= 21'h0009b2; 
        10'b0111011000: data <= 21'h1ffd22; 
        10'b0111011001: data <= 21'h1ffe10; 
        10'b0111011010: data <= 21'h1fffbc; 
        10'b0111011011: data <= 21'h1fff48; 
        10'b0111011100: data <= 21'h1fff1e; 
        10'b0111011101: data <= 21'h0000ef; 
        10'b0111011110: data <= 21'h00001f; 
        10'b0111011111: data <= 21'h000df4; 
        10'b0111100000: data <= 21'h0007b6; 
        10'b0111100001: data <= 21'h00026a; 
        10'b0111100010: data <= 21'h1ff89e; 
        10'b0111100011: data <= 21'h1fe6e4; 
        10'b0111100100: data <= 21'h1fd34a; 
        10'b0111100101: data <= 21'h1fb91b; 
        10'b0111100110: data <= 21'h1fa7c5; 
        10'b0111100111: data <= 21'h1faf78; 
        10'b0111101000: data <= 21'h1fc2dc; 
        10'b0111101001: data <= 21'h1fdd2a; 
        10'b0111101010: data <= 21'h1fdfac; 
        10'b0111101011: data <= 21'h1fe326; 
        10'b0111101100: data <= 21'h1ffeda; 
        10'b0111101101: data <= 21'h0008e8; 
        10'b0111101110: data <= 21'h001050; 
        10'b0111101111: data <= 21'h0019d2; 
        10'b0111110000: data <= 21'h00055a; 
        10'b0111110001: data <= 21'h001f3f; 
        10'b0111110010: data <= 21'h001f31; 
        10'b0111110011: data <= 21'h000963; 
        10'b0111110100: data <= 21'h1ffb63; 
        10'b0111110101: data <= 21'h1ff95b; 
        10'b0111110110: data <= 21'h1ff9f1; 
        10'b0111110111: data <= 21'h1ffa77; 
        10'b0111111000: data <= 21'h1ffc95; 
        10'b0111111001: data <= 21'h1ffccb; 
        10'b0111111010: data <= 21'h0002b5; 
        10'b0111111011: data <= 21'h0014a3; 
        10'b0111111100: data <= 21'h000edc; 
        10'b0111111101: data <= 21'h0008f6; 
        10'b0111111110: data <= 21'h0004b2; 
        10'b0111111111: data <= 21'h1ffa8d; 
        10'b1000000000: data <= 21'h1ff01b; 
        10'b1000000001: data <= 21'h1fcc1a; 
        10'b1000000010: data <= 21'h1fb38f; 
        10'b1000000011: data <= 21'h1fb7ad; 
        10'b1000000100: data <= 21'h1fa8aa; 
        10'b1000000101: data <= 21'h1fb8b8; 
        10'b1000000110: data <= 21'h1fd2e9; 
        10'b1000000111: data <= 21'h1ff5bf; 
        10'b1000001000: data <= 21'h001234; 
        10'b1000001001: data <= 21'h00188a; 
        10'b1000001010: data <= 21'h001a71; 
        10'b1000001011: data <= 21'h001a24; 
        10'b1000001100: data <= 21'h00124e; 
        10'b1000001101: data <= 21'h00247d; 
        10'b1000001110: data <= 21'h00220e; 
        10'b1000001111: data <= 21'h000d03; 
        10'b1000010000: data <= 21'h1ff404; 
        10'b1000010001: data <= 21'h1ff7e2; 
        10'b1000010010: data <= 21'h1ffa18; 
        10'b1000010011: data <= 21'h1fff0f; 
        10'b1000010100: data <= 21'h1fff11; 
        10'b1000010101: data <= 21'h1ffa08; 
        10'b1000010110: data <= 21'h1ffc2d; 
        10'b1000010111: data <= 21'h0019e0; 
        10'b1000011000: data <= 21'h001a64; 
        10'b1000011001: data <= 21'h001f01; 
        10'b1000011010: data <= 21'h001ab8; 
        10'b1000011011: data <= 21'h0009ce; 
        10'b1000011100: data <= 21'h0002f1; 
        10'b1000011101: data <= 21'h1ff51a; 
        10'b1000011110: data <= 21'h1ff825; 
        10'b1000011111: data <= 21'h1fe75d; 
        10'b1000100000: data <= 21'h1fdc02; 
        10'b1000100001: data <= 21'h1fd9b7; 
        10'b1000100010: data <= 21'h1fe5ea; 
        10'b1000100011: data <= 21'h000931; 
        10'b1000100100: data <= 21'h0018a2; 
        10'b1000100101: data <= 21'h001ecc; 
        10'b1000100110: data <= 21'h002284; 
        10'b1000100111: data <= 21'h001edf; 
        10'b1000101000: data <= 21'h001b54; 
        10'b1000101001: data <= 21'h001fe1; 
        10'b1000101010: data <= 21'h000c38; 
        10'b1000101011: data <= 21'h00016c; 
        10'b1000101100: data <= 21'h1ff5dd; 
        10'b1000101101: data <= 21'h1ffe20; 
        10'b1000101110: data <= 21'h1ffefd; 
        10'b1000101111: data <= 21'h1ffdd5; 
        10'b1000110000: data <= 21'h1ffeb1; 
        10'b1000110001: data <= 21'h1ff820; 
        10'b1000110010: data <= 21'h0004a8; 
        10'b1000110011: data <= 21'h001bc4; 
        10'b1000110100: data <= 21'h002221; 
        10'b1000110101: data <= 21'h0024f1; 
        10'b1000110110: data <= 21'h00271f; 
        10'b1000110111: data <= 21'h0013bd; 
        10'b1000111000: data <= 21'h00173a; 
        10'b1000111001: data <= 21'h001a48; 
        10'b1000111010: data <= 21'h0009b4; 
        10'b1000111011: data <= 21'h1ffd5a; 
        10'b1000111100: data <= 21'h1ff72d; 
        10'b1000111101: data <= 21'h1ff27e; 
        10'b1000111110: data <= 21'h000416; 
        10'b1000111111: data <= 21'h000748; 
        10'b1001000000: data <= 21'h000de5; 
        10'b1001000001: data <= 21'h0018c2; 
        10'b1001000010: data <= 21'h0019ef; 
        10'b1001000011: data <= 21'h0011a6; 
        10'b1001000100: data <= 21'h001ebc; 
        10'b1001000101: data <= 21'h001176; 
        10'b1001000110: data <= 21'h1ffcbf; 
        10'b1001000111: data <= 21'h1ff900; 
        10'b1001001000: data <= 21'h1ff7e0; 
        10'b1001001001: data <= 21'h1ffd9a; 
        10'b1001001010: data <= 21'h1ffd7f; 
        10'b1001001011: data <= 21'h1ffd35; 
        10'b1001001100: data <= 21'h1ffab4; 
        10'b1001001101: data <= 21'h1fffa3; 
        10'b1001001110: data <= 21'h1ffe14; 
        10'b1001001111: data <= 21'h000dce; 
        10'b1001010000: data <= 21'h0020f4; 
        10'b1001010001: data <= 21'h0020e8; 
        10'b1001010010: data <= 21'h001cbe; 
        10'b1001010011: data <= 21'h001037; 
        10'b1001010100: data <= 21'h00114d; 
        10'b1001010101: data <= 21'h0005b9; 
        10'b1001010110: data <= 21'h1ffdb9; 
        10'b1001010111: data <= 21'h1ff839; 
        10'b1001011000: data <= 21'h00027e; 
        10'b1001011001: data <= 21'h1ffe9a; 
        10'b1001011010: data <= 21'h1ffdf6; 
        10'b1001011011: data <= 21'h1ffc34; 
        10'b1001011100: data <= 21'h000812; 
        10'b1001011101: data <= 21'h0002f2; 
        10'b1001011110: data <= 21'h000fd4; 
        10'b1001011111: data <= 21'h001973; 
        10'b1001100000: data <= 21'h000ecd; 
        10'b1001100001: data <= 21'h0005a9; 
        10'b1001100010: data <= 21'h1ffa44; 
        10'b1001100011: data <= 21'h1ff138; 
        10'b1001100100: data <= 21'h1ffb32; 
        10'b1001100101: data <= 21'h1ff9e7; 
        10'b1001100110: data <= 21'h1ff7f8; 
        10'b1001100111: data <= 21'h1ff879; 
        10'b1001101000: data <= 21'h1ffcaf; 
        10'b1001101001: data <= 21'h1ffdb1; 
        10'b1001101010: data <= 21'h1ffe77; 
        10'b1001101011: data <= 21'h000896; 
        10'b1001101100: data <= 21'h00108c; 
        10'b1001101101: data <= 21'h001687; 
        10'b1001101110: data <= 21'h001419; 
        10'b1001101111: data <= 21'h000b72; 
        10'b1001110000: data <= 21'h0000e4; 
        10'b1001110001: data <= 21'h000848; 
        10'b1001110010: data <= 21'h000a00; 
        10'b1001110011: data <= 21'h000c28; 
        10'b1001110100: data <= 21'h00035d; 
        10'b1001110101: data <= 21'h1ffb93; 
        10'b1001110110: data <= 21'h1ffb4a; 
        10'b1001110111: data <= 21'h1ff94d; 
        10'b1001111000: data <= 21'h00053d; 
        10'b1001111001: data <= 21'h0003ff; 
        10'b1001111010: data <= 21'h0003ef; 
        10'b1001111011: data <= 21'h001196; 
        10'b1001111100: data <= 21'h000888; 
        10'b1001111101: data <= 21'h1ffcf9; 
        10'b1001111110: data <= 21'h1ffc10; 
        10'b1001111111: data <= 21'h1ffadb; 
        10'b1010000000: data <= 21'h1ff4b2; 
        10'b1010000001: data <= 21'h1ff788; 
        10'b1010000010: data <= 21'h1ffe77; 
        10'b1010000011: data <= 21'h1fffc4; 
        10'b1010000100: data <= 21'h1ffda5; 
        10'b1010000101: data <= 21'h1ff9a6; 
        10'b1010000110: data <= 21'h1ffaba; 
        10'b1010000111: data <= 21'h0005a7; 
        10'b1010001000: data <= 21'h001213; 
        10'b1010001001: data <= 21'h001b4c; 
        10'b1010001010: data <= 21'h001457; 
        10'b1010001011: data <= 21'h00157a; 
        10'b1010001100: data <= 21'h000532; 
        10'b1010001101: data <= 21'h000dc1; 
        10'b1010001110: data <= 21'h0008be; 
        10'b1010001111: data <= 21'h1fffdd; 
        10'b1010010000: data <= 21'h1ff91c; 
        10'b1010010001: data <= 21'h00011a; 
        10'b1010010010: data <= 21'h0002cc; 
        10'b1010010011: data <= 21'h0006e1; 
        10'b1010010100: data <= 21'h00051f; 
        10'b1010010101: data <= 21'h000aa2; 
        10'b1010010110: data <= 21'h0010ee; 
        10'b1010010111: data <= 21'h1ffd24; 
        10'b1010011000: data <= 21'h1ff4ad; 
        10'b1010011001: data <= 21'h1ff4cb; 
        10'b1010011010: data <= 21'h1ffa18; 
        10'b1010011011: data <= 21'h1ff89b; 
        10'b1010011100: data <= 21'h1fff58; 
        10'b1010011101: data <= 21'h1ffe16; 
        10'b1010011110: data <= 21'h1ff8f9; 
        10'b1010011111: data <= 21'h1ff994; 
        10'b1010100000: data <= 21'h1ffaf1; 
        10'b1010100001: data <= 21'h0000cd; 
        10'b1010100010: data <= 21'h0000d9; 
        10'b1010100011: data <= 21'h00001b; 
        10'b1010100100: data <= 21'h000b9e; 
        10'b1010100101: data <= 21'h0012b6; 
        10'b1010100110: data <= 21'h00160b; 
        10'b1010100111: data <= 21'h001a04; 
        10'b1010101000: data <= 21'h001a6d; 
        10'b1010101001: data <= 21'h0015ad; 
        10'b1010101010: data <= 21'h001f96; 
        10'b1010101011: data <= 21'h00215b; 
        10'b1010101100: data <= 21'h00222a; 
        10'b1010101101: data <= 21'h001ae9; 
        10'b1010101110: data <= 21'h0017bc; 
        10'b1010101111: data <= 21'h00118e; 
        10'b1010110000: data <= 21'h0010c2; 
        10'b1010110001: data <= 21'h1ffe8b; 
        10'b1010110010: data <= 21'h1ff262; 
        10'b1010110011: data <= 21'h1fed28; 
        10'b1010110100: data <= 21'h1fef12; 
        10'b1010110101: data <= 21'h1ff5ab; 
        10'b1010110110: data <= 21'h1ff659; 
        10'b1010110111: data <= 21'h1ffd26; 
        10'b1010111000: data <= 21'h1ffb34; 
        10'b1010111001: data <= 21'h1fffe0; 
        10'b1010111010: data <= 21'h1ffb17; 
        10'b1010111011: data <= 21'h0000e2; 
        10'b1010111100: data <= 21'h1fff40; 
        10'b1010111101: data <= 21'h1ff7e4; 
        10'b1010111110: data <= 21'h00009f; 
        10'b1010111111: data <= 21'h000150; 
        10'b1011000000: data <= 21'h1ffdfe; 
        10'b1011000001: data <= 21'h00074e; 
        10'b1011000010: data <= 21'h000afe; 
        10'b1011000011: data <= 21'h000625; 
        10'b1011000100: data <= 21'h000ecf; 
        10'b1011000101: data <= 21'h000efa; 
        10'b1011000110: data <= 21'h001bfe; 
        10'b1011000111: data <= 21'h001fff; 
        10'b1011001000: data <= 21'h00225a; 
        10'b1011001001: data <= 21'h001ae6; 
        10'b1011001010: data <= 21'h00131f; 
        10'b1011001011: data <= 21'h0007ae; 
        10'b1011001100: data <= 21'h1ffcea; 
        10'b1011001101: data <= 21'h1ff3e2; 
        10'b1011001110: data <= 21'h1ff3d2; 
        10'b1011001111: data <= 21'h1ff605; 
        10'b1011010000: data <= 21'h1ff618; 
        10'b1011010001: data <= 21'h1ffb03; 
        10'b1011010010: data <= 21'h1ffb02; 
        10'b1011010011: data <= 21'h1fff76; 
        10'b1011010100: data <= 21'h1ff9f2; 
        10'b1011010101: data <= 21'h0000c5; 
        10'b1011010110: data <= 21'h1ff80f; 
        10'b1011010111: data <= 21'h1ffee2; 
        10'b1011011000: data <= 21'h1ffa41; 
        10'b1011011001: data <= 21'h1ff7d1; 
        10'b1011011010: data <= 21'h1ff832; 
        10'b1011011011: data <= 21'h1ffe00; 
        10'b1011011100: data <= 21'h1ffe1d; 
        10'b1011011101: data <= 21'h1ffa9b; 
        10'b1011011110: data <= 21'h1ff9b8; 
        10'b1011011111: data <= 21'h1ffdd2; 
        10'b1011100000: data <= 21'h1ffe01; 
        10'b1011100001: data <= 21'h1ffd61; 
        10'b1011100010: data <= 21'h1ffc55; 
        10'b1011100011: data <= 21'h1ffcf0; 
        10'b1011100100: data <= 21'h1ffb75; 
        10'b1011100101: data <= 21'h1ffd8d; 
        10'b1011100110: data <= 21'h1ffb6a; 
        10'b1011100111: data <= 21'h1ff726; 
        10'b1011101000: data <= 21'h1ffa92; 
        10'b1011101001: data <= 21'h1ffd6c; 
        10'b1011101010: data <= 21'h1ffc70; 
        10'b1011101011: data <= 21'h1ffdae; 
        10'b1011101100: data <= 21'h1ff85b; 
        10'b1011101101: data <= 21'h1ff87e; 
        10'b1011101110: data <= 21'h1ffedb; 
        10'b1011101111: data <= 21'h1ffba2; 
        10'b1011110000: data <= 21'h000034; 
        10'b1011110001: data <= 21'h1ffa1f; 
        10'b1011110010: data <= 21'h1fff5b; 
        10'b1011110011: data <= 21'h0000e9; 
        10'b1011110100: data <= 21'h1ffc18; 
        10'b1011110101: data <= 21'h1ff9e3; 
        10'b1011110110: data <= 21'h1ffd4d; 
        10'b1011110111: data <= 21'h1ff855; 
        10'b1011111000: data <= 21'h000065; 
        10'b1011111001: data <= 21'h1ffdea; 
        10'b1011111010: data <= 21'h1fff9b; 
        10'b1011111011: data <= 21'h1ffd90; 
        10'b1011111100: data <= 21'h1ffec0; 
        10'b1011111101: data <= 21'h1ff83c; 
        10'b1011111110: data <= 21'h1ff9a2; 
        10'b1011111111: data <= 21'h1ffe53; 
        10'b1100000000: data <= 21'h1ff999; 
        10'b1100000001: data <= 21'h1ffecd; 
        10'b1100000010: data <= 21'h1ffb3a; 
        10'b1100000011: data <= 21'h1ffd31; 
        10'b1100000100: data <= 21'h1ffb71; 
        10'b1100000101: data <= 21'h1fffda; 
        10'b1100000110: data <= 21'h1ff8a8; 
        10'b1100000111: data <= 21'h1ff9ee; 
        10'b1100001000: data <= 21'h1fff7d; 
        10'b1100001001: data <= 21'h1ffd57; 
        10'b1100001010: data <= 21'h1ff9df; 
        10'b1100001011: data <= 21'h1ffe18; 
        10'b1100001100: data <= 21'h1ff8c3; 
        10'b1100001101: data <= 21'h1ff826; 
        10'b1100001110: data <= 21'h1fff8e; 
        10'b1100001111: data <= 21'h1ffc59; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 16) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 22'h3ffaf6; 
        10'b0000000001: data <= 22'h3ff38a; 
        10'b0000000010: data <= 22'h3fff62; 
        10'b0000000011: data <= 22'h000090; 
        10'b0000000100: data <= 22'h000141; 
        10'b0000000101: data <= 22'h3ffee8; 
        10'b0000000110: data <= 22'h3ffb43; 
        10'b0000000111: data <= 22'h00014c; 
        10'b0000001000: data <= 22'h3ff5f1; 
        10'b0000001001: data <= 22'h0000cb; 
        10'b0000001010: data <= 22'h0000d9; 
        10'b0000001011: data <= 22'h3ff76d; 
        10'b0000001100: data <= 22'h3ff738; 
        10'b0000001101: data <= 22'h3ff700; 
        10'b0000001110: data <= 22'h3ff7ad; 
        10'b0000001111: data <= 22'h3ff8c3; 
        10'b0000010000: data <= 22'h00002c; 
        10'b0000010001: data <= 22'h00008e; 
        10'b0000010010: data <= 22'h3ff391; 
        10'b0000010011: data <= 22'h000145; 
        10'b0000010100: data <= 22'h3ffbf6; 
        10'b0000010101: data <= 22'h3ffc81; 
        10'b0000010110: data <= 22'h3fefac; 
        10'b0000010111: data <= 22'h3fff1a; 
        10'b0000011000: data <= 22'h3fff64; 
        10'b0000011001: data <= 22'h3ff0a5; 
        10'b0000011010: data <= 22'h3ff871; 
        10'b0000011011: data <= 22'h000073; 
        10'b0000011100: data <= 22'h3ff327; 
        10'b0000011101: data <= 22'h3ff7f3; 
        10'b0000011110: data <= 22'h3ff35d; 
        10'b0000011111: data <= 22'h3ffb9a; 
        10'b0000100000: data <= 22'h3ff181; 
        10'b0000100001: data <= 22'h3ff911; 
        10'b0000100010: data <= 22'h0001aa; 
        10'b0000100011: data <= 22'h0000ec; 
        10'b0000100100: data <= 22'h3ff08f; 
        10'b0000100101: data <= 22'h3fefda; 
        10'b0000100110: data <= 22'h3ff17c; 
        10'b0000100111: data <= 22'h3ffb3c; 
        10'b0000101000: data <= 22'h3ffc8f; 
        10'b0000101001: data <= 22'h3ff89d; 
        10'b0000101010: data <= 22'h3ff75f; 
        10'b0000101011: data <= 22'h3ff463; 
        10'b0000101100: data <= 22'h000197; 
        10'b0000101101: data <= 22'h3ff398; 
        10'b0000101110: data <= 22'h3ffd3f; 
        10'b0000101111: data <= 22'h3ff68b; 
        10'b0000110000: data <= 22'h3ff6bd; 
        10'b0000110001: data <= 22'h3ff0fd; 
        10'b0000110010: data <= 22'h3ff9bd; 
        10'b0000110011: data <= 22'h3ffe83; 
        10'b0000110100: data <= 22'h3ff271; 
        10'b0000110101: data <= 22'h3fff37; 
        10'b0000110110: data <= 22'h3ffaa4; 
        10'b0000110111: data <= 22'h3ff291; 
        10'b0000111000: data <= 22'h3ff4b2; 
        10'b0000111001: data <= 22'h3ff9aa; 
        10'b0000111010: data <= 22'h3ff93a; 
        10'b0000111011: data <= 22'h3ff39b; 
        10'b0000111100: data <= 22'h3ffc0d; 
        10'b0000111101: data <= 22'h3ffd57; 
        10'b0000111110: data <= 22'h3ff570; 
        10'b0000111111: data <= 22'h3ffd21; 
        10'b0001000000: data <= 22'h3ffe9a; 
        10'b0001000001: data <= 22'h3ff89e; 
        10'b0001000010: data <= 22'h3ff232; 
        10'b0001000011: data <= 22'h3ff291; 
        10'b0001000100: data <= 22'h3ff0e0; 
        10'b0001000101: data <= 22'h3ff2e1; 
        10'b0001000110: data <= 22'h3ff7b2; 
        10'b0001000111: data <= 22'h3ff680; 
        10'b0001001000: data <= 22'h3ff541; 
        10'b0001001001: data <= 22'h3ff4dd; 
        10'b0001001010: data <= 22'h3ffd23; 
        10'b0001001011: data <= 22'h3fffac; 
        10'b0001001100: data <= 22'h3ff84a; 
        10'b0001001101: data <= 22'h3ff348; 
        10'b0001001110: data <= 22'h000166; 
        10'b0001001111: data <= 22'h3ffef5; 
        10'b0001010000: data <= 22'h00000a; 
        10'b0001010001: data <= 22'h3ff613; 
        10'b0001010010: data <= 22'h3ff050; 
        10'b0001010011: data <= 22'h3ff8b4; 
        10'b0001010100: data <= 22'h0001bc; 
        10'b0001010101: data <= 22'h3ffd02; 
        10'b0001010110: data <= 22'h3ff8e6; 
        10'b0001010111: data <= 22'h3ffe18; 
        10'b0001011000: data <= 22'h3ffcd2; 
        10'b0001011001: data <= 22'h000011; 
        10'b0001011010: data <= 22'h3ffb50; 
        10'b0001011011: data <= 22'h3fff1e; 
        10'b0001011100: data <= 22'h3ffe30; 
        10'b0001011101: data <= 22'h3ffa05; 
        10'b0001011110: data <= 22'h00058f; 
        10'b0001011111: data <= 22'h001286; 
        10'b0001100000: data <= 22'h00271d; 
        10'b0001100001: data <= 22'h00207e; 
        10'b0001100010: data <= 22'h00211e; 
        10'b0001100011: data <= 22'h00248f; 
        10'b0001100100: data <= 22'h00195a; 
        10'b0001100101: data <= 22'h001c95; 
        10'b0001100110: data <= 22'h001654; 
        10'b0001100111: data <= 22'h0001ac; 
        10'b0001101000: data <= 22'h3ffdc7; 
        10'b0001101001: data <= 22'h3fe4b9; 
        10'b0001101010: data <= 22'h3ff03a; 
        10'b0001101011: data <= 22'h3ffea4; 
        10'b0001101100: data <= 22'h0000c4; 
        10'b0001101101: data <= 22'h3ff407; 
        10'b0001101110: data <= 22'h3ffa8d; 
        10'b0001101111: data <= 22'h3ff57f; 
        10'b0001110000: data <= 22'h3ffa62; 
        10'b0001110001: data <= 22'h3fff17; 
        10'b0001110010: data <= 22'h3ffbc0; 
        10'b0001110011: data <= 22'h000079; 
        10'b0001110100: data <= 22'h0005f2; 
        10'b0001110101: data <= 22'h3ffff3; 
        10'b0001110110: data <= 22'h0016fa; 
        10'b0001110111: data <= 22'h001365; 
        10'b0001111000: data <= 22'h0034e3; 
        10'b0001111001: data <= 22'h002d70; 
        10'b0001111010: data <= 22'h003856; 
        10'b0001111011: data <= 22'h0043c5; 
        10'b0001111100: data <= 22'h004ea0; 
        10'b0001111101: data <= 22'h005444; 
        10'b0001111110: data <= 22'h004bc3; 
        10'b0001111111: data <= 22'h00378b; 
        10'b0010000000: data <= 22'h001f52; 
        10'b0010000001: data <= 22'h001910; 
        10'b0010000010: data <= 22'h0028f5; 
        10'b0010000011: data <= 22'h000507; 
        10'b0010000100: data <= 22'h3fe3f4; 
        10'b0010000101: data <= 22'h3fd443; 
        10'b0010000110: data <= 22'h3fda9f; 
        10'b0010000111: data <= 22'h3fdb6c; 
        10'b0010001000: data <= 22'h3ffb8e; 
        10'b0010001001: data <= 22'h3ff959; 
        10'b0010001010: data <= 22'h3ff677; 
        10'b0010001011: data <= 22'h3ffd81; 
        10'b0010001100: data <= 22'h3ff236; 
        10'b0010001101: data <= 22'h3ff036; 
        10'b0010001110: data <= 22'h3ff435; 
        10'b0010001111: data <= 22'h3ff439; 
        10'b0010010000: data <= 22'h0002f4; 
        10'b0010010001: data <= 22'h0017e4; 
        10'b0010010010: data <= 22'h002bac; 
        10'b0010010011: data <= 22'h0022e5; 
        10'b0010010100: data <= 22'h0027f1; 
        10'b0010010101: data <= 22'h00233e; 
        10'b0010010110: data <= 22'h001fe6; 
        10'b0010010111: data <= 22'h002988; 
        10'b0010011000: data <= 22'h002a2a; 
        10'b0010011001: data <= 22'h003295; 
        10'b0010011010: data <= 22'h0008a5; 
        10'b0010011011: data <= 22'h0021b2; 
        10'b0010011100: data <= 22'h0026e9; 
        10'b0010011101: data <= 22'h3ffd02; 
        10'b0010011110: data <= 22'h3ffdec; 
        10'b0010011111: data <= 22'h3fee5c; 
        10'b0010100000: data <= 22'h3fe77b; 
        10'b0010100001: data <= 22'h3fcbf3; 
        10'b0010100010: data <= 22'h3fbd6e; 
        10'b0010100011: data <= 22'h3fc7a8; 
        10'b0010100100: data <= 22'h3fefab; 
        10'b0010100101: data <= 22'h000012; 
        10'b0010100110: data <= 22'h3ff4c5; 
        10'b0010100111: data <= 22'h3ff91b; 
        10'b0010101000: data <= 22'h3ff3a1; 
        10'b0010101001: data <= 22'h3ff647; 
        10'b0010101010: data <= 22'h3ff538; 
        10'b0010101011: data <= 22'h000509; 
        10'b0010101100: data <= 22'h001d95; 
        10'b0010101101: data <= 22'h003700; 
        10'b0010101110: data <= 22'h002a10; 
        10'b0010101111: data <= 22'h00203b; 
        10'b0010110000: data <= 22'h0030d0; 
        10'b0010110001: data <= 22'h0027d3; 
        10'b0010110010: data <= 22'h002365; 
        10'b0010110011: data <= 22'h0021dd; 
        10'b0010110100: data <= 22'h002d4a; 
        10'b0010110101: data <= 22'h0040f7; 
        10'b0010110110: data <= 22'h002d2a; 
        10'b0010110111: data <= 22'h00104f; 
        10'b0010111000: data <= 22'h002afa; 
        10'b0010111001: data <= 22'h002767; 
        10'b0010111010: data <= 22'h002582; 
        10'b0010111011: data <= 22'h3fef3a; 
        10'b0010111100: data <= 22'h001000; 
        10'b0010111101: data <= 22'h3ff024; 
        10'b0010111110: data <= 22'h3fc6df; 
        10'b0010111111: data <= 22'h3fc6de; 
        10'b0011000000: data <= 22'h3fdd02; 
        10'b0011000001: data <= 22'h3ff8f6; 
        10'b0011000010: data <= 22'h3ffe71; 
        10'b0011000011: data <= 22'h3ffa80; 
        10'b0011000100: data <= 22'h0000ac; 
        10'b0011000101: data <= 22'h3ffe12; 
        10'b0011000110: data <= 22'h00035b; 
        10'b0011000111: data <= 22'h0018b1; 
        10'b0011001000: data <= 22'h0040f0; 
        10'b0011001001: data <= 22'h004099; 
        10'b0011001010: data <= 22'h002d85; 
        10'b0011001011: data <= 22'h000ccc; 
        10'b0011001100: data <= 22'h000db8; 
        10'b0011001101: data <= 22'h001cf0; 
        10'b0011001110: data <= 22'h0008e1; 
        10'b0011001111: data <= 22'h000d30; 
        10'b0011010000: data <= 22'h002618; 
        10'b0011010001: data <= 22'h002413; 
        10'b0011010010: data <= 22'h003bc7; 
        10'b0011010011: data <= 22'h00231f; 
        10'b0011010100: data <= 22'h000ac3; 
        10'b0011010101: data <= 22'h001e01; 
        10'b0011010110: data <= 22'h0018df; 
        10'b0011010111: data <= 22'h001b05; 
        10'b0011011000: data <= 22'h001b63; 
        10'b0011011001: data <= 22'h0003df; 
        10'b0011011010: data <= 22'h3fe46a; 
        10'b0011011011: data <= 22'h3fbfe4; 
        10'b0011011100: data <= 22'h3fd207; 
        10'b0011011101: data <= 22'h3ff3ed; 
        10'b0011011110: data <= 22'h3ff047; 
        10'b0011011111: data <= 22'h3ff79d; 
        10'b0011100000: data <= 22'h3ff9e8; 
        10'b0011100001: data <= 22'h3ff696; 
        10'b0011100010: data <= 22'h0002ba; 
        10'b0011100011: data <= 22'h00170e; 
        10'b0011100100: data <= 22'h003588; 
        10'b0011100101: data <= 22'h0032dd; 
        10'b0011100110: data <= 22'h00263a; 
        10'b0011100111: data <= 22'h000f9d; 
        10'b0011101000: data <= 22'h0019e4; 
        10'b0011101001: data <= 22'h000c57; 
        10'b0011101010: data <= 22'h0020b4; 
        10'b0011101011: data <= 22'h000a7f; 
        10'b0011101100: data <= 22'h0008ef; 
        10'b0011101101: data <= 22'h000ffd; 
        10'b0011101110: data <= 22'h0040ff; 
        10'b0011101111: data <= 22'h0035ed; 
        10'b0011110000: data <= 22'h000c71; 
        10'b0011110001: data <= 22'h001df8; 
        10'b0011110010: data <= 22'h002b11; 
        10'b0011110011: data <= 22'h001c11; 
        10'b0011110100: data <= 22'h002913; 
        10'b0011110101: data <= 22'h001526; 
        10'b0011110110: data <= 22'h3ff501; 
        10'b0011110111: data <= 22'h3fc495; 
        10'b0011111000: data <= 22'h3fd383; 
        10'b0011111001: data <= 22'h3fefc4; 
        10'b0011111010: data <= 22'h3ff231; 
        10'b0011111011: data <= 22'h3ff612; 
        10'b0011111100: data <= 22'h3ff835; 
        10'b0011111101: data <= 22'h3ff0bc; 
        10'b0011111110: data <= 22'h3ffb21; 
        10'b0011111111: data <= 22'h0009f0; 
        10'b0100000000: data <= 22'h001ba9; 
        10'b0100000001: data <= 22'h0024b3; 
        10'b0100000010: data <= 22'h001e64; 
        10'b0100000011: data <= 22'h000762; 
        10'b0100000100: data <= 22'h3ffc25; 
        10'b0100000101: data <= 22'h3fe3a7; 
        10'b0100000110: data <= 22'h3fc9f5; 
        10'b0100000111: data <= 22'h3f9cc2; 
        10'b0100001000: data <= 22'h3faf79; 
        10'b0100001001: data <= 22'h3ff546; 
        10'b0100001010: data <= 22'h004d6b; 
        10'b0100001011: data <= 22'h0076ff; 
        10'b0100001100: data <= 22'h0044be; 
        10'b0100001101: data <= 22'h002833; 
        10'b0100001110: data <= 22'h002bb1; 
        10'b0100001111: data <= 22'h002862; 
        10'b0100010000: data <= 22'h003c7d; 
        10'b0100010001: data <= 22'h00269a; 
        10'b0100010010: data <= 22'h3ff44e; 
        10'b0100010011: data <= 22'h3fc4fd; 
        10'b0100010100: data <= 22'h3fe24e; 
        10'b0100010101: data <= 22'h3fef41; 
        10'b0100010110: data <= 22'h3ff368; 
        10'b0100010111: data <= 22'h3ff57e; 
        10'b0100011000: data <= 22'h3ffe50; 
        10'b0100011001: data <= 22'h3ffd7c; 
        10'b0100011010: data <= 22'h0000d4; 
        10'b0100011011: data <= 22'h000eea; 
        10'b0100011100: data <= 22'h000d69; 
        10'b0100011101: data <= 22'h0005b5; 
        10'b0100011110: data <= 22'h3feeb4; 
        10'b0100011111: data <= 22'h3fd42d; 
        10'b0100100000: data <= 22'h3fafd8; 
        10'b0100100001: data <= 22'h3f8d6b; 
        10'b0100100010: data <= 22'h3f7396; 
        10'b0100100011: data <= 22'h3f6ffd; 
        10'b0100100100: data <= 22'h3f95ea; 
        10'b0100100101: data <= 22'h3fe53a; 
        10'b0100100110: data <= 22'h003f7a; 
        10'b0100100111: data <= 22'h004961; 
        10'b0100101000: data <= 22'h003e79; 
        10'b0100101001: data <= 22'h003a3f; 
        10'b0100101010: data <= 22'h0023f4; 
        10'b0100101011: data <= 22'h003e5e; 
        10'b0100101100: data <= 22'h0039e3; 
        10'b0100101101: data <= 22'h001731; 
        10'b0100101110: data <= 22'h3feb3f; 
        10'b0100101111: data <= 22'h3fd9b8; 
        10'b0100110000: data <= 22'h3ff1b0; 
        10'b0100110001: data <= 22'h3fefcb; 
        10'b0100110010: data <= 22'h3ff924; 
        10'b0100110011: data <= 22'h3ffe41; 
        10'b0100110100: data <= 22'h0001e3; 
        10'b0100110101: data <= 22'h3ffe43; 
        10'b0100110110: data <= 22'h3ff2bd; 
        10'b0100110111: data <= 22'h000e87; 
        10'b0100111000: data <= 22'h3ff768; 
        10'b0100111001: data <= 22'h3fd312; 
        10'b0100111010: data <= 22'h3fbc9a; 
        10'b0100111011: data <= 22'h3f9ced; 
        10'b0100111100: data <= 22'h3f8425; 
        10'b0100111101: data <= 22'h3f94f9; 
        10'b0100111110: data <= 22'h3fae83; 
        10'b0100111111: data <= 22'h3fd995; 
        10'b0101000000: data <= 22'h3feb31; 
        10'b0101000001: data <= 22'h001ae6; 
        10'b0101000010: data <= 22'h002a3e; 
        10'b0101000011: data <= 22'h002a77; 
        10'b0101000100: data <= 22'h001362; 
        10'b0101000101: data <= 22'h002bfb; 
        10'b0101000110: data <= 22'h00366b; 
        10'b0101000111: data <= 22'h003510; 
        10'b0101001000: data <= 22'h002e52; 
        10'b0101001001: data <= 22'h000038; 
        10'b0101001010: data <= 22'h3feb9b; 
        10'b0101001011: data <= 22'h3feeef; 
        10'b0101001100: data <= 22'h3ff0f9; 
        10'b0101001101: data <= 22'h3ff71a; 
        10'b0101001110: data <= 22'h3ff3ae; 
        10'b0101001111: data <= 22'h3ff233; 
        10'b0101010000: data <= 22'h000088; 
        10'b0101010001: data <= 22'h3ff598; 
        10'b0101010010: data <= 22'h3ffd59; 
        10'b0101010011: data <= 22'h3fff31; 
        10'b0101010100: data <= 22'h3fefab; 
        10'b0101010101: data <= 22'h3fd2e7; 
        10'b0101010110: data <= 22'h3fb10b; 
        10'b0101010111: data <= 22'h3f9d38; 
        10'b0101011000: data <= 22'h3fa6ad; 
        10'b0101011001: data <= 22'h3fd06d; 
        10'b0101011010: data <= 22'h0000f0; 
        10'b0101011011: data <= 22'h0007ee; 
        10'b0101011100: data <= 22'h000c92; 
        10'b0101011101: data <= 22'h001c89; 
        10'b0101011110: data <= 22'h0046b3; 
        10'b0101011111: data <= 22'h002488; 
        10'b0101100000: data <= 22'h0018f3; 
        10'b0101100001: data <= 22'h00234d; 
        10'b0101100010: data <= 22'h001c48; 
        10'b0101100011: data <= 22'h3ffd88; 
        10'b0101100100: data <= 22'h3fdb65; 
        10'b0101100101: data <= 22'h3fcdbc; 
        10'b0101100110: data <= 22'h3fcb62; 
        10'b0101100111: data <= 22'h3fde8c; 
        10'b0101101000: data <= 22'h3ffa20; 
        10'b0101101001: data <= 22'h3ff5dc; 
        10'b0101101010: data <= 22'h3ffa88; 
        10'b0101101011: data <= 22'h3ffc26; 
        10'b0101101100: data <= 22'h3ff8de; 
        10'b0101101101: data <= 22'h3ff530; 
        10'b0101101110: data <= 22'h3ff95c; 
        10'b0101101111: data <= 22'h3ffb8e; 
        10'b0101110000: data <= 22'h3feb1c; 
        10'b0101110001: data <= 22'h3fe12b; 
        10'b0101110010: data <= 22'h3fbfc8; 
        10'b0101110011: data <= 22'h3fb5dd; 
        10'b0101110100: data <= 22'h3fcdb6; 
        10'b0101110101: data <= 22'h3ff61a; 
        10'b0101110110: data <= 22'h3fefa8; 
        10'b0101110111: data <= 22'h3fd560; 
        10'b0101111000: data <= 22'h000364; 
        10'b0101111001: data <= 22'h003cdb; 
        10'b0101111010: data <= 22'h003d78; 
        10'b0101111011: data <= 22'h000b38; 
        10'b0101111100: data <= 22'h001be7; 
        10'b0101111101: data <= 22'h001dc0; 
        10'b0101111110: data <= 22'h000fca; 
        10'b0101111111: data <= 22'h3feb0f; 
        10'b0110000000: data <= 22'h3fc7e5; 
        10'b0110000001: data <= 22'h3fc79e; 
        10'b0110000010: data <= 22'h3fd378; 
        10'b0110000011: data <= 22'h3fe0b9; 
        10'b0110000100: data <= 22'h3fee0a; 
        10'b0110000101: data <= 22'h3fff9e; 
        10'b0110000110: data <= 22'h3ffcba; 
        10'b0110000111: data <= 22'h3ff671; 
        10'b0110001000: data <= 22'h00017c; 
        10'b0110001001: data <= 22'h3ff3cb; 
        10'b0110001010: data <= 22'h3ff830; 
        10'b0110001011: data <= 22'h3ffaea; 
        10'b0110001100: data <= 22'h3ffc22; 
        10'b0110001101: data <= 22'h3fe637; 
        10'b0110001110: data <= 22'h3fc60d; 
        10'b0110001111: data <= 22'h3fcb9f; 
        10'b0110010000: data <= 22'h3fdc6e; 
        10'b0110010001: data <= 22'h3ffb0f; 
        10'b0110010010: data <= 22'h3fdab3; 
        10'b0110010011: data <= 22'h3fd83b; 
        10'b0110010100: data <= 22'h000b45; 
        10'b0110010101: data <= 22'h001d72; 
        10'b0110010110: data <= 22'h001f70; 
        10'b0110010111: data <= 22'h3ffb54; 
        10'b0110011000: data <= 22'h3ff339; 
        10'b0110011001: data <= 22'h3ff67c; 
        10'b0110011010: data <= 22'h00044b; 
        10'b0110011011: data <= 22'h3fe79a; 
        10'b0110011100: data <= 22'h3fdef9; 
        10'b0110011101: data <= 22'h3fefff; 
        10'b0110011110: data <= 22'h3fe946; 
        10'b0110011111: data <= 22'h3ff0a8; 
        10'b0110100000: data <= 22'h3febcd; 
        10'b0110100001: data <= 22'h3fedd7; 
        10'b0110100010: data <= 22'h000074; 
        10'b0110100011: data <= 22'h0000e7; 
        10'b0110100100: data <= 22'h000154; 
        10'b0110100101: data <= 22'h3ff3fb; 
        10'b0110100110: data <= 22'h0001cf; 
        10'b0110100111: data <= 22'h000472; 
        10'b0110101000: data <= 22'h3ffad1; 
        10'b0110101001: data <= 22'h3fe308; 
        10'b0110101010: data <= 22'h3fca3e; 
        10'b0110101011: data <= 22'h3fc679; 
        10'b0110101100: data <= 22'h3fd4f6; 
        10'b0110101101: data <= 22'h3fe6c4; 
        10'b0110101110: data <= 22'h3fe40d; 
        10'b0110101111: data <= 22'h3ff68f; 
        10'b0110110000: data <= 22'h000b9e; 
        10'b0110110001: data <= 22'h002fdd; 
        10'b0110110010: data <= 22'h001b7b; 
        10'b0110110011: data <= 22'h3ffd4a; 
        10'b0110110100: data <= 22'h3fd80c; 
        10'b0110110101: data <= 22'h3ff466; 
        10'b0110110110: data <= 22'h3ffc10; 
        10'b0110110111: data <= 22'h000a83; 
        10'b0110111000: data <= 22'h0018cf; 
        10'b0110111001: data <= 22'h00183a; 
        10'b0110111010: data <= 22'h00085f; 
        10'b0110111011: data <= 22'h00032e; 
        10'b0110111100: data <= 22'h3ff0d7; 
        10'b0110111101: data <= 22'h3ffc99; 
        10'b0110111110: data <= 22'h3ffb33; 
        10'b0110111111: data <= 22'h3ff3ef; 
        10'b0111000000: data <= 22'h3ffb76; 
        10'b0111000001: data <= 22'h3ffd6f; 
        10'b0111000010: data <= 22'h000b06; 
        10'b0111000011: data <= 22'h0001f5; 
        10'b0111000100: data <= 22'h000814; 
        10'b0111000101: data <= 22'h3ff29f; 
        10'b0111000110: data <= 22'h3fea09; 
        10'b0111000111: data <= 22'h3fd9f9; 
        10'b0111001000: data <= 22'h3fad3e; 
        10'b0111001001: data <= 22'h3fa8ca; 
        10'b0111001010: data <= 22'h3fb2b5; 
        10'b0111001011: data <= 22'h3fec6c; 
        10'b0111001100: data <= 22'h00170f; 
        10'b0111001101: data <= 22'h003bb4; 
        10'b0111001110: data <= 22'h3ff98c; 
        10'b0111001111: data <= 22'h3fd46f; 
        10'b0111010000: data <= 22'h3fd1eb; 
        10'b0111010001: data <= 22'h3ff0ff; 
        10'b0111010010: data <= 22'h001370; 
        10'b0111010011: data <= 22'h0032ec; 
        10'b0111010100: data <= 22'h0023d6; 
        10'b0111010101: data <= 22'h002d1a; 
        10'b0111010110: data <= 22'h002bce; 
        10'b0111010111: data <= 22'h001365; 
        10'b0111011000: data <= 22'h3ffa44; 
        10'b0111011001: data <= 22'h3ffc21; 
        10'b0111011010: data <= 22'h3fff78; 
        10'b0111011011: data <= 22'h3ffe90; 
        10'b0111011100: data <= 22'h3ffe3c; 
        10'b0111011101: data <= 22'h0001de; 
        10'b0111011110: data <= 22'h00003d; 
        10'b0111011111: data <= 22'h001be7; 
        10'b0111100000: data <= 22'h000f6c; 
        10'b0111100001: data <= 22'h0004d3; 
        10'b0111100010: data <= 22'h3ff13b; 
        10'b0111100011: data <= 22'h3fcdc8; 
        10'b0111100100: data <= 22'h3fa694; 
        10'b0111100101: data <= 22'h3f7236; 
        10'b0111100110: data <= 22'h3f4f8b; 
        10'b0111100111: data <= 22'h3f5ef0; 
        10'b0111101000: data <= 22'h3f85b8; 
        10'b0111101001: data <= 22'h3fba55; 
        10'b0111101010: data <= 22'h3fbf58; 
        10'b0111101011: data <= 22'h3fc64b; 
        10'b0111101100: data <= 22'h3ffdb5; 
        10'b0111101101: data <= 22'h0011cf; 
        10'b0111101110: data <= 22'h0020a0; 
        10'b0111101111: data <= 22'h0033a5; 
        10'b0111110000: data <= 22'h000ab3; 
        10'b0111110001: data <= 22'h003e7e; 
        10'b0111110010: data <= 22'h003e62; 
        10'b0111110011: data <= 22'h0012c7; 
        10'b0111110100: data <= 22'h3ff6c5; 
        10'b0111110101: data <= 22'h3ff2b6; 
        10'b0111110110: data <= 22'h3ff3e3; 
        10'b0111110111: data <= 22'h3ff4ee; 
        10'b0111111000: data <= 22'h3ff929; 
        10'b0111111001: data <= 22'h3ff996; 
        10'b0111111010: data <= 22'h00056b; 
        10'b0111111011: data <= 22'h002947; 
        10'b0111111100: data <= 22'h001db8; 
        10'b0111111101: data <= 22'h0011ec; 
        10'b0111111110: data <= 22'h000964; 
        10'b0111111111: data <= 22'h3ff51b; 
        10'b1000000000: data <= 22'h3fe035; 
        10'b1000000001: data <= 22'h3f9833; 
        10'b1000000010: data <= 22'h3f671d; 
        10'b1000000011: data <= 22'h3f6f5a; 
        10'b1000000100: data <= 22'h3f5155; 
        10'b1000000101: data <= 22'h3f7170; 
        10'b1000000110: data <= 22'h3fa5d1; 
        10'b1000000111: data <= 22'h3feb7d; 
        10'b1000001000: data <= 22'h002468; 
        10'b1000001001: data <= 22'h003113; 
        10'b1000001010: data <= 22'h0034e3; 
        10'b1000001011: data <= 22'h003449; 
        10'b1000001100: data <= 22'h00249c; 
        10'b1000001101: data <= 22'h0048fa; 
        10'b1000001110: data <= 22'h00441c; 
        10'b1000001111: data <= 22'h001a06; 
        10'b1000010000: data <= 22'h3fe807; 
        10'b1000010001: data <= 22'h3fefc5; 
        10'b1000010010: data <= 22'h3ff430; 
        10'b1000010011: data <= 22'h3ffe1e; 
        10'b1000010100: data <= 22'h3ffe22; 
        10'b1000010101: data <= 22'h3ff411; 
        10'b1000010110: data <= 22'h3ff85a; 
        10'b1000010111: data <= 22'h0033c0; 
        10'b1000011000: data <= 22'h0034c9; 
        10'b1000011001: data <= 22'h003e02; 
        10'b1000011010: data <= 22'h00356f; 
        10'b1000011011: data <= 22'h00139c; 
        10'b1000011100: data <= 22'h0005e3; 
        10'b1000011101: data <= 22'h3fea35; 
        10'b1000011110: data <= 22'h3ff049; 
        10'b1000011111: data <= 22'h3fcebb; 
        10'b1000100000: data <= 22'h3fb803; 
        10'b1000100001: data <= 22'h3fb36f; 
        10'b1000100010: data <= 22'h3fcbd4; 
        10'b1000100011: data <= 22'h001261; 
        10'b1000100100: data <= 22'h003145; 
        10'b1000100101: data <= 22'h003d98; 
        10'b1000100110: data <= 22'h004508; 
        10'b1000100111: data <= 22'h003dbd; 
        10'b1000101000: data <= 22'h0036a7; 
        10'b1000101001: data <= 22'h003fc1; 
        10'b1000101010: data <= 22'h00186f; 
        10'b1000101011: data <= 22'h0002d9; 
        10'b1000101100: data <= 22'h3febbb; 
        10'b1000101101: data <= 22'h3ffc41; 
        10'b1000101110: data <= 22'h3ffdfb; 
        10'b1000101111: data <= 22'h3ffbab; 
        10'b1000110000: data <= 22'h3ffd62; 
        10'b1000110001: data <= 22'h3ff041; 
        10'b1000110010: data <= 22'h000950; 
        10'b1000110011: data <= 22'h003789; 
        10'b1000110100: data <= 22'h004441; 
        10'b1000110101: data <= 22'h0049e2; 
        10'b1000110110: data <= 22'h004e3f; 
        10'b1000110111: data <= 22'h00277b; 
        10'b1000111000: data <= 22'h002e74; 
        10'b1000111001: data <= 22'h003491; 
        10'b1000111010: data <= 22'h001367; 
        10'b1000111011: data <= 22'h3ffab4; 
        10'b1000111100: data <= 22'h3fee5b; 
        10'b1000111101: data <= 22'h3fe4fb; 
        10'b1000111110: data <= 22'h00082c; 
        10'b1000111111: data <= 22'h000e8f; 
        10'b1001000000: data <= 22'h001bc9; 
        10'b1001000001: data <= 22'h003185; 
        10'b1001000010: data <= 22'h0033dd; 
        10'b1001000011: data <= 22'h00234c; 
        10'b1001000100: data <= 22'h003d77; 
        10'b1001000101: data <= 22'h0022ed; 
        10'b1001000110: data <= 22'h3ff97d; 
        10'b1001000111: data <= 22'h3ff201; 
        10'b1001001000: data <= 22'h3fefc0; 
        10'b1001001001: data <= 22'h3ffb34; 
        10'b1001001010: data <= 22'h3ffafe; 
        10'b1001001011: data <= 22'h3ffa6a; 
        10'b1001001100: data <= 22'h3ff568; 
        10'b1001001101: data <= 22'h3fff47; 
        10'b1001001110: data <= 22'h3ffc27; 
        10'b1001001111: data <= 22'h001b9c; 
        10'b1001010000: data <= 22'h0041e8; 
        10'b1001010001: data <= 22'h0041d1; 
        10'b1001010010: data <= 22'h00397d; 
        10'b1001010011: data <= 22'h00206e; 
        10'b1001010100: data <= 22'h00229a; 
        10'b1001010101: data <= 22'h000b71; 
        10'b1001010110: data <= 22'h3ffb72; 
        10'b1001010111: data <= 22'h3ff071; 
        10'b1001011000: data <= 22'h0004fd; 
        10'b1001011001: data <= 22'h3ffd33; 
        10'b1001011010: data <= 22'h3ffbed; 
        10'b1001011011: data <= 22'h3ff868; 
        10'b1001011100: data <= 22'h001023; 
        10'b1001011101: data <= 22'h0005e4; 
        10'b1001011110: data <= 22'h001fa8; 
        10'b1001011111: data <= 22'h0032e6; 
        10'b1001100000: data <= 22'h001d9b; 
        10'b1001100001: data <= 22'h000b52; 
        10'b1001100010: data <= 22'h3ff488; 
        10'b1001100011: data <= 22'h3fe270; 
        10'b1001100100: data <= 22'h3ff664; 
        10'b1001100101: data <= 22'h3ff3ce; 
        10'b1001100110: data <= 22'h3fefef; 
        10'b1001100111: data <= 22'h3ff0f2; 
        10'b1001101000: data <= 22'h3ff95e; 
        10'b1001101001: data <= 22'h3ffb62; 
        10'b1001101010: data <= 22'h3ffced; 
        10'b1001101011: data <= 22'h00112b; 
        10'b1001101100: data <= 22'h002119; 
        10'b1001101101: data <= 22'h002d0d; 
        10'b1001101110: data <= 22'h002832; 
        10'b1001101111: data <= 22'h0016e4; 
        10'b1001110000: data <= 22'h0001c8; 
        10'b1001110001: data <= 22'h001090; 
        10'b1001110010: data <= 22'h001401; 
        10'b1001110011: data <= 22'h00184f; 
        10'b1001110100: data <= 22'h0006bb; 
        10'b1001110101: data <= 22'h3ff726; 
        10'b1001110110: data <= 22'h3ff694; 
        10'b1001110111: data <= 22'h3ff29a; 
        10'b1001111000: data <= 22'h000a7b; 
        10'b1001111001: data <= 22'h0007ff; 
        10'b1001111010: data <= 22'h0007dd; 
        10'b1001111011: data <= 22'h00232d; 
        10'b1001111100: data <= 22'h001111; 
        10'b1001111101: data <= 22'h3ff9f1; 
        10'b1001111110: data <= 22'h3ff820; 
        10'b1001111111: data <= 22'h3ff5b6; 
        10'b1010000000: data <= 22'h3fe963; 
        10'b1010000001: data <= 22'h3fef10; 
        10'b1010000010: data <= 22'h3ffced; 
        10'b1010000011: data <= 22'h3fff88; 
        10'b1010000100: data <= 22'h3ffb4b; 
        10'b1010000101: data <= 22'h3ff34c; 
        10'b1010000110: data <= 22'h3ff574; 
        10'b1010000111: data <= 22'h000b4e; 
        10'b1010001000: data <= 22'h002427; 
        10'b1010001001: data <= 22'h003698; 
        10'b1010001010: data <= 22'h0028ae; 
        10'b1010001011: data <= 22'h002af4; 
        10'b1010001100: data <= 22'h000a64; 
        10'b1010001101: data <= 22'h001b83; 
        10'b1010001110: data <= 22'h00117b; 
        10'b1010001111: data <= 22'h3fffba; 
        10'b1010010000: data <= 22'h3ff237; 
        10'b1010010001: data <= 22'h000234; 
        10'b1010010010: data <= 22'h000597; 
        10'b1010010011: data <= 22'h000dc3; 
        10'b1010010100: data <= 22'h000a3e; 
        10'b1010010101: data <= 22'h001545; 
        10'b1010010110: data <= 22'h0021dc; 
        10'b1010010111: data <= 22'h3ffa48; 
        10'b1010011000: data <= 22'h3fe95b; 
        10'b1010011001: data <= 22'h3fe996; 
        10'b1010011010: data <= 22'h3ff431; 
        10'b1010011011: data <= 22'h3ff136; 
        10'b1010011100: data <= 22'h3ffeb0; 
        10'b1010011101: data <= 22'h3ffc2c; 
        10'b1010011110: data <= 22'h3ff1f2; 
        10'b1010011111: data <= 22'h3ff329; 
        10'b1010100000: data <= 22'h3ff5e2; 
        10'b1010100001: data <= 22'h00019a; 
        10'b1010100010: data <= 22'h0001b3; 
        10'b1010100011: data <= 22'h000036; 
        10'b1010100100: data <= 22'h00173c; 
        10'b1010100101: data <= 22'h00256c; 
        10'b1010100110: data <= 22'h002c17; 
        10'b1010100111: data <= 22'h003407; 
        10'b1010101000: data <= 22'h0034db; 
        10'b1010101001: data <= 22'h002b5a; 
        10'b1010101010: data <= 22'h003f2d; 
        10'b1010101011: data <= 22'h0042b6; 
        10'b1010101100: data <= 22'h004455; 
        10'b1010101101: data <= 22'h0035d2; 
        10'b1010101110: data <= 22'h002f78; 
        10'b1010101111: data <= 22'h00231b; 
        10'b1010110000: data <= 22'h002184; 
        10'b1010110001: data <= 22'h3ffd17; 
        10'b1010110010: data <= 22'h3fe4c3; 
        10'b1010110011: data <= 22'h3fda50; 
        10'b1010110100: data <= 22'h3fde23; 
        10'b1010110101: data <= 22'h3feb56; 
        10'b1010110110: data <= 22'h3fecb2; 
        10'b1010110111: data <= 22'h3ffa4c; 
        10'b1010111000: data <= 22'h3ff667; 
        10'b1010111001: data <= 22'h3fffc0; 
        10'b1010111010: data <= 22'h3ff62f; 
        10'b1010111011: data <= 22'h0001c5; 
        10'b1010111100: data <= 22'h3ffe7f; 
        10'b1010111101: data <= 22'h3fefc9; 
        10'b1010111110: data <= 22'h00013f; 
        10'b1010111111: data <= 22'h00029f; 
        10'b1011000000: data <= 22'h3ffbfd; 
        10'b1011000001: data <= 22'h000e9c; 
        10'b1011000010: data <= 22'h0015fc; 
        10'b1011000011: data <= 22'h000c4a; 
        10'b1011000100: data <= 22'h001d9f; 
        10'b1011000101: data <= 22'h001df3; 
        10'b1011000110: data <= 22'h0037fd; 
        10'b1011000111: data <= 22'h003ffe; 
        10'b1011001000: data <= 22'h0044b4; 
        10'b1011001001: data <= 22'h0035cc; 
        10'b1011001010: data <= 22'h00263d; 
        10'b1011001011: data <= 22'h000f5d; 
        10'b1011001100: data <= 22'h3ff9d3; 
        10'b1011001101: data <= 22'h3fe7c4; 
        10'b1011001110: data <= 22'h3fe7a3; 
        10'b1011001111: data <= 22'h3fec0a; 
        10'b1011010000: data <= 22'h3fec31; 
        10'b1011010001: data <= 22'h3ff605; 
        10'b1011010010: data <= 22'h3ff604; 
        10'b1011010011: data <= 22'h3ffeeb; 
        10'b1011010100: data <= 22'h3ff3e3; 
        10'b1011010101: data <= 22'h00018a; 
        10'b1011010110: data <= 22'h3ff01e; 
        10'b1011010111: data <= 22'h3ffdc4; 
        10'b1011011000: data <= 22'h3ff482; 
        10'b1011011001: data <= 22'h3fefa3; 
        10'b1011011010: data <= 22'h3ff064; 
        10'b1011011011: data <= 22'h3ffc00; 
        10'b1011011100: data <= 22'h3ffc3a; 
        10'b1011011101: data <= 22'h3ff537; 
        10'b1011011110: data <= 22'h3ff371; 
        10'b1011011111: data <= 22'h3ffba5; 
        10'b1011100000: data <= 22'h3ffc02; 
        10'b1011100001: data <= 22'h3ffac2; 
        10'b1011100010: data <= 22'h3ff8a9; 
        10'b1011100011: data <= 22'h3ff9df; 
        10'b1011100100: data <= 22'h3ff6ea; 
        10'b1011100101: data <= 22'h3ffb1b; 
        10'b1011100110: data <= 22'h3ff6d4; 
        10'b1011100111: data <= 22'h3fee4d; 
        10'b1011101000: data <= 22'h3ff524; 
        10'b1011101001: data <= 22'h3ffad9; 
        10'b1011101010: data <= 22'h3ff8e0; 
        10'b1011101011: data <= 22'h3ffb5c; 
        10'b1011101100: data <= 22'h3ff0b7; 
        10'b1011101101: data <= 22'h3ff0fb; 
        10'b1011101110: data <= 22'h3ffdb5; 
        10'b1011101111: data <= 22'h3ff744; 
        10'b1011110000: data <= 22'h000067; 
        10'b1011110001: data <= 22'h3ff43d; 
        10'b1011110010: data <= 22'h3ffeb5; 
        10'b1011110011: data <= 22'h0001d2; 
        10'b1011110100: data <= 22'h3ff830; 
        10'b1011110101: data <= 22'h3ff3c6; 
        10'b1011110110: data <= 22'h3ffa9a; 
        10'b1011110111: data <= 22'h3ff0ab; 
        10'b1011111000: data <= 22'h0000ca; 
        10'b1011111001: data <= 22'h3ffbd4; 
        10'b1011111010: data <= 22'h3fff37; 
        10'b1011111011: data <= 22'h3ffb20; 
        10'b1011111100: data <= 22'h3ffd80; 
        10'b1011111101: data <= 22'h3ff078; 
        10'b1011111110: data <= 22'h3ff344; 
        10'b1011111111: data <= 22'h3ffca5; 
        10'b1100000000: data <= 22'h3ff333; 
        10'b1100000001: data <= 22'h3ffd99; 
        10'b1100000010: data <= 22'h3ff673; 
        10'b1100000011: data <= 22'h3ffa63; 
        10'b1100000100: data <= 22'h3ff6e3; 
        10'b1100000101: data <= 22'h3fffb4; 
        10'b1100000110: data <= 22'h3ff150; 
        10'b1100000111: data <= 22'h3ff3dd; 
        10'b1100001000: data <= 22'h3ffef9; 
        10'b1100001001: data <= 22'h3ffaaf; 
        10'b1100001010: data <= 22'h3ff3bf; 
        10'b1100001011: data <= 22'h3ffc31; 
        10'b1100001100: data <= 22'h3ff186; 
        10'b1100001101: data <= 22'h3ff04c; 
        10'b1100001110: data <= 22'h3fff1c; 
        10'b1100001111: data <= 22'h3ff8b3; 
      endcase 
    end 
  end 
endgenerate 
assign dout = data; 
endmodule
