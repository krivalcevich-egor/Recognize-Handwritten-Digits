`timescale 1ns / 1ps 
 
////////////////////////////////////////////////////////////////////////////////// 
// WEIGHT MEMORY (ROM) 
////////////////////////////////////////////////////////////////////////////////// 
module ROM_weights_9 #( 
    parameter int WGHT_INT = 6, // integer part 
    parameter int WGHT_FRC = 16 // fractional part 
)( 
    input logic clk, // clock 
    input logic [9:0] address,
    output [WGHT_INT + WGHT_FRC-1:0] dout 
); 

(* rom_style = "block" *) reg [WGHT_INT + WGHT_FRC-1:0] data;
generate 
  if (WGHT_FRC == 1) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 7'h00; 
        10'b0000000001: data <= 7'h00; 
        10'b0000000010: data <= 7'h00; 
        10'b0000000011: data <= 7'h00; 
        10'b0000000100: data <= 7'h00; 
        10'b0000000101: data <= 7'h00; 
        10'b0000000110: data <= 7'h00; 
        10'b0000000111: data <= 7'h00; 
        10'b0000001000: data <= 7'h00; 
        10'b0000001001: data <= 7'h00; 
        10'b0000001010: data <= 7'h00; 
        10'b0000001011: data <= 7'h00; 
        10'b0000001100: data <= 7'h00; 
        10'b0000001101: data <= 7'h00; 
        10'b0000001110: data <= 7'h00; 
        10'b0000001111: data <= 7'h00; 
        10'b0000010000: data <= 7'h00; 
        10'b0000010001: data <= 7'h00; 
        10'b0000010010: data <= 7'h00; 
        10'b0000010011: data <= 7'h00; 
        10'b0000010100: data <= 7'h00; 
        10'b0000010101: data <= 7'h00; 
        10'b0000010110: data <= 7'h00; 
        10'b0000010111: data <= 7'h00; 
        10'b0000011000: data <= 7'h00; 
        10'b0000011001: data <= 7'h00; 
        10'b0000011010: data <= 7'h00; 
        10'b0000011011: data <= 7'h00; 
        10'b0000011100: data <= 7'h00; 
        10'b0000011101: data <= 7'h00; 
        10'b0000011110: data <= 7'h00; 
        10'b0000011111: data <= 7'h00; 
        10'b0000100000: data <= 7'h00; 
        10'b0000100001: data <= 7'h00; 
        10'b0000100010: data <= 7'h00; 
        10'b0000100011: data <= 7'h00; 
        10'b0000100100: data <= 7'h00; 
        10'b0000100101: data <= 7'h00; 
        10'b0000100110: data <= 7'h00; 
        10'b0000100111: data <= 7'h00; 
        10'b0000101000: data <= 7'h00; 
        10'b0000101001: data <= 7'h00; 
        10'b0000101010: data <= 7'h00; 
        10'b0000101011: data <= 7'h00; 
        10'b0000101100: data <= 7'h00; 
        10'b0000101101: data <= 7'h00; 
        10'b0000101110: data <= 7'h00; 
        10'b0000101111: data <= 7'h00; 
        10'b0000110000: data <= 7'h00; 
        10'b0000110001: data <= 7'h00; 
        10'b0000110010: data <= 7'h00; 
        10'b0000110011: data <= 7'h00; 
        10'b0000110100: data <= 7'h00; 
        10'b0000110101: data <= 7'h00; 
        10'b0000110110: data <= 7'h00; 
        10'b0000110111: data <= 7'h00; 
        10'b0000111000: data <= 7'h00; 
        10'b0000111001: data <= 7'h00; 
        10'b0000111010: data <= 7'h00; 
        10'b0000111011: data <= 7'h00; 
        10'b0000111100: data <= 7'h00; 
        10'b0000111101: data <= 7'h00; 
        10'b0000111110: data <= 7'h00; 
        10'b0000111111: data <= 7'h00; 
        10'b0001000000: data <= 7'h00; 
        10'b0001000001: data <= 7'h00; 
        10'b0001000010: data <= 7'h00; 
        10'b0001000011: data <= 7'h00; 
        10'b0001000100: data <= 7'h00; 
        10'b0001000101: data <= 7'h00; 
        10'b0001000110: data <= 7'h00; 
        10'b0001000111: data <= 7'h00; 
        10'b0001001000: data <= 7'h00; 
        10'b0001001001: data <= 7'h00; 
        10'b0001001010: data <= 7'h00; 
        10'b0001001011: data <= 7'h00; 
        10'b0001001100: data <= 7'h00; 
        10'b0001001101: data <= 7'h00; 
        10'b0001001110: data <= 7'h00; 
        10'b0001001111: data <= 7'h00; 
        10'b0001010000: data <= 7'h00; 
        10'b0001010001: data <= 7'h00; 
        10'b0001010010: data <= 7'h00; 
        10'b0001010011: data <= 7'h00; 
        10'b0001010100: data <= 7'h00; 
        10'b0001010101: data <= 7'h00; 
        10'b0001010110: data <= 7'h00; 
        10'b0001010111: data <= 7'h00; 
        10'b0001011000: data <= 7'h00; 
        10'b0001011001: data <= 7'h00; 
        10'b0001011010: data <= 7'h00; 
        10'b0001011011: data <= 7'h00; 
        10'b0001011100: data <= 7'h00; 
        10'b0001011101: data <= 7'h00; 
        10'b0001011110: data <= 7'h00; 
        10'b0001011111: data <= 7'h00; 
        10'b0001100000: data <= 7'h00; 
        10'b0001100001: data <= 7'h00; 
        10'b0001100010: data <= 7'h00; 
        10'b0001100011: data <= 7'h00; 
        10'b0001100100: data <= 7'h00; 
        10'b0001100101: data <= 7'h00; 
        10'b0001100110: data <= 7'h00; 
        10'b0001100111: data <= 7'h00; 
        10'b0001101000: data <= 7'h00; 
        10'b0001101001: data <= 7'h00; 
        10'b0001101010: data <= 7'h00; 
        10'b0001101011: data <= 7'h00; 
        10'b0001101100: data <= 7'h00; 
        10'b0001101101: data <= 7'h00; 
        10'b0001101110: data <= 7'h00; 
        10'b0001101111: data <= 7'h00; 
        10'b0001110000: data <= 7'h00; 
        10'b0001110001: data <= 7'h00; 
        10'b0001110010: data <= 7'h00; 
        10'b0001110011: data <= 7'h00; 
        10'b0001110100: data <= 7'h00; 
        10'b0001110101: data <= 7'h00; 
        10'b0001110110: data <= 7'h00; 
        10'b0001110111: data <= 7'h00; 
        10'b0001111000: data <= 7'h00; 
        10'b0001111001: data <= 7'h00; 
        10'b0001111010: data <= 7'h00; 
        10'b0001111011: data <= 7'h00; 
        10'b0001111100: data <= 7'h00; 
        10'b0001111101: data <= 7'h00; 
        10'b0001111110: data <= 7'h00; 
        10'b0001111111: data <= 7'h7f; 
        10'b0010000000: data <= 7'h00; 
        10'b0010000001: data <= 7'h00; 
        10'b0010000010: data <= 7'h00; 
        10'b0010000011: data <= 7'h00; 
        10'b0010000100: data <= 7'h00; 
        10'b0010000101: data <= 7'h00; 
        10'b0010000110: data <= 7'h00; 
        10'b0010000111: data <= 7'h00; 
        10'b0010001000: data <= 7'h00; 
        10'b0010001001: data <= 7'h00; 
        10'b0010001010: data <= 7'h00; 
        10'b0010001011: data <= 7'h00; 
        10'b0010001100: data <= 7'h00; 
        10'b0010001101: data <= 7'h00; 
        10'b0010001110: data <= 7'h00; 
        10'b0010001111: data <= 7'h00; 
        10'b0010010000: data <= 7'h00; 
        10'b0010010001: data <= 7'h00; 
        10'b0010010010: data <= 7'h00; 
        10'b0010010011: data <= 7'h00; 
        10'b0010010100: data <= 7'h00; 
        10'b0010010101: data <= 7'h00; 
        10'b0010010110: data <= 7'h00; 
        10'b0010010111: data <= 7'h00; 
        10'b0010011000: data <= 7'h00; 
        10'b0010011001: data <= 7'h00; 
        10'b0010011010: data <= 7'h7f; 
        10'b0010011011: data <= 7'h7f; 
        10'b0010011100: data <= 7'h7f; 
        10'b0010011101: data <= 7'h7f; 
        10'b0010011110: data <= 7'h00; 
        10'b0010011111: data <= 7'h00; 
        10'b0010100000: data <= 7'h00; 
        10'b0010100001: data <= 7'h00; 
        10'b0010100010: data <= 7'h00; 
        10'b0010100011: data <= 7'h00; 
        10'b0010100100: data <= 7'h00; 
        10'b0010100101: data <= 7'h00; 
        10'b0010100110: data <= 7'h00; 
        10'b0010100111: data <= 7'h00; 
        10'b0010101000: data <= 7'h00; 
        10'b0010101001: data <= 7'h00; 
        10'b0010101010: data <= 7'h00; 
        10'b0010101011: data <= 7'h00; 
        10'b0010101100: data <= 7'h00; 
        10'b0010101101: data <= 7'h00; 
        10'b0010101110: data <= 7'h00; 
        10'b0010101111: data <= 7'h00; 
        10'b0010110000: data <= 7'h00; 
        10'b0010110001: data <= 7'h00; 
        10'b0010110010: data <= 7'h00; 
        10'b0010110011: data <= 7'h00; 
        10'b0010110100: data <= 7'h00; 
        10'b0010110101: data <= 7'h00; 
        10'b0010110110: data <= 7'h01; 
        10'b0010110111: data <= 7'h00; 
        10'b0010111000: data <= 7'h00; 
        10'b0010111001: data <= 7'h00; 
        10'b0010111010: data <= 7'h00; 
        10'b0010111011: data <= 7'h00; 
        10'b0010111100: data <= 7'h00; 
        10'b0010111101: data <= 7'h00; 
        10'b0010111110: data <= 7'h00; 
        10'b0010111111: data <= 7'h00; 
        10'b0011000000: data <= 7'h00; 
        10'b0011000001: data <= 7'h00; 
        10'b0011000010: data <= 7'h00; 
        10'b0011000011: data <= 7'h00; 
        10'b0011000100: data <= 7'h00; 
        10'b0011000101: data <= 7'h00; 
        10'b0011000110: data <= 7'h00; 
        10'b0011000111: data <= 7'h00; 
        10'b0011001000: data <= 7'h00; 
        10'b0011001001: data <= 7'h00; 
        10'b0011001010: data <= 7'h00; 
        10'b0011001011: data <= 7'h00; 
        10'b0011001100: data <= 7'h00; 
        10'b0011001101: data <= 7'h00; 
        10'b0011001110: data <= 7'h00; 
        10'b0011001111: data <= 7'h00; 
        10'b0011010000: data <= 7'h00; 
        10'b0011010001: data <= 7'h01; 
        10'b0011010010: data <= 7'h01; 
        10'b0011010011: data <= 7'h01; 
        10'b0011010100: data <= 7'h01; 
        10'b0011010101: data <= 7'h00; 
        10'b0011010110: data <= 7'h00; 
        10'b0011010111: data <= 7'h00; 
        10'b0011011000: data <= 7'h00; 
        10'b0011011001: data <= 7'h00; 
        10'b0011011010: data <= 7'h00; 
        10'b0011011011: data <= 7'h00; 
        10'b0011011100: data <= 7'h00; 
        10'b0011011101: data <= 7'h00; 
        10'b0011011110: data <= 7'h00; 
        10'b0011011111: data <= 7'h00; 
        10'b0011100000: data <= 7'h00; 
        10'b0011100001: data <= 7'h00; 
        10'b0011100010: data <= 7'h00; 
        10'b0011100011: data <= 7'h00; 
        10'b0011100100: data <= 7'h00; 
        10'b0011100101: data <= 7'h00; 
        10'b0011100110: data <= 7'h00; 
        10'b0011100111: data <= 7'h7f; 
        10'b0011101000: data <= 7'h00; 
        10'b0011101001: data <= 7'h00; 
        10'b0011101010: data <= 7'h00; 
        10'b0011101011: data <= 7'h00; 
        10'b0011101100: data <= 7'h00; 
        10'b0011101101: data <= 7'h00; 
        10'b0011101110: data <= 7'h01; 
        10'b0011101111: data <= 7'h00; 
        10'b0011110000: data <= 7'h00; 
        10'b0011110001: data <= 7'h00; 
        10'b0011110010: data <= 7'h00; 
        10'b0011110011: data <= 7'h00; 
        10'b0011110100: data <= 7'h00; 
        10'b0011110101: data <= 7'h00; 
        10'b0011110110: data <= 7'h00; 
        10'b0011110111: data <= 7'h00; 
        10'b0011111000: data <= 7'h00; 
        10'b0011111001: data <= 7'h00; 
        10'b0011111010: data <= 7'h00; 
        10'b0011111011: data <= 7'h00; 
        10'b0011111100: data <= 7'h00; 
        10'b0011111101: data <= 7'h00; 
        10'b0011111110: data <= 7'h00; 
        10'b0011111111: data <= 7'h00; 
        10'b0100000000: data <= 7'h00; 
        10'b0100000001: data <= 7'h00; 
        10'b0100000010: data <= 7'h00; 
        10'b0100000011: data <= 7'h00; 
        10'b0100000100: data <= 7'h00; 
        10'b0100000101: data <= 7'h00; 
        10'b0100000110: data <= 7'h00; 
        10'b0100000111: data <= 7'h00; 
        10'b0100001000: data <= 7'h00; 
        10'b0100001001: data <= 7'h00; 
        10'b0100001010: data <= 7'h00; 
        10'b0100001011: data <= 7'h00; 
        10'b0100001100: data <= 7'h00; 
        10'b0100001101: data <= 7'h00; 
        10'b0100001110: data <= 7'h00; 
        10'b0100001111: data <= 7'h00; 
        10'b0100010000: data <= 7'h00; 
        10'b0100010001: data <= 7'h00; 
        10'b0100010010: data <= 7'h00; 
        10'b0100010011: data <= 7'h00; 
        10'b0100010100: data <= 7'h00; 
        10'b0100010101: data <= 7'h00; 
        10'b0100010110: data <= 7'h00; 
        10'b0100010111: data <= 7'h00; 
        10'b0100011000: data <= 7'h00; 
        10'b0100011001: data <= 7'h00; 
        10'b0100011010: data <= 7'h00; 
        10'b0100011011: data <= 7'h00; 
        10'b0100011100: data <= 7'h00; 
        10'b0100011101: data <= 7'h00; 
        10'b0100011110: data <= 7'h00; 
        10'b0100011111: data <= 7'h00; 
        10'b0100100000: data <= 7'h00; 
        10'b0100100001: data <= 7'h00; 
        10'b0100100010: data <= 7'h00; 
        10'b0100100011: data <= 7'h00; 
        10'b0100100100: data <= 7'h00; 
        10'b0100100101: data <= 7'h00; 
        10'b0100100110: data <= 7'h00; 
        10'b0100100111: data <= 7'h00; 
        10'b0100101000: data <= 7'h00; 
        10'b0100101001: data <= 7'h00; 
        10'b0100101010: data <= 7'h00; 
        10'b0100101011: data <= 7'h00; 
        10'b0100101100: data <= 7'h00; 
        10'b0100101101: data <= 7'h00; 
        10'b0100101110: data <= 7'h00; 
        10'b0100101111: data <= 7'h00; 
        10'b0100110000: data <= 7'h00; 
        10'b0100110001: data <= 7'h00; 
        10'b0100110010: data <= 7'h00; 
        10'b0100110011: data <= 7'h00; 
        10'b0100110100: data <= 7'h00; 
        10'b0100110101: data <= 7'h00; 
        10'b0100110110: data <= 7'h00; 
        10'b0100110111: data <= 7'h00; 
        10'b0100111000: data <= 7'h00; 
        10'b0100111001: data <= 7'h00; 
        10'b0100111010: data <= 7'h01; 
        10'b0100111011: data <= 7'h00; 
        10'b0100111100: data <= 7'h01; 
        10'b0100111101: data <= 7'h00; 
        10'b0100111110: data <= 7'h00; 
        10'b0100111111: data <= 7'h00; 
        10'b0101000000: data <= 7'h00; 
        10'b0101000001: data <= 7'h00; 
        10'b0101000010: data <= 7'h00; 
        10'b0101000011: data <= 7'h00; 
        10'b0101000100: data <= 7'h00; 
        10'b0101000101: data <= 7'h01; 
        10'b0101000110: data <= 7'h00; 
        10'b0101000111: data <= 7'h00; 
        10'b0101001000: data <= 7'h01; 
        10'b0101001001: data <= 7'h00; 
        10'b0101001010: data <= 7'h00; 
        10'b0101001011: data <= 7'h00; 
        10'b0101001100: data <= 7'h00; 
        10'b0101001101: data <= 7'h00; 
        10'b0101001110: data <= 7'h00; 
        10'b0101001111: data <= 7'h00; 
        10'b0101010000: data <= 7'h00; 
        10'b0101010001: data <= 7'h00; 
        10'b0101010010: data <= 7'h00; 
        10'b0101010011: data <= 7'h00; 
        10'b0101010100: data <= 7'h00; 
        10'b0101010101: data <= 7'h01; 
        10'b0101010110: data <= 7'h01; 
        10'b0101010111: data <= 7'h00; 
        10'b0101011000: data <= 7'h00; 
        10'b0101011001: data <= 7'h01; 
        10'b0101011010: data <= 7'h00; 
        10'b0101011011: data <= 7'h00; 
        10'b0101011100: data <= 7'h00; 
        10'b0101011101: data <= 7'h00; 
        10'b0101011110: data <= 7'h01; 
        10'b0101011111: data <= 7'h01; 
        10'b0101100000: data <= 7'h00; 
        10'b0101100001: data <= 7'h01; 
        10'b0101100010: data <= 7'h01; 
        10'b0101100011: data <= 7'h01; 
        10'b0101100100: data <= 7'h01; 
        10'b0101100101: data <= 7'h01; 
        10'b0101100110: data <= 7'h00; 
        10'b0101100111: data <= 7'h00; 
        10'b0101101000: data <= 7'h00; 
        10'b0101101001: data <= 7'h00; 
        10'b0101101010: data <= 7'h00; 
        10'b0101101011: data <= 7'h00; 
        10'b0101101100: data <= 7'h00; 
        10'b0101101101: data <= 7'h00; 
        10'b0101101110: data <= 7'h00; 
        10'b0101101111: data <= 7'h00; 
        10'b0101110000: data <= 7'h00; 
        10'b0101110001: data <= 7'h00; 
        10'b0101110010: data <= 7'h00; 
        10'b0101110011: data <= 7'h00; 
        10'b0101110100: data <= 7'h00; 
        10'b0101110101: data <= 7'h00; 
        10'b0101110110: data <= 7'h00; 
        10'b0101110111: data <= 7'h00; 
        10'b0101111000: data <= 7'h00; 
        10'b0101111001: data <= 7'h00; 
        10'b0101111010: data <= 7'h01; 
        10'b0101111011: data <= 7'h00; 
        10'b0101111100: data <= 7'h01; 
        10'b0101111101: data <= 7'h01; 
        10'b0101111110: data <= 7'h01; 
        10'b0101111111: data <= 7'h01; 
        10'b0110000000: data <= 7'h01; 
        10'b0110000001: data <= 7'h00; 
        10'b0110000010: data <= 7'h00; 
        10'b0110000011: data <= 7'h00; 
        10'b0110000100: data <= 7'h00; 
        10'b0110000101: data <= 7'h00; 
        10'b0110000110: data <= 7'h00; 
        10'b0110000111: data <= 7'h00; 
        10'b0110001000: data <= 7'h00; 
        10'b0110001001: data <= 7'h00; 
        10'b0110001010: data <= 7'h00; 
        10'b0110001011: data <= 7'h00; 
        10'b0110001100: data <= 7'h00; 
        10'b0110001101: data <= 7'h00; 
        10'b0110001110: data <= 7'h00; 
        10'b0110001111: data <= 7'h00; 
        10'b0110010000: data <= 7'h00; 
        10'b0110010001: data <= 7'h00; 
        10'b0110010010: data <= 7'h00; 
        10'b0110010011: data <= 7'h00; 
        10'b0110010100: data <= 7'h00; 
        10'b0110010101: data <= 7'h00; 
        10'b0110010110: data <= 7'h00; 
        10'b0110010111: data <= 7'h00; 
        10'b0110011000: data <= 7'h00; 
        10'b0110011001: data <= 7'h00; 
        10'b0110011010: data <= 7'h00; 
        10'b0110011011: data <= 7'h00; 
        10'b0110011100: data <= 7'h00; 
        10'b0110011101: data <= 7'h00; 
        10'b0110011110: data <= 7'h00; 
        10'b0110011111: data <= 7'h00; 
        10'b0110100000: data <= 7'h00; 
        10'b0110100001: data <= 7'h00; 
        10'b0110100010: data <= 7'h00; 
        10'b0110100011: data <= 7'h00; 
        10'b0110100100: data <= 7'h00; 
        10'b0110100101: data <= 7'h00; 
        10'b0110100110: data <= 7'h00; 
        10'b0110100111: data <= 7'h00; 
        10'b0110101000: data <= 7'h00; 
        10'b0110101001: data <= 7'h00; 
        10'b0110101010: data <= 7'h00; 
        10'b0110101011: data <= 7'h00; 
        10'b0110101100: data <= 7'h00; 
        10'b0110101101: data <= 7'h00; 
        10'b0110101110: data <= 7'h00; 
        10'b0110101111: data <= 7'h00; 
        10'b0110110000: data <= 7'h00; 
        10'b0110110001: data <= 7'h00; 
        10'b0110110010: data <= 7'h00; 
        10'b0110110011: data <= 7'h00; 
        10'b0110110100: data <= 7'h01; 
        10'b0110110101: data <= 7'h01; 
        10'b0110110110: data <= 7'h00; 
        10'b0110110111: data <= 7'h00; 
        10'b0110111000: data <= 7'h00; 
        10'b0110111001: data <= 7'h00; 
        10'b0110111010: data <= 7'h00; 
        10'b0110111011: data <= 7'h00; 
        10'b0110111100: data <= 7'h00; 
        10'b0110111101: data <= 7'h00; 
        10'b0110111110: data <= 7'h00; 
        10'b0110111111: data <= 7'h00; 
        10'b0111000000: data <= 7'h00; 
        10'b0111000001: data <= 7'h00; 
        10'b0111000010: data <= 7'h00; 
        10'b0111000011: data <= 7'h00; 
        10'b0111000100: data <= 7'h00; 
        10'b0111000101: data <= 7'h00; 
        10'b0111000110: data <= 7'h00; 
        10'b0111000111: data <= 7'h00; 
        10'b0111001000: data <= 7'h00; 
        10'b0111001001: data <= 7'h00; 
        10'b0111001010: data <= 7'h00; 
        10'b0111001011: data <= 7'h00; 
        10'b0111001100: data <= 7'h00; 
        10'b0111001101: data <= 7'h00; 
        10'b0111001110: data <= 7'h00; 
        10'b0111001111: data <= 7'h00; 
        10'b0111010000: data <= 7'h00; 
        10'b0111010001: data <= 7'h00; 
        10'b0111010010: data <= 7'h00; 
        10'b0111010011: data <= 7'h00; 
        10'b0111010100: data <= 7'h00; 
        10'b0111010101: data <= 7'h7f; 
        10'b0111010110: data <= 7'h00; 
        10'b0111010111: data <= 7'h00; 
        10'b0111011000: data <= 7'h00; 
        10'b0111011001: data <= 7'h00; 
        10'b0111011010: data <= 7'h00; 
        10'b0111011011: data <= 7'h00; 
        10'b0111011100: data <= 7'h00; 
        10'b0111011101: data <= 7'h00; 
        10'b0111011110: data <= 7'h00; 
        10'b0111011111: data <= 7'h00; 
        10'b0111100000: data <= 7'h00; 
        10'b0111100001: data <= 7'h00; 
        10'b0111100010: data <= 7'h00; 
        10'b0111100011: data <= 7'h00; 
        10'b0111100100: data <= 7'h00; 
        10'b0111100101: data <= 7'h00; 
        10'b0111100110: data <= 7'h00; 
        10'b0111100111: data <= 7'h00; 
        10'b0111101000: data <= 7'h00; 
        10'b0111101001: data <= 7'h00; 
        10'b0111101010: data <= 7'h00; 
        10'b0111101011: data <= 7'h00; 
        10'b0111101100: data <= 7'h00; 
        10'b0111101101: data <= 7'h00; 
        10'b0111101110: data <= 7'h00; 
        10'b0111101111: data <= 7'h00; 
        10'b0111110000: data <= 7'h00; 
        10'b0111110001: data <= 7'h00; 
        10'b0111110010: data <= 7'h00; 
        10'b0111110011: data <= 7'h00; 
        10'b0111110100: data <= 7'h00; 
        10'b0111110101: data <= 7'h00; 
        10'b0111110110: data <= 7'h00; 
        10'b0111110111: data <= 7'h00; 
        10'b0111111000: data <= 7'h00; 
        10'b0111111001: data <= 7'h00; 
        10'b0111111010: data <= 7'h00; 
        10'b0111111011: data <= 7'h00; 
        10'b0111111100: data <= 7'h00; 
        10'b0111111101: data <= 7'h00; 
        10'b0111111110: data <= 7'h00; 
        10'b0111111111: data <= 7'h00; 
        10'b1000000000: data <= 7'h00; 
        10'b1000000001: data <= 7'h00; 
        10'b1000000010: data <= 7'h00; 
        10'b1000000011: data <= 7'h00; 
        10'b1000000100: data <= 7'h00; 
        10'b1000000101: data <= 7'h00; 
        10'b1000000110: data <= 7'h00; 
        10'b1000000111: data <= 7'h00; 
        10'b1000001000: data <= 7'h00; 
        10'b1000001001: data <= 7'h00; 
        10'b1000001010: data <= 7'h00; 
        10'b1000001011: data <= 7'h00; 
        10'b1000001100: data <= 7'h00; 
        10'b1000001101: data <= 7'h00; 
        10'b1000001110: data <= 7'h00; 
        10'b1000001111: data <= 7'h00; 
        10'b1000010000: data <= 7'h00; 
        10'b1000010001: data <= 7'h00; 
        10'b1000010010: data <= 7'h00; 
        10'b1000010011: data <= 7'h00; 
        10'b1000010100: data <= 7'h00; 
        10'b1000010101: data <= 7'h00; 
        10'b1000010110: data <= 7'h00; 
        10'b1000010111: data <= 7'h00; 
        10'b1000011000: data <= 7'h00; 
        10'b1000011001: data <= 7'h00; 
        10'b1000011010: data <= 7'h00; 
        10'b1000011011: data <= 7'h00; 
        10'b1000011100: data <= 7'h00; 
        10'b1000011101: data <= 7'h00; 
        10'b1000011110: data <= 7'h00; 
        10'b1000011111: data <= 7'h00; 
        10'b1000100000: data <= 7'h7f; 
        10'b1000100001: data <= 7'h00; 
        10'b1000100010: data <= 7'h00; 
        10'b1000100011: data <= 7'h00; 
        10'b1000100100: data <= 7'h00; 
        10'b1000100101: data <= 7'h00; 
        10'b1000100110: data <= 7'h00; 
        10'b1000100111: data <= 7'h00; 
        10'b1000101000: data <= 7'h00; 
        10'b1000101001: data <= 7'h00; 
        10'b1000101010: data <= 7'h00; 
        10'b1000101011: data <= 7'h00; 
        10'b1000101100: data <= 7'h00; 
        10'b1000101101: data <= 7'h00; 
        10'b1000101110: data <= 7'h00; 
        10'b1000101111: data <= 7'h00; 
        10'b1000110000: data <= 7'h00; 
        10'b1000110001: data <= 7'h00; 
        10'b1000110010: data <= 7'h00; 
        10'b1000110011: data <= 7'h00; 
        10'b1000110100: data <= 7'h00; 
        10'b1000110101: data <= 7'h00; 
        10'b1000110110: data <= 7'h00; 
        10'b1000110111: data <= 7'h7f; 
        10'b1000111000: data <= 7'h7f; 
        10'b1000111001: data <= 7'h7f; 
        10'b1000111010: data <= 7'h7f; 
        10'b1000111011: data <= 7'h7f; 
        10'b1000111100: data <= 7'h7f; 
        10'b1000111101: data <= 7'h00; 
        10'b1000111110: data <= 7'h00; 
        10'b1000111111: data <= 7'h00; 
        10'b1001000000: data <= 7'h00; 
        10'b1001000001: data <= 7'h00; 
        10'b1001000010: data <= 7'h00; 
        10'b1001000011: data <= 7'h00; 
        10'b1001000100: data <= 7'h00; 
        10'b1001000101: data <= 7'h00; 
        10'b1001000110: data <= 7'h00; 
        10'b1001000111: data <= 7'h00; 
        10'b1001001000: data <= 7'h00; 
        10'b1001001001: data <= 7'h00; 
        10'b1001001010: data <= 7'h00; 
        10'b1001001011: data <= 7'h00; 
        10'b1001001100: data <= 7'h00; 
        10'b1001001101: data <= 7'h00; 
        10'b1001001110: data <= 7'h00; 
        10'b1001001111: data <= 7'h00; 
        10'b1001010000: data <= 7'h00; 
        10'b1001010001: data <= 7'h00; 
        10'b1001010010: data <= 7'h00; 
        10'b1001010011: data <= 7'h7f; 
        10'b1001010100: data <= 7'h7f; 
        10'b1001010101: data <= 7'h7f; 
        10'b1001010110: data <= 7'h7f; 
        10'b1001010111: data <= 7'h7f; 
        10'b1001011000: data <= 7'h00; 
        10'b1001011001: data <= 7'h00; 
        10'b1001011010: data <= 7'h00; 
        10'b1001011011: data <= 7'h00; 
        10'b1001011100: data <= 7'h00; 
        10'b1001011101: data <= 7'h00; 
        10'b1001011110: data <= 7'h00; 
        10'b1001011111: data <= 7'h00; 
        10'b1001100000: data <= 7'h00; 
        10'b1001100001: data <= 7'h00; 
        10'b1001100010: data <= 7'h00; 
        10'b1001100011: data <= 7'h00; 
        10'b1001100100: data <= 7'h00; 
        10'b1001100101: data <= 7'h00; 
        10'b1001100110: data <= 7'h00; 
        10'b1001100111: data <= 7'h00; 
        10'b1001101000: data <= 7'h00; 
        10'b1001101001: data <= 7'h00; 
        10'b1001101010: data <= 7'h00; 
        10'b1001101011: data <= 7'h00; 
        10'b1001101100: data <= 7'h00; 
        10'b1001101101: data <= 7'h00; 
        10'b1001101110: data <= 7'h00; 
        10'b1001101111: data <= 7'h00; 
        10'b1001110000: data <= 7'h00; 
        10'b1001110001: data <= 7'h00; 
        10'b1001110010: data <= 7'h00; 
        10'b1001110011: data <= 7'h00; 
        10'b1001110100: data <= 7'h00; 
        10'b1001110101: data <= 7'h00; 
        10'b1001110110: data <= 7'h00; 
        10'b1001110111: data <= 7'h00; 
        10'b1001111000: data <= 7'h00; 
        10'b1001111001: data <= 7'h00; 
        10'b1001111010: data <= 7'h00; 
        10'b1001111011: data <= 7'h00; 
        10'b1001111100: data <= 7'h00; 
        10'b1001111101: data <= 7'h00; 
        10'b1001111110: data <= 7'h00; 
        10'b1001111111: data <= 7'h00; 
        10'b1010000000: data <= 7'h00; 
        10'b1010000001: data <= 7'h00; 
        10'b1010000010: data <= 7'h00; 
        10'b1010000011: data <= 7'h00; 
        10'b1010000100: data <= 7'h00; 
        10'b1010000101: data <= 7'h00; 
        10'b1010000110: data <= 7'h00; 
        10'b1010000111: data <= 7'h00; 
        10'b1010001000: data <= 7'h00; 
        10'b1010001001: data <= 7'h00; 
        10'b1010001010: data <= 7'h00; 
        10'b1010001011: data <= 7'h00; 
        10'b1010001100: data <= 7'h00; 
        10'b1010001101: data <= 7'h00; 
        10'b1010001110: data <= 7'h00; 
        10'b1010001111: data <= 7'h00; 
        10'b1010010000: data <= 7'h00; 
        10'b1010010001: data <= 7'h00; 
        10'b1010010010: data <= 7'h00; 
        10'b1010010011: data <= 7'h00; 
        10'b1010010100: data <= 7'h00; 
        10'b1010010101: data <= 7'h00; 
        10'b1010010110: data <= 7'h00; 
        10'b1010010111: data <= 7'h00; 
        10'b1010011000: data <= 7'h00; 
        10'b1010011001: data <= 7'h00; 
        10'b1010011010: data <= 7'h00; 
        10'b1010011011: data <= 7'h00; 
        10'b1010011100: data <= 7'h00; 
        10'b1010011101: data <= 7'h00; 
        10'b1010011110: data <= 7'h00; 
        10'b1010011111: data <= 7'h00; 
        10'b1010100000: data <= 7'h00; 
        10'b1010100001: data <= 7'h00; 
        10'b1010100010: data <= 7'h00; 
        10'b1010100011: data <= 7'h00; 
        10'b1010100100: data <= 7'h00; 
        10'b1010100101: data <= 7'h00; 
        10'b1010100110: data <= 7'h00; 
        10'b1010100111: data <= 7'h00; 
        10'b1010101000: data <= 7'h00; 
        10'b1010101001: data <= 7'h00; 
        10'b1010101010: data <= 7'h00; 
        10'b1010101011: data <= 7'h00; 
        10'b1010101100: data <= 7'h00; 
        10'b1010101101: data <= 7'h00; 
        10'b1010101110: data <= 7'h00; 
        10'b1010101111: data <= 7'h00; 
        10'b1010110000: data <= 7'h00; 
        10'b1010110001: data <= 7'h00; 
        10'b1010110010: data <= 7'h00; 
        10'b1010110011: data <= 7'h00; 
        10'b1010110100: data <= 7'h00; 
        10'b1010110101: data <= 7'h00; 
        10'b1010110110: data <= 7'h00; 
        10'b1010110111: data <= 7'h00; 
        10'b1010111000: data <= 7'h00; 
        10'b1010111001: data <= 7'h00; 
        10'b1010111010: data <= 7'h00; 
        10'b1010111011: data <= 7'h00; 
        10'b1010111100: data <= 7'h00; 
        10'b1010111101: data <= 7'h00; 
        10'b1010111110: data <= 7'h00; 
        10'b1010111111: data <= 7'h00; 
        10'b1011000000: data <= 7'h00; 
        10'b1011000001: data <= 7'h00; 
        10'b1011000010: data <= 7'h00; 
        10'b1011000011: data <= 7'h00; 
        10'b1011000100: data <= 7'h00; 
        10'b1011000101: data <= 7'h00; 
        10'b1011000110: data <= 7'h00; 
        10'b1011000111: data <= 7'h00; 
        10'b1011001000: data <= 7'h00; 
        10'b1011001001: data <= 7'h00; 
        10'b1011001010: data <= 7'h00; 
        10'b1011001011: data <= 7'h00; 
        10'b1011001100: data <= 7'h00; 
        10'b1011001101: data <= 7'h01; 
        10'b1011001110: data <= 7'h01; 
        10'b1011001111: data <= 7'h01; 
        10'b1011010000: data <= 7'h01; 
        10'b1011010001: data <= 7'h00; 
        10'b1011010010: data <= 7'h00; 
        10'b1011010011: data <= 7'h00; 
        10'b1011010100: data <= 7'h00; 
        10'b1011010101: data <= 7'h00; 
        10'b1011010110: data <= 7'h00; 
        10'b1011010111: data <= 7'h00; 
        10'b1011011000: data <= 7'h00; 
        10'b1011011001: data <= 7'h00; 
        10'b1011011010: data <= 7'h00; 
        10'b1011011011: data <= 7'h00; 
        10'b1011011100: data <= 7'h00; 
        10'b1011011101: data <= 7'h00; 
        10'b1011011110: data <= 7'h00; 
        10'b1011011111: data <= 7'h00; 
        10'b1011100000: data <= 7'h00; 
        10'b1011100001: data <= 7'h00; 
        10'b1011100010: data <= 7'h00; 
        10'b1011100011: data <= 7'h00; 
        10'b1011100100: data <= 7'h01; 
        10'b1011100101: data <= 7'h01; 
        10'b1011100110: data <= 7'h01; 
        10'b1011100111: data <= 7'h00; 
        10'b1011101000: data <= 7'h00; 
        10'b1011101001: data <= 7'h00; 
        10'b1011101010: data <= 7'h00; 
        10'b1011101011: data <= 7'h00; 
        10'b1011101100: data <= 7'h00; 
        10'b1011101101: data <= 7'h00; 
        10'b1011101110: data <= 7'h00; 
        10'b1011101111: data <= 7'h00; 
        10'b1011110000: data <= 7'h00; 
        10'b1011110001: data <= 7'h00; 
        10'b1011110010: data <= 7'h00; 
        10'b1011110011: data <= 7'h00; 
        10'b1011110100: data <= 7'h00; 
        10'b1011110101: data <= 7'h00; 
        10'b1011110110: data <= 7'h00; 
        10'b1011110111: data <= 7'h00; 
        10'b1011111000: data <= 7'h00; 
        10'b1011111001: data <= 7'h00; 
        10'b1011111010: data <= 7'h00; 
        10'b1011111011: data <= 7'h00; 
        10'b1011111100: data <= 7'h00; 
        10'b1011111101: data <= 7'h00; 
        10'b1011111110: data <= 7'h00; 
        10'b1011111111: data <= 7'h00; 
        10'b1100000000: data <= 7'h00; 
        10'b1100000001: data <= 7'h00; 
        10'b1100000010: data <= 7'h00; 
        10'b1100000011: data <= 7'h00; 
        10'b1100000100: data <= 7'h00; 
        10'b1100000101: data <= 7'h00; 
        10'b1100000110: data <= 7'h00; 
        10'b1100000111: data <= 7'h00; 
        10'b1100001000: data <= 7'h00; 
        10'b1100001001: data <= 7'h00; 
        10'b1100001010: data <= 7'h00; 
        10'b1100001011: data <= 7'h00; 
        10'b1100001100: data <= 7'h00; 
        10'b1100001101: data <= 7'h00; 
        10'b1100001110: data <= 7'h00; 
        10'b1100001111: data <= 7'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 2) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 8'h00; 
        10'b0000000001: data <= 8'h00; 
        10'b0000000010: data <= 8'h00; 
        10'b0000000011: data <= 8'h00; 
        10'b0000000100: data <= 8'h00; 
        10'b0000000101: data <= 8'h00; 
        10'b0000000110: data <= 8'h00; 
        10'b0000000111: data <= 8'h00; 
        10'b0000001000: data <= 8'h00; 
        10'b0000001001: data <= 8'h00; 
        10'b0000001010: data <= 8'h00; 
        10'b0000001011: data <= 8'h00; 
        10'b0000001100: data <= 8'h00; 
        10'b0000001101: data <= 8'h00; 
        10'b0000001110: data <= 8'h00; 
        10'b0000001111: data <= 8'h00; 
        10'b0000010000: data <= 8'h00; 
        10'b0000010001: data <= 8'h00; 
        10'b0000010010: data <= 8'h00; 
        10'b0000010011: data <= 8'h00; 
        10'b0000010100: data <= 8'h00; 
        10'b0000010101: data <= 8'h00; 
        10'b0000010110: data <= 8'h00; 
        10'b0000010111: data <= 8'h00; 
        10'b0000011000: data <= 8'h00; 
        10'b0000011001: data <= 8'h00; 
        10'b0000011010: data <= 8'h00; 
        10'b0000011011: data <= 8'h00; 
        10'b0000011100: data <= 8'h00; 
        10'b0000011101: data <= 8'h00; 
        10'b0000011110: data <= 8'h00; 
        10'b0000011111: data <= 8'h00; 
        10'b0000100000: data <= 8'h00; 
        10'b0000100001: data <= 8'h00; 
        10'b0000100010: data <= 8'h00; 
        10'b0000100011: data <= 8'h00; 
        10'b0000100100: data <= 8'h00; 
        10'b0000100101: data <= 8'h00; 
        10'b0000100110: data <= 8'h00; 
        10'b0000100111: data <= 8'h00; 
        10'b0000101000: data <= 8'h00; 
        10'b0000101001: data <= 8'h00; 
        10'b0000101010: data <= 8'h00; 
        10'b0000101011: data <= 8'h00; 
        10'b0000101100: data <= 8'h00; 
        10'b0000101101: data <= 8'h00; 
        10'b0000101110: data <= 8'h00; 
        10'b0000101111: data <= 8'h00; 
        10'b0000110000: data <= 8'h00; 
        10'b0000110001: data <= 8'h00; 
        10'b0000110010: data <= 8'h00; 
        10'b0000110011: data <= 8'h00; 
        10'b0000110100: data <= 8'h00; 
        10'b0000110101: data <= 8'h00; 
        10'b0000110110: data <= 8'h00; 
        10'b0000110111: data <= 8'h00; 
        10'b0000111000: data <= 8'h00; 
        10'b0000111001: data <= 8'h00; 
        10'b0000111010: data <= 8'h00; 
        10'b0000111011: data <= 8'h00; 
        10'b0000111100: data <= 8'h00; 
        10'b0000111101: data <= 8'h00; 
        10'b0000111110: data <= 8'h00; 
        10'b0000111111: data <= 8'h00; 
        10'b0001000000: data <= 8'h00; 
        10'b0001000001: data <= 8'h00; 
        10'b0001000010: data <= 8'h00; 
        10'b0001000011: data <= 8'h00; 
        10'b0001000100: data <= 8'h00; 
        10'b0001000101: data <= 8'h00; 
        10'b0001000110: data <= 8'h00; 
        10'b0001000111: data <= 8'h00; 
        10'b0001001000: data <= 8'h00; 
        10'b0001001001: data <= 8'h00; 
        10'b0001001010: data <= 8'h00; 
        10'b0001001011: data <= 8'h00; 
        10'b0001001100: data <= 8'h00; 
        10'b0001001101: data <= 8'h00; 
        10'b0001001110: data <= 8'h00; 
        10'b0001001111: data <= 8'h00; 
        10'b0001010000: data <= 8'h00; 
        10'b0001010001: data <= 8'h00; 
        10'b0001010010: data <= 8'h00; 
        10'b0001010011: data <= 8'h00; 
        10'b0001010100: data <= 8'h00; 
        10'b0001010101: data <= 8'h00; 
        10'b0001010110: data <= 8'h00; 
        10'b0001010111: data <= 8'h00; 
        10'b0001011000: data <= 8'h00; 
        10'b0001011001: data <= 8'h00; 
        10'b0001011010: data <= 8'h00; 
        10'b0001011011: data <= 8'h00; 
        10'b0001011100: data <= 8'h00; 
        10'b0001011101: data <= 8'h00; 
        10'b0001011110: data <= 8'h00; 
        10'b0001011111: data <= 8'h00; 
        10'b0001100000: data <= 8'h00; 
        10'b0001100001: data <= 8'h00; 
        10'b0001100010: data <= 8'h00; 
        10'b0001100011: data <= 8'h00; 
        10'b0001100100: data <= 8'h00; 
        10'b0001100101: data <= 8'h00; 
        10'b0001100110: data <= 8'h00; 
        10'b0001100111: data <= 8'h00; 
        10'b0001101000: data <= 8'h00; 
        10'b0001101001: data <= 8'h00; 
        10'b0001101010: data <= 8'h00; 
        10'b0001101011: data <= 8'h00; 
        10'b0001101100: data <= 8'h00; 
        10'b0001101101: data <= 8'h00; 
        10'b0001101110: data <= 8'h00; 
        10'b0001101111: data <= 8'h00; 
        10'b0001110000: data <= 8'h00; 
        10'b0001110001: data <= 8'h00; 
        10'b0001110010: data <= 8'h00; 
        10'b0001110011: data <= 8'h00; 
        10'b0001110100: data <= 8'h00; 
        10'b0001110101: data <= 8'h00; 
        10'b0001110110: data <= 8'h00; 
        10'b0001110111: data <= 8'h00; 
        10'b0001111000: data <= 8'h00; 
        10'b0001111001: data <= 8'h00; 
        10'b0001111010: data <= 8'h00; 
        10'b0001111011: data <= 8'h00; 
        10'b0001111100: data <= 8'h00; 
        10'b0001111101: data <= 8'hff; 
        10'b0001111110: data <= 8'hff; 
        10'b0001111111: data <= 8'hff; 
        10'b0010000000: data <= 8'hff; 
        10'b0010000001: data <= 8'hff; 
        10'b0010000010: data <= 8'hff; 
        10'b0010000011: data <= 8'h00; 
        10'b0010000100: data <= 8'h00; 
        10'b0010000101: data <= 8'h00; 
        10'b0010000110: data <= 8'h00; 
        10'b0010000111: data <= 8'h00; 
        10'b0010001000: data <= 8'h00; 
        10'b0010001001: data <= 8'h00; 
        10'b0010001010: data <= 8'h00; 
        10'b0010001011: data <= 8'h00; 
        10'b0010001100: data <= 8'h00; 
        10'b0010001101: data <= 8'h00; 
        10'b0010001110: data <= 8'h00; 
        10'b0010001111: data <= 8'h00; 
        10'b0010010000: data <= 8'h00; 
        10'b0010010001: data <= 8'h00; 
        10'b0010010010: data <= 8'h00; 
        10'b0010010011: data <= 8'h00; 
        10'b0010010100: data <= 8'h00; 
        10'b0010010101: data <= 8'h00; 
        10'b0010010110: data <= 8'h00; 
        10'b0010010111: data <= 8'h00; 
        10'b0010011000: data <= 8'hff; 
        10'b0010011001: data <= 8'hff; 
        10'b0010011010: data <= 8'hff; 
        10'b0010011011: data <= 8'hff; 
        10'b0010011100: data <= 8'hfe; 
        10'b0010011101: data <= 8'hff; 
        10'b0010011110: data <= 8'hff; 
        10'b0010011111: data <= 8'h00; 
        10'b0010100000: data <= 8'h00; 
        10'b0010100001: data <= 8'h00; 
        10'b0010100010: data <= 8'h00; 
        10'b0010100011: data <= 8'h00; 
        10'b0010100100: data <= 8'h00; 
        10'b0010100101: data <= 8'h00; 
        10'b0010100110: data <= 8'h00; 
        10'b0010100111: data <= 8'h00; 
        10'b0010101000: data <= 8'h00; 
        10'b0010101001: data <= 8'h00; 
        10'b0010101010: data <= 8'h00; 
        10'b0010101011: data <= 8'h00; 
        10'b0010101100: data <= 8'h00; 
        10'b0010101101: data <= 8'h00; 
        10'b0010101110: data <= 8'h00; 
        10'b0010101111: data <= 8'hff; 
        10'b0010110000: data <= 8'hff; 
        10'b0010110001: data <= 8'hff; 
        10'b0010110010: data <= 8'hff; 
        10'b0010110011: data <= 8'h00; 
        10'b0010110100: data <= 8'h00; 
        10'b0010110101: data <= 8'h01; 
        10'b0010110110: data <= 8'h01; 
        10'b0010110111: data <= 8'h01; 
        10'b0010111000: data <= 8'h01; 
        10'b0010111001: data <= 8'h00; 
        10'b0010111010: data <= 8'h01; 
        10'b0010111011: data <= 8'h00; 
        10'b0010111100: data <= 8'h00; 
        10'b0010111101: data <= 8'h00; 
        10'b0010111110: data <= 8'hff; 
        10'b0010111111: data <= 8'hff; 
        10'b0011000000: data <= 8'h00; 
        10'b0011000001: data <= 8'h00; 
        10'b0011000010: data <= 8'h00; 
        10'b0011000011: data <= 8'h00; 
        10'b0011000100: data <= 8'h00; 
        10'b0011000101: data <= 8'h00; 
        10'b0011000110: data <= 8'h00; 
        10'b0011000111: data <= 8'h00; 
        10'b0011001000: data <= 8'h00; 
        10'b0011001001: data <= 8'hff; 
        10'b0011001010: data <= 8'hff; 
        10'b0011001011: data <= 8'hff; 
        10'b0011001100: data <= 8'hff; 
        10'b0011001101: data <= 8'h00; 
        10'b0011001110: data <= 8'h00; 
        10'b0011001111: data <= 8'h00; 
        10'b0011010000: data <= 8'h01; 
        10'b0011010001: data <= 8'h01; 
        10'b0011010010: data <= 8'h01; 
        10'b0011010011: data <= 8'h02; 
        10'b0011010100: data <= 8'h02; 
        10'b0011010101: data <= 8'h01; 
        10'b0011010110: data <= 8'h01; 
        10'b0011010111: data <= 8'h00; 
        10'b0011011000: data <= 8'h00; 
        10'b0011011001: data <= 8'h00; 
        10'b0011011010: data <= 8'hff; 
        10'b0011011011: data <= 8'hff; 
        10'b0011011100: data <= 8'hff; 
        10'b0011011101: data <= 8'h00; 
        10'b0011011110: data <= 8'h00; 
        10'b0011011111: data <= 8'h00; 
        10'b0011100000: data <= 8'h00; 
        10'b0011100001: data <= 8'h00; 
        10'b0011100010: data <= 8'h00; 
        10'b0011100011: data <= 8'h00; 
        10'b0011100100: data <= 8'h00; 
        10'b0011100101: data <= 8'hff; 
        10'b0011100110: data <= 8'hff; 
        10'b0011100111: data <= 8'hff; 
        10'b0011101000: data <= 8'h00; 
        10'b0011101001: data <= 8'h00; 
        10'b0011101010: data <= 8'h00; 
        10'b0011101011: data <= 8'h00; 
        10'b0011101100: data <= 8'h00; 
        10'b0011101101: data <= 8'h00; 
        10'b0011101110: data <= 8'h01; 
        10'b0011101111: data <= 8'h01; 
        10'b0011110000: data <= 8'h01; 
        10'b0011110001: data <= 8'h00; 
        10'b0011110010: data <= 8'h00; 
        10'b0011110011: data <= 8'h00; 
        10'b0011110100: data <= 8'h00; 
        10'b0011110101: data <= 8'h00; 
        10'b0011110110: data <= 8'h00; 
        10'b0011110111: data <= 8'hff; 
        10'b0011111000: data <= 8'hff; 
        10'b0011111001: data <= 8'h00; 
        10'b0011111010: data <= 8'h00; 
        10'b0011111011: data <= 8'h00; 
        10'b0011111100: data <= 8'h00; 
        10'b0011111101: data <= 8'h00; 
        10'b0011111110: data <= 8'h00; 
        10'b0011111111: data <= 8'h00; 
        10'b0100000000: data <= 8'hff; 
        10'b0100000001: data <= 8'hff; 
        10'b0100000010: data <= 8'h00; 
        10'b0100000011: data <= 8'h00; 
        10'b0100000100: data <= 8'h00; 
        10'b0100000101: data <= 8'h00; 
        10'b0100000110: data <= 8'h00; 
        10'b0100000111: data <= 8'h00; 
        10'b0100001000: data <= 8'h00; 
        10'b0100001001: data <= 8'h01; 
        10'b0100001010: data <= 8'h01; 
        10'b0100001011: data <= 8'h01; 
        10'b0100001100: data <= 8'h00; 
        10'b0100001101: data <= 8'h00; 
        10'b0100001110: data <= 8'h00; 
        10'b0100001111: data <= 8'h00; 
        10'b0100010000: data <= 8'h00; 
        10'b0100010001: data <= 8'h00; 
        10'b0100010010: data <= 8'hff; 
        10'b0100010011: data <= 8'hff; 
        10'b0100010100: data <= 8'h00; 
        10'b0100010101: data <= 8'h00; 
        10'b0100010110: data <= 8'h00; 
        10'b0100010111: data <= 8'h00; 
        10'b0100011000: data <= 8'h00; 
        10'b0100011001: data <= 8'h00; 
        10'b0100011010: data <= 8'h00; 
        10'b0100011011: data <= 8'h00; 
        10'b0100011100: data <= 8'hff; 
        10'b0100011101: data <= 8'h00; 
        10'b0100011110: data <= 8'h00; 
        10'b0100011111: data <= 8'h00; 
        10'b0100100000: data <= 8'h01; 
        10'b0100100001: data <= 8'h01; 
        10'b0100100010: data <= 8'h01; 
        10'b0100100011: data <= 8'h01; 
        10'b0100100100: data <= 8'h00; 
        10'b0100100101: data <= 8'h00; 
        10'b0100100110: data <= 8'h00; 
        10'b0100100111: data <= 8'h00; 
        10'b0100101000: data <= 8'h00; 
        10'b0100101001: data <= 8'h00; 
        10'b0100101010: data <= 8'h00; 
        10'b0100101011: data <= 8'h00; 
        10'b0100101100: data <= 8'h00; 
        10'b0100101101: data <= 8'h00; 
        10'b0100101110: data <= 8'h00; 
        10'b0100101111: data <= 8'h00; 
        10'b0100110000: data <= 8'h00; 
        10'b0100110001: data <= 8'h00; 
        10'b0100110010: data <= 8'h00; 
        10'b0100110011: data <= 8'h00; 
        10'b0100110100: data <= 8'h00; 
        10'b0100110101: data <= 8'h00; 
        10'b0100110110: data <= 8'h00; 
        10'b0100110111: data <= 8'h00; 
        10'b0100111000: data <= 8'h00; 
        10'b0100111001: data <= 8'h00; 
        10'b0100111010: data <= 8'h01; 
        10'b0100111011: data <= 8'h01; 
        10'b0100111100: data <= 8'h01; 
        10'b0100111101: data <= 8'h01; 
        10'b0100111110: data <= 8'h01; 
        10'b0100111111: data <= 8'h01; 
        10'b0101000000: data <= 8'h00; 
        10'b0101000001: data <= 8'h00; 
        10'b0101000010: data <= 8'h00; 
        10'b0101000011: data <= 8'h00; 
        10'b0101000100: data <= 8'h00; 
        10'b0101000101: data <= 8'h01; 
        10'b0101000110: data <= 8'h01; 
        10'b0101000111: data <= 8'h01; 
        10'b0101001000: data <= 8'h01; 
        10'b0101001001: data <= 8'h01; 
        10'b0101001010: data <= 8'h00; 
        10'b0101001011: data <= 8'h00; 
        10'b0101001100: data <= 8'h00; 
        10'b0101001101: data <= 8'h00; 
        10'b0101001110: data <= 8'h00; 
        10'b0101001111: data <= 8'h00; 
        10'b0101010000: data <= 8'h00; 
        10'b0101010001: data <= 8'h00; 
        10'b0101010010: data <= 8'h00; 
        10'b0101010011: data <= 8'h00; 
        10'b0101010100: data <= 8'h00; 
        10'b0101010101: data <= 8'h01; 
        10'b0101010110: data <= 8'h01; 
        10'b0101010111: data <= 8'h01; 
        10'b0101011000: data <= 8'h01; 
        10'b0101011001: data <= 8'h01; 
        10'b0101011010: data <= 8'h01; 
        10'b0101011011: data <= 8'h00; 
        10'b0101011100: data <= 8'hff; 
        10'b0101011101: data <= 8'h01; 
        10'b0101011110: data <= 8'h01; 
        10'b0101011111: data <= 8'h01; 
        10'b0101100000: data <= 8'h01; 
        10'b0101100001: data <= 8'h01; 
        10'b0101100010: data <= 8'h01; 
        10'b0101100011: data <= 8'h01; 
        10'b0101100100: data <= 8'h02; 
        10'b0101100101: data <= 8'h01; 
        10'b0101100110: data <= 8'h00; 
        10'b0101100111: data <= 8'h00; 
        10'b0101101000: data <= 8'h00; 
        10'b0101101001: data <= 8'h00; 
        10'b0101101010: data <= 8'h00; 
        10'b0101101011: data <= 8'h00; 
        10'b0101101100: data <= 8'h00; 
        10'b0101101101: data <= 8'h00; 
        10'b0101101110: data <= 8'h00; 
        10'b0101101111: data <= 8'h00; 
        10'b0101110000: data <= 8'h01; 
        10'b0101110001: data <= 8'h01; 
        10'b0101110010: data <= 8'h01; 
        10'b0101110011: data <= 8'h01; 
        10'b0101110100: data <= 8'h01; 
        10'b0101110101: data <= 8'h00; 
        10'b0101110110: data <= 8'h00; 
        10'b0101110111: data <= 8'h00; 
        10'b0101111000: data <= 8'h00; 
        10'b0101111001: data <= 8'h01; 
        10'b0101111010: data <= 8'h01; 
        10'b0101111011: data <= 8'h01; 
        10'b0101111100: data <= 8'h01; 
        10'b0101111101: data <= 8'h01; 
        10'b0101111110: data <= 8'h01; 
        10'b0101111111: data <= 8'h01; 
        10'b0110000000: data <= 8'h01; 
        10'b0110000001: data <= 8'h01; 
        10'b0110000010: data <= 8'h00; 
        10'b0110000011: data <= 8'h00; 
        10'b0110000100: data <= 8'h00; 
        10'b0110000101: data <= 8'h00; 
        10'b0110000110: data <= 8'h00; 
        10'b0110000111: data <= 8'h00; 
        10'b0110001000: data <= 8'h00; 
        10'b0110001001: data <= 8'h00; 
        10'b0110001010: data <= 8'h00; 
        10'b0110001011: data <= 8'h00; 
        10'b0110001100: data <= 8'h00; 
        10'b0110001101: data <= 8'h00; 
        10'b0110001110: data <= 8'h01; 
        10'b0110001111: data <= 8'h01; 
        10'b0110010000: data <= 8'h00; 
        10'b0110010001: data <= 8'h00; 
        10'b0110010010: data <= 8'h00; 
        10'b0110010011: data <= 8'h00; 
        10'b0110010100: data <= 8'h00; 
        10'b0110010101: data <= 8'h00; 
        10'b0110010110: data <= 8'h00; 
        10'b0110010111: data <= 8'h01; 
        10'b0110011000: data <= 8'h01; 
        10'b0110011001: data <= 8'h01; 
        10'b0110011010: data <= 8'h01; 
        10'b0110011011: data <= 8'h00; 
        10'b0110011100: data <= 8'h01; 
        10'b0110011101: data <= 8'h00; 
        10'b0110011110: data <= 8'hff; 
        10'b0110011111: data <= 8'hff; 
        10'b0110100000: data <= 8'h00; 
        10'b0110100001: data <= 8'h00; 
        10'b0110100010: data <= 8'h00; 
        10'b0110100011: data <= 8'h00; 
        10'b0110100100: data <= 8'h00; 
        10'b0110100101: data <= 8'h00; 
        10'b0110100110: data <= 8'h00; 
        10'b0110100111: data <= 8'h00; 
        10'b0110101000: data <= 8'h00; 
        10'b0110101001: data <= 8'h00; 
        10'b0110101010: data <= 8'h00; 
        10'b0110101011: data <= 8'h00; 
        10'b0110101100: data <= 8'h00; 
        10'b0110101101: data <= 8'h00; 
        10'b0110101110: data <= 8'h00; 
        10'b0110101111: data <= 8'h00; 
        10'b0110110000: data <= 8'h00; 
        10'b0110110001: data <= 8'h00; 
        10'b0110110010: data <= 8'h00; 
        10'b0110110011: data <= 8'h01; 
        10'b0110110100: data <= 8'h01; 
        10'b0110110101: data <= 8'h01; 
        10'b0110110110: data <= 8'h01; 
        10'b0110110111: data <= 8'h00; 
        10'b0110111000: data <= 8'h00; 
        10'b0110111001: data <= 8'hff; 
        10'b0110111010: data <= 8'hff; 
        10'b0110111011: data <= 8'hff; 
        10'b0110111100: data <= 8'h00; 
        10'b0110111101: data <= 8'h00; 
        10'b0110111110: data <= 8'h00; 
        10'b0110111111: data <= 8'h00; 
        10'b0111000000: data <= 8'h00; 
        10'b0111000001: data <= 8'h00; 
        10'b0111000010: data <= 8'h00; 
        10'b0111000011: data <= 8'h00; 
        10'b0111000100: data <= 8'h00; 
        10'b0111000101: data <= 8'h00; 
        10'b0111000110: data <= 8'h00; 
        10'b0111000111: data <= 8'h00; 
        10'b0111001000: data <= 8'h01; 
        10'b0111001001: data <= 8'h00; 
        10'b0111001010: data <= 8'h00; 
        10'b0111001011: data <= 8'h00; 
        10'b0111001100: data <= 8'h00; 
        10'b0111001101: data <= 8'hff; 
        10'b0111001110: data <= 8'h00; 
        10'b0111001111: data <= 8'h01; 
        10'b0111010000: data <= 8'h01; 
        10'b0111010001: data <= 8'h01; 
        10'b0111010010: data <= 8'h00; 
        10'b0111010011: data <= 8'hff; 
        10'b0111010100: data <= 8'hff; 
        10'b0111010101: data <= 8'hff; 
        10'b0111010110: data <= 8'hff; 
        10'b0111010111: data <= 8'hff; 
        10'b0111011000: data <= 8'h00; 
        10'b0111011001: data <= 8'h00; 
        10'b0111011010: data <= 8'h00; 
        10'b0111011011: data <= 8'h00; 
        10'b0111011100: data <= 8'h00; 
        10'b0111011101: data <= 8'h00; 
        10'b0111011110: data <= 8'h00; 
        10'b0111011111: data <= 8'h00; 
        10'b0111100000: data <= 8'h00; 
        10'b0111100001: data <= 8'h00; 
        10'b0111100010: data <= 8'h00; 
        10'b0111100011: data <= 8'h00; 
        10'b0111100100: data <= 8'h00; 
        10'b0111100101: data <= 8'h00; 
        10'b0111100110: data <= 8'h01; 
        10'b0111100111: data <= 8'h01; 
        10'b0111101000: data <= 8'h00; 
        10'b0111101001: data <= 8'h00; 
        10'b0111101010: data <= 8'h00; 
        10'b0111101011: data <= 8'h01; 
        10'b0111101100: data <= 8'h00; 
        10'b0111101101: data <= 8'h00; 
        10'b0111101110: data <= 8'h00; 
        10'b0111101111: data <= 8'hff; 
        10'b0111110000: data <= 8'hff; 
        10'b0111110001: data <= 8'hff; 
        10'b0111110010: data <= 8'hff; 
        10'b0111110011: data <= 8'hff; 
        10'b0111110100: data <= 8'h00; 
        10'b0111110101: data <= 8'h00; 
        10'b0111110110: data <= 8'h00; 
        10'b0111110111: data <= 8'h00; 
        10'b0111111000: data <= 8'h00; 
        10'b0111111001: data <= 8'h00; 
        10'b0111111010: data <= 8'h00; 
        10'b0111111011: data <= 8'h00; 
        10'b0111111100: data <= 8'h00; 
        10'b0111111101: data <= 8'hff; 
        10'b0111111110: data <= 8'hff; 
        10'b0111111111: data <= 8'hff; 
        10'b1000000000: data <= 8'h00; 
        10'b1000000001: data <= 8'h00; 
        10'b1000000010: data <= 8'h01; 
        10'b1000000011: data <= 8'h01; 
        10'b1000000100: data <= 8'h00; 
        10'b1000000101: data <= 8'h00; 
        10'b1000000110: data <= 8'h00; 
        10'b1000000111: data <= 8'h01; 
        10'b1000001000: data <= 8'h00; 
        10'b1000001001: data <= 8'h00; 
        10'b1000001010: data <= 8'hff; 
        10'b1000001011: data <= 8'h00; 
        10'b1000001100: data <= 8'h00; 
        10'b1000001101: data <= 8'hff; 
        10'b1000001110: data <= 8'hff; 
        10'b1000001111: data <= 8'hff; 
        10'b1000010000: data <= 8'h00; 
        10'b1000010001: data <= 8'h00; 
        10'b1000010010: data <= 8'h00; 
        10'b1000010011: data <= 8'h00; 
        10'b1000010100: data <= 8'h00; 
        10'b1000010101: data <= 8'h00; 
        10'b1000010110: data <= 8'h00; 
        10'b1000010111: data <= 8'h00; 
        10'b1000011000: data <= 8'h00; 
        10'b1000011001: data <= 8'hff; 
        10'b1000011010: data <= 8'hff; 
        10'b1000011011: data <= 8'hff; 
        10'b1000011100: data <= 8'hff; 
        10'b1000011101: data <= 8'hff; 
        10'b1000011110: data <= 8'hff; 
        10'b1000011111: data <= 8'hff; 
        10'b1000100000: data <= 8'hff; 
        10'b1000100001: data <= 8'hff; 
        10'b1000100010: data <= 8'hff; 
        10'b1000100011: data <= 8'hff; 
        10'b1000100100: data <= 8'hff; 
        10'b1000100101: data <= 8'h00; 
        10'b1000100110: data <= 8'h00; 
        10'b1000100111: data <= 8'h00; 
        10'b1000101000: data <= 8'h00; 
        10'b1000101001: data <= 8'h00; 
        10'b1000101010: data <= 8'h00; 
        10'b1000101011: data <= 8'h00; 
        10'b1000101100: data <= 8'h00; 
        10'b1000101101: data <= 8'h00; 
        10'b1000101110: data <= 8'h00; 
        10'b1000101111: data <= 8'h00; 
        10'b1000110000: data <= 8'h00; 
        10'b1000110001: data <= 8'h00; 
        10'b1000110010: data <= 8'h00; 
        10'b1000110011: data <= 8'h00; 
        10'b1000110100: data <= 8'h00; 
        10'b1000110101: data <= 8'h00; 
        10'b1000110110: data <= 8'hff; 
        10'b1000110111: data <= 8'hff; 
        10'b1000111000: data <= 8'hff; 
        10'b1000111001: data <= 8'hff; 
        10'b1000111010: data <= 8'hfe; 
        10'b1000111011: data <= 8'hfe; 
        10'b1000111100: data <= 8'hff; 
        10'b1000111101: data <= 8'h00; 
        10'b1000111110: data <= 8'hff; 
        10'b1000111111: data <= 8'h00; 
        10'b1001000000: data <= 8'h00; 
        10'b1001000001: data <= 8'h00; 
        10'b1001000010: data <= 8'hff; 
        10'b1001000011: data <= 8'h00; 
        10'b1001000100: data <= 8'h00; 
        10'b1001000101: data <= 8'h00; 
        10'b1001000110: data <= 8'h00; 
        10'b1001000111: data <= 8'h00; 
        10'b1001001000: data <= 8'h00; 
        10'b1001001001: data <= 8'h00; 
        10'b1001001010: data <= 8'h00; 
        10'b1001001011: data <= 8'h00; 
        10'b1001001100: data <= 8'h00; 
        10'b1001001101: data <= 8'h00; 
        10'b1001001110: data <= 8'h00; 
        10'b1001001111: data <= 8'h00; 
        10'b1001010000: data <= 8'h00; 
        10'b1001010001: data <= 8'h00; 
        10'b1001010010: data <= 8'hff; 
        10'b1001010011: data <= 8'hff; 
        10'b1001010100: data <= 8'hff; 
        10'b1001010101: data <= 8'hff; 
        10'b1001010110: data <= 8'hff; 
        10'b1001010111: data <= 8'hff; 
        10'b1001011000: data <= 8'hff; 
        10'b1001011001: data <= 8'hff; 
        10'b1001011010: data <= 8'hff; 
        10'b1001011011: data <= 8'h00; 
        10'b1001011100: data <= 8'h00; 
        10'b1001011101: data <= 8'hff; 
        10'b1001011110: data <= 8'hff; 
        10'b1001011111: data <= 8'h00; 
        10'b1001100000: data <= 8'h00; 
        10'b1001100001: data <= 8'h00; 
        10'b1001100010: data <= 8'h00; 
        10'b1001100011: data <= 8'h00; 
        10'b1001100100: data <= 8'h00; 
        10'b1001100101: data <= 8'h00; 
        10'b1001100110: data <= 8'h00; 
        10'b1001100111: data <= 8'h00; 
        10'b1001101000: data <= 8'h00; 
        10'b1001101001: data <= 8'h00; 
        10'b1001101010: data <= 8'h00; 
        10'b1001101011: data <= 8'h00; 
        10'b1001101100: data <= 8'h00; 
        10'b1001101101: data <= 8'h00; 
        10'b1001101110: data <= 8'hff; 
        10'b1001101111: data <= 8'hff; 
        10'b1001110000: data <= 8'hff; 
        10'b1001110001: data <= 8'hff; 
        10'b1001110010: data <= 8'hff; 
        10'b1001110011: data <= 8'h00; 
        10'b1001110100: data <= 8'hff; 
        10'b1001110101: data <= 8'hff; 
        10'b1001110110: data <= 8'hff; 
        10'b1001110111: data <= 8'hff; 
        10'b1001111000: data <= 8'hff; 
        10'b1001111001: data <= 8'hff; 
        10'b1001111010: data <= 8'hff; 
        10'b1001111011: data <= 8'hff; 
        10'b1001111100: data <= 8'h00; 
        10'b1001111101: data <= 8'h00; 
        10'b1001111110: data <= 8'h00; 
        10'b1001111111: data <= 8'h00; 
        10'b1010000000: data <= 8'h00; 
        10'b1010000001: data <= 8'h00; 
        10'b1010000010: data <= 8'h00; 
        10'b1010000011: data <= 8'h00; 
        10'b1010000100: data <= 8'h00; 
        10'b1010000101: data <= 8'h00; 
        10'b1010000110: data <= 8'h00; 
        10'b1010000111: data <= 8'h00; 
        10'b1010001000: data <= 8'h00; 
        10'b1010001001: data <= 8'h00; 
        10'b1010001010: data <= 8'h00; 
        10'b1010001011: data <= 8'hff; 
        10'b1010001100: data <= 8'h00; 
        10'b1010001101: data <= 8'h00; 
        10'b1010001110: data <= 8'h00; 
        10'b1010001111: data <= 8'hff; 
        10'b1010010000: data <= 8'hff; 
        10'b1010010001: data <= 8'hff; 
        10'b1010010010: data <= 8'hff; 
        10'b1010010011: data <= 8'hff; 
        10'b1010010100: data <= 8'hff; 
        10'b1010010101: data <= 8'hff; 
        10'b1010010110: data <= 8'hff; 
        10'b1010010111: data <= 8'h00; 
        10'b1010011000: data <= 8'h00; 
        10'b1010011001: data <= 8'h00; 
        10'b1010011010: data <= 8'h01; 
        10'b1010011011: data <= 8'h01; 
        10'b1010011100: data <= 8'h00; 
        10'b1010011101: data <= 8'h00; 
        10'b1010011110: data <= 8'h00; 
        10'b1010011111: data <= 8'h00; 
        10'b1010100000: data <= 8'h00; 
        10'b1010100001: data <= 8'h00; 
        10'b1010100010: data <= 8'h00; 
        10'b1010100011: data <= 8'h00; 
        10'b1010100100: data <= 8'h00; 
        10'b1010100101: data <= 8'h00; 
        10'b1010100110: data <= 8'h00; 
        10'b1010100111: data <= 8'h00; 
        10'b1010101000: data <= 8'h00; 
        10'b1010101001: data <= 8'h00; 
        10'b1010101010: data <= 8'h00; 
        10'b1010101011: data <= 8'h00; 
        10'b1010101100: data <= 8'h00; 
        10'b1010101101: data <= 8'h00; 
        10'b1010101110: data <= 8'hff; 
        10'b1010101111: data <= 8'hff; 
        10'b1010110000: data <= 8'h00; 
        10'b1010110001: data <= 8'h00; 
        10'b1010110010: data <= 8'h00; 
        10'b1010110011: data <= 8'h00; 
        10'b1010110100: data <= 8'h01; 
        10'b1010110101: data <= 8'h01; 
        10'b1010110110: data <= 8'h01; 
        10'b1010110111: data <= 8'h00; 
        10'b1010111000: data <= 8'h00; 
        10'b1010111001: data <= 8'h00; 
        10'b1010111010: data <= 8'h00; 
        10'b1010111011: data <= 8'h00; 
        10'b1010111100: data <= 8'h00; 
        10'b1010111101: data <= 8'h00; 
        10'b1010111110: data <= 8'h00; 
        10'b1010111111: data <= 8'h00; 
        10'b1011000000: data <= 8'h00; 
        10'b1011000001: data <= 8'h00; 
        10'b1011000010: data <= 8'h00; 
        10'b1011000011: data <= 8'h01; 
        10'b1011000100: data <= 8'h01; 
        10'b1011000101: data <= 8'h01; 
        10'b1011000110: data <= 8'h01; 
        10'b1011000111: data <= 8'h00; 
        10'b1011001000: data <= 8'h01; 
        10'b1011001001: data <= 8'h01; 
        10'b1011001010: data <= 8'h01; 
        10'b1011001011: data <= 8'h01; 
        10'b1011001100: data <= 8'h01; 
        10'b1011001101: data <= 8'h01; 
        10'b1011001110: data <= 8'h01; 
        10'b1011001111: data <= 8'h01; 
        10'b1011010000: data <= 8'h01; 
        10'b1011010001: data <= 8'h01; 
        10'b1011010010: data <= 8'h00; 
        10'b1011010011: data <= 8'h00; 
        10'b1011010100: data <= 8'h00; 
        10'b1011010101: data <= 8'h00; 
        10'b1011010110: data <= 8'h00; 
        10'b1011010111: data <= 8'h00; 
        10'b1011011000: data <= 8'h00; 
        10'b1011011001: data <= 8'h00; 
        10'b1011011010: data <= 8'h00; 
        10'b1011011011: data <= 8'h00; 
        10'b1011011100: data <= 8'h00; 
        10'b1011011101: data <= 8'h00; 
        10'b1011011110: data <= 8'h00; 
        10'b1011011111: data <= 8'h00; 
        10'b1011100000: data <= 8'h01; 
        10'b1011100001: data <= 8'h01; 
        10'b1011100010: data <= 8'h01; 
        10'b1011100011: data <= 8'h01; 
        10'b1011100100: data <= 8'h01; 
        10'b1011100101: data <= 8'h01; 
        10'b1011100110: data <= 8'h01; 
        10'b1011100111: data <= 8'h01; 
        10'b1011101000: data <= 8'h01; 
        10'b1011101001: data <= 8'h00; 
        10'b1011101010: data <= 8'h01; 
        10'b1011101011: data <= 8'h01; 
        10'b1011101100: data <= 8'h01; 
        10'b1011101101: data <= 8'h00; 
        10'b1011101110: data <= 8'h00; 
        10'b1011101111: data <= 8'h00; 
        10'b1011110000: data <= 8'h00; 
        10'b1011110001: data <= 8'h00; 
        10'b1011110010: data <= 8'h00; 
        10'b1011110011: data <= 8'h00; 
        10'b1011110100: data <= 8'h00; 
        10'b1011110101: data <= 8'h00; 
        10'b1011110110: data <= 8'h00; 
        10'b1011110111: data <= 8'h00; 
        10'b1011111000: data <= 8'h00; 
        10'b1011111001: data <= 8'h00; 
        10'b1011111010: data <= 8'h00; 
        10'b1011111011: data <= 8'h00; 
        10'b1011111100: data <= 8'h00; 
        10'b1011111101: data <= 8'h00; 
        10'b1011111110: data <= 8'h00; 
        10'b1011111111: data <= 8'h00; 
        10'b1100000000: data <= 8'h00; 
        10'b1100000001: data <= 8'h00; 
        10'b1100000010: data <= 8'h00; 
        10'b1100000011: data <= 8'h00; 
        10'b1100000100: data <= 8'h00; 
        10'b1100000101: data <= 8'h00; 
        10'b1100000110: data <= 8'h00; 
        10'b1100000111: data <= 8'h00; 
        10'b1100001000: data <= 8'h00; 
        10'b1100001001: data <= 8'h00; 
        10'b1100001010: data <= 8'h00; 
        10'b1100001011: data <= 8'h00; 
        10'b1100001100: data <= 8'h00; 
        10'b1100001101: data <= 8'h00; 
        10'b1100001110: data <= 8'h00; 
        10'b1100001111: data <= 8'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 3) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 9'h000; 
        10'b0000000001: data <= 9'h000; 
        10'b0000000010: data <= 9'h000; 
        10'b0000000011: data <= 9'h000; 
        10'b0000000100: data <= 9'h000; 
        10'b0000000101: data <= 9'h000; 
        10'b0000000110: data <= 9'h000; 
        10'b0000000111: data <= 9'h000; 
        10'b0000001000: data <= 9'h000; 
        10'b0000001001: data <= 9'h000; 
        10'b0000001010: data <= 9'h000; 
        10'b0000001011: data <= 9'h000; 
        10'b0000001100: data <= 9'h000; 
        10'b0000001101: data <= 9'h000; 
        10'b0000001110: data <= 9'h000; 
        10'b0000001111: data <= 9'h000; 
        10'b0000010000: data <= 9'h000; 
        10'b0000010001: data <= 9'h000; 
        10'b0000010010: data <= 9'h000; 
        10'b0000010011: data <= 9'h000; 
        10'b0000010100: data <= 9'h000; 
        10'b0000010101: data <= 9'h000; 
        10'b0000010110: data <= 9'h000; 
        10'b0000010111: data <= 9'h000; 
        10'b0000011000: data <= 9'h000; 
        10'b0000011001: data <= 9'h000; 
        10'b0000011010: data <= 9'h000; 
        10'b0000011011: data <= 9'h000; 
        10'b0000011100: data <= 9'h000; 
        10'b0000011101: data <= 9'h000; 
        10'b0000011110: data <= 9'h000; 
        10'b0000011111: data <= 9'h000; 
        10'b0000100000: data <= 9'h000; 
        10'b0000100001: data <= 9'h000; 
        10'b0000100010: data <= 9'h000; 
        10'b0000100011: data <= 9'h000; 
        10'b0000100100: data <= 9'h000; 
        10'b0000100101: data <= 9'h000; 
        10'b0000100110: data <= 9'h000; 
        10'b0000100111: data <= 9'h000; 
        10'b0000101000: data <= 9'h000; 
        10'b0000101001: data <= 9'h000; 
        10'b0000101010: data <= 9'h000; 
        10'b0000101011: data <= 9'h000; 
        10'b0000101100: data <= 9'h000; 
        10'b0000101101: data <= 9'h000; 
        10'b0000101110: data <= 9'h000; 
        10'b0000101111: data <= 9'h000; 
        10'b0000110000: data <= 9'h000; 
        10'b0000110001: data <= 9'h000; 
        10'b0000110010: data <= 9'h000; 
        10'b0000110011: data <= 9'h000; 
        10'b0000110100: data <= 9'h000; 
        10'b0000110101: data <= 9'h000; 
        10'b0000110110: data <= 9'h000; 
        10'b0000110111: data <= 9'h000; 
        10'b0000111000: data <= 9'h000; 
        10'b0000111001: data <= 9'h000; 
        10'b0000111010: data <= 9'h000; 
        10'b0000111011: data <= 9'h000; 
        10'b0000111100: data <= 9'h000; 
        10'b0000111101: data <= 9'h000; 
        10'b0000111110: data <= 9'h000; 
        10'b0000111111: data <= 9'h000; 
        10'b0001000000: data <= 9'h000; 
        10'b0001000001: data <= 9'h000; 
        10'b0001000010: data <= 9'h000; 
        10'b0001000011: data <= 9'h000; 
        10'b0001000100: data <= 9'h000; 
        10'b0001000101: data <= 9'h000; 
        10'b0001000110: data <= 9'h000; 
        10'b0001000111: data <= 9'h000; 
        10'b0001001000: data <= 9'h000; 
        10'b0001001001: data <= 9'h000; 
        10'b0001001010: data <= 9'h000; 
        10'b0001001011: data <= 9'h000; 
        10'b0001001100: data <= 9'h000; 
        10'b0001001101: data <= 9'h000; 
        10'b0001001110: data <= 9'h000; 
        10'b0001001111: data <= 9'h000; 
        10'b0001010000: data <= 9'h000; 
        10'b0001010001: data <= 9'h000; 
        10'b0001010010: data <= 9'h000; 
        10'b0001010011: data <= 9'h000; 
        10'b0001010100: data <= 9'h000; 
        10'b0001010101: data <= 9'h000; 
        10'b0001010110: data <= 9'h000; 
        10'b0001010111: data <= 9'h000; 
        10'b0001011000: data <= 9'h000; 
        10'b0001011001: data <= 9'h000; 
        10'b0001011010: data <= 9'h000; 
        10'b0001011011: data <= 9'h000; 
        10'b0001011100: data <= 9'h000; 
        10'b0001011101: data <= 9'h000; 
        10'b0001011110: data <= 9'h000; 
        10'b0001011111: data <= 9'h000; 
        10'b0001100000: data <= 9'h000; 
        10'b0001100001: data <= 9'h000; 
        10'b0001100010: data <= 9'h000; 
        10'b0001100011: data <= 9'h000; 
        10'b0001100100: data <= 9'h000; 
        10'b0001100101: data <= 9'h000; 
        10'b0001100110: data <= 9'h000; 
        10'b0001100111: data <= 9'h000; 
        10'b0001101000: data <= 9'h000; 
        10'b0001101001: data <= 9'h000; 
        10'b0001101010: data <= 9'h000; 
        10'b0001101011: data <= 9'h000; 
        10'b0001101100: data <= 9'h000; 
        10'b0001101101: data <= 9'h000; 
        10'b0001101110: data <= 9'h000; 
        10'b0001101111: data <= 9'h000; 
        10'b0001110000: data <= 9'h000; 
        10'b0001110001: data <= 9'h000; 
        10'b0001110010: data <= 9'h000; 
        10'b0001110011: data <= 9'h000; 
        10'b0001110100: data <= 9'h000; 
        10'b0001110101: data <= 9'h000; 
        10'b0001110110: data <= 9'h000; 
        10'b0001110111: data <= 9'h000; 
        10'b0001111000: data <= 9'h000; 
        10'b0001111001: data <= 9'h000; 
        10'b0001111010: data <= 9'h000; 
        10'b0001111011: data <= 9'h000; 
        10'b0001111100: data <= 9'h1ff; 
        10'b0001111101: data <= 9'h1ff; 
        10'b0001111110: data <= 9'h1fe; 
        10'b0001111111: data <= 9'h1fe; 
        10'b0010000000: data <= 9'h1fe; 
        10'b0010000001: data <= 9'h1fe; 
        10'b0010000010: data <= 9'h1ff; 
        10'b0010000011: data <= 9'h1ff; 
        10'b0010000100: data <= 9'h000; 
        10'b0010000101: data <= 9'h000; 
        10'b0010000110: data <= 9'h000; 
        10'b0010000111: data <= 9'h000; 
        10'b0010001000: data <= 9'h000; 
        10'b0010001001: data <= 9'h000; 
        10'b0010001010: data <= 9'h000; 
        10'b0010001011: data <= 9'h000; 
        10'b0010001100: data <= 9'h000; 
        10'b0010001101: data <= 9'h000; 
        10'b0010001110: data <= 9'h000; 
        10'b0010001111: data <= 9'h000; 
        10'b0010010000: data <= 9'h000; 
        10'b0010010001: data <= 9'h000; 
        10'b0010010010: data <= 9'h000; 
        10'b0010010011: data <= 9'h000; 
        10'b0010010100: data <= 9'h1ff; 
        10'b0010010101: data <= 9'h1ff; 
        10'b0010010110: data <= 9'h1ff; 
        10'b0010010111: data <= 9'h1ff; 
        10'b0010011000: data <= 9'h1ff; 
        10'b0010011001: data <= 9'h1ff; 
        10'b0010011010: data <= 9'h1fe; 
        10'b0010011011: data <= 9'h1fe; 
        10'b0010011100: data <= 9'h1fd; 
        10'b0010011101: data <= 9'h1fe; 
        10'b0010011110: data <= 9'h1ff; 
        10'b0010011111: data <= 9'h1ff; 
        10'b0010100000: data <= 9'h1ff; 
        10'b0010100001: data <= 9'h1ff; 
        10'b0010100010: data <= 9'h1ff; 
        10'b0010100011: data <= 9'h1ff; 
        10'b0010100100: data <= 9'h000; 
        10'b0010100101: data <= 9'h000; 
        10'b0010100110: data <= 9'h000; 
        10'b0010100111: data <= 9'h000; 
        10'b0010101000: data <= 9'h000; 
        10'b0010101001: data <= 9'h000; 
        10'b0010101010: data <= 9'h000; 
        10'b0010101011: data <= 9'h000; 
        10'b0010101100: data <= 9'h000; 
        10'b0010101101: data <= 9'h1ff; 
        10'b0010101110: data <= 9'h1ff; 
        10'b0010101111: data <= 9'h1ff; 
        10'b0010110000: data <= 9'h1ff; 
        10'b0010110001: data <= 9'h1ff; 
        10'b0010110010: data <= 9'h1ff; 
        10'b0010110011: data <= 9'h000; 
        10'b0010110100: data <= 9'h000; 
        10'b0010110101: data <= 9'h001; 
        10'b0010110110: data <= 9'h002; 
        10'b0010110111: data <= 9'h002; 
        10'b0010111000: data <= 9'h001; 
        10'b0010111001: data <= 9'h001; 
        10'b0010111010: data <= 9'h001; 
        10'b0010111011: data <= 9'h000; 
        10'b0010111100: data <= 9'h000; 
        10'b0010111101: data <= 9'h1ff; 
        10'b0010111110: data <= 9'h1fe; 
        10'b0010111111: data <= 9'h1fe; 
        10'b0011000000: data <= 9'h1ff; 
        10'b0011000001: data <= 9'h000; 
        10'b0011000010: data <= 9'h000; 
        10'b0011000011: data <= 9'h000; 
        10'b0011000100: data <= 9'h000; 
        10'b0011000101: data <= 9'h000; 
        10'b0011000110: data <= 9'h000; 
        10'b0011000111: data <= 9'h000; 
        10'b0011001000: data <= 9'h1ff; 
        10'b0011001001: data <= 9'h1ff; 
        10'b0011001010: data <= 9'h1fe; 
        10'b0011001011: data <= 9'h1fe; 
        10'b0011001100: data <= 9'h1fe; 
        10'b0011001101: data <= 9'h1ff; 
        10'b0011001110: data <= 9'h000; 
        10'b0011001111: data <= 9'h000; 
        10'b0011010000: data <= 9'h002; 
        10'b0011010001: data <= 9'h002; 
        10'b0011010010: data <= 9'h003; 
        10'b0011010011: data <= 9'h003; 
        10'b0011010100: data <= 9'h003; 
        10'b0011010101: data <= 9'h001; 
        10'b0011010110: data <= 9'h001; 
        10'b0011010111: data <= 9'h000; 
        10'b0011011000: data <= 9'h000; 
        10'b0011011001: data <= 9'h000; 
        10'b0011011010: data <= 9'h1ff; 
        10'b0011011011: data <= 9'h1fe; 
        10'b0011011100: data <= 9'h1ff; 
        10'b0011011101: data <= 9'h000; 
        10'b0011011110: data <= 9'h000; 
        10'b0011011111: data <= 9'h000; 
        10'b0011100000: data <= 9'h000; 
        10'b0011100001: data <= 9'h000; 
        10'b0011100010: data <= 9'h000; 
        10'b0011100011: data <= 9'h000; 
        10'b0011100100: data <= 9'h1ff; 
        10'b0011100101: data <= 9'h1ff; 
        10'b0011100110: data <= 9'h1fe; 
        10'b0011100111: data <= 9'h1fe; 
        10'b0011101000: data <= 9'h1ff; 
        10'b0011101001: data <= 9'h000; 
        10'b0011101010: data <= 9'h000; 
        10'b0011101011: data <= 9'h1ff; 
        10'b0011101100: data <= 9'h000; 
        10'b0011101101: data <= 9'h001; 
        10'b0011101110: data <= 9'h003; 
        10'b0011101111: data <= 9'h001; 
        10'b0011110000: data <= 9'h001; 
        10'b0011110001: data <= 9'h000; 
        10'b0011110010: data <= 9'h000; 
        10'b0011110011: data <= 9'h000; 
        10'b0011110100: data <= 9'h000; 
        10'b0011110101: data <= 9'h000; 
        10'b0011110110: data <= 9'h1ff; 
        10'b0011110111: data <= 9'h1fe; 
        10'b0011111000: data <= 9'h1ff; 
        10'b0011111001: data <= 9'h1ff; 
        10'b0011111010: data <= 9'h000; 
        10'b0011111011: data <= 9'h000; 
        10'b0011111100: data <= 9'h000; 
        10'b0011111101: data <= 9'h000; 
        10'b0011111110: data <= 9'h000; 
        10'b0011111111: data <= 9'h1ff; 
        10'b0100000000: data <= 9'h1ff; 
        10'b0100000001: data <= 9'h1ff; 
        10'b0100000010: data <= 9'h000; 
        10'b0100000011: data <= 9'h1ff; 
        10'b0100000100: data <= 9'h000; 
        10'b0100000101: data <= 9'h000; 
        10'b0100000110: data <= 9'h001; 
        10'b0100000111: data <= 9'h000; 
        10'b0100001000: data <= 9'h000; 
        10'b0100001001: data <= 9'h001; 
        10'b0100001010: data <= 9'h002; 
        10'b0100001011: data <= 9'h002; 
        10'b0100001100: data <= 9'h000; 
        10'b0100001101: data <= 9'h000; 
        10'b0100001110: data <= 9'h000; 
        10'b0100001111: data <= 9'h1ff; 
        10'b0100010000: data <= 9'h000; 
        10'b0100010001: data <= 9'h1ff; 
        10'b0100010010: data <= 9'h1ff; 
        10'b0100010011: data <= 9'h1ff; 
        10'b0100010100: data <= 9'h1ff; 
        10'b0100010101: data <= 9'h000; 
        10'b0100010110: data <= 9'h000; 
        10'b0100010111: data <= 9'h000; 
        10'b0100011000: data <= 9'h000; 
        10'b0100011001: data <= 9'h000; 
        10'b0100011010: data <= 9'h000; 
        10'b0100011011: data <= 9'h000; 
        10'b0100011100: data <= 9'h1ff; 
        10'b0100011101: data <= 9'h1ff; 
        10'b0100011110: data <= 9'h001; 
        10'b0100011111: data <= 9'h001; 
        10'b0100100000: data <= 9'h001; 
        10'b0100100001: data <= 9'h001; 
        10'b0100100010: data <= 9'h001; 
        10'b0100100011: data <= 9'h002; 
        10'b0100100100: data <= 9'h001; 
        10'b0100100101: data <= 9'h000; 
        10'b0100100110: data <= 9'h000; 
        10'b0100100111: data <= 9'h1ff; 
        10'b0100101000: data <= 9'h1ff; 
        10'b0100101001: data <= 9'h000; 
        10'b0100101010: data <= 9'h001; 
        10'b0100101011: data <= 9'h000; 
        10'b0100101100: data <= 9'h001; 
        10'b0100101101: data <= 9'h000; 
        10'b0100101110: data <= 9'h1ff; 
        10'b0100101111: data <= 9'h1ff; 
        10'b0100110000: data <= 9'h1ff; 
        10'b0100110001: data <= 9'h000; 
        10'b0100110010: data <= 9'h000; 
        10'b0100110011: data <= 9'h000; 
        10'b0100110100: data <= 9'h000; 
        10'b0100110101: data <= 9'h000; 
        10'b0100110110: data <= 9'h000; 
        10'b0100110111: data <= 9'h000; 
        10'b0100111000: data <= 9'h000; 
        10'b0100111001: data <= 9'h001; 
        10'b0100111010: data <= 9'h002; 
        10'b0100111011: data <= 9'h002; 
        10'b0100111100: data <= 9'h003; 
        10'b0100111101: data <= 9'h001; 
        10'b0100111110: data <= 9'h001; 
        10'b0100111111: data <= 9'h002; 
        10'b0101000000: data <= 9'h1ff; 
        10'b0101000001: data <= 9'h1ff; 
        10'b0101000010: data <= 9'h000; 
        10'b0101000011: data <= 9'h000; 
        10'b0101000100: data <= 9'h001; 
        10'b0101000101: data <= 9'h003; 
        10'b0101000110: data <= 9'h001; 
        10'b0101000111: data <= 9'h001; 
        10'b0101001000: data <= 9'h002; 
        10'b0101001001: data <= 9'h001; 
        10'b0101001010: data <= 9'h001; 
        10'b0101001011: data <= 9'h000; 
        10'b0101001100: data <= 9'h000; 
        10'b0101001101: data <= 9'h000; 
        10'b0101001110: data <= 9'h000; 
        10'b0101001111: data <= 9'h000; 
        10'b0101010000: data <= 9'h000; 
        10'b0101010001: data <= 9'h000; 
        10'b0101010010: data <= 9'h000; 
        10'b0101010011: data <= 9'h000; 
        10'b0101010100: data <= 9'h001; 
        10'b0101010101: data <= 9'h002; 
        10'b0101010110: data <= 9'h003; 
        10'b0101010111: data <= 9'h001; 
        10'b0101011000: data <= 9'h002; 
        10'b0101011001: data <= 9'h002; 
        10'b0101011010: data <= 9'h001; 
        10'b0101011011: data <= 9'h000; 
        10'b0101011100: data <= 9'h1ff; 
        10'b0101011101: data <= 9'h001; 
        10'b0101011110: data <= 9'h003; 
        10'b0101011111: data <= 9'h002; 
        10'b0101100000: data <= 9'h002; 
        10'b0101100001: data <= 9'h003; 
        10'b0101100010: data <= 9'h003; 
        10'b0101100011: data <= 9'h003; 
        10'b0101100100: data <= 9'h003; 
        10'b0101100101: data <= 9'h002; 
        10'b0101100110: data <= 9'h001; 
        10'b0101100111: data <= 9'h000; 
        10'b0101101000: data <= 9'h000; 
        10'b0101101001: data <= 9'h000; 
        10'b0101101010: data <= 9'h000; 
        10'b0101101011: data <= 9'h000; 
        10'b0101101100: data <= 9'h000; 
        10'b0101101101: data <= 9'h000; 
        10'b0101101110: data <= 9'h000; 
        10'b0101101111: data <= 9'h000; 
        10'b0101110000: data <= 9'h001; 
        10'b0101110001: data <= 9'h002; 
        10'b0101110010: data <= 9'h002; 
        10'b0101110011: data <= 9'h001; 
        10'b0101110100: data <= 9'h001; 
        10'b0101110101: data <= 9'h001; 
        10'b0101110110: data <= 9'h001; 
        10'b0101110111: data <= 9'h000; 
        10'b0101111000: data <= 9'h1ff; 
        10'b0101111001: data <= 9'h002; 
        10'b0101111010: data <= 9'h003; 
        10'b0101111011: data <= 9'h002; 
        10'b0101111100: data <= 9'h002; 
        10'b0101111101: data <= 9'h002; 
        10'b0101111110: data <= 9'h003; 
        10'b0101111111: data <= 9'h003; 
        10'b0110000000: data <= 9'h002; 
        10'b0110000001: data <= 9'h001; 
        10'b0110000010: data <= 9'h000; 
        10'b0110000011: data <= 9'h1ff; 
        10'b0110000100: data <= 9'h1ff; 
        10'b0110000101: data <= 9'h000; 
        10'b0110000110: data <= 9'h000; 
        10'b0110000111: data <= 9'h000; 
        10'b0110001000: data <= 9'h000; 
        10'b0110001001: data <= 9'h000; 
        10'b0110001010: data <= 9'h000; 
        10'b0110001011: data <= 9'h000; 
        10'b0110001100: data <= 9'h001; 
        10'b0110001101: data <= 9'h001; 
        10'b0110001110: data <= 9'h001; 
        10'b0110001111: data <= 9'h001; 
        10'b0110010000: data <= 9'h001; 
        10'b0110010001: data <= 9'h000; 
        10'b0110010010: data <= 9'h000; 
        10'b0110010011: data <= 9'h000; 
        10'b0110010100: data <= 9'h1ff; 
        10'b0110010101: data <= 9'h001; 
        10'b0110010110: data <= 9'h000; 
        10'b0110010111: data <= 9'h002; 
        10'b0110011000: data <= 9'h002; 
        10'b0110011001: data <= 9'h002; 
        10'b0110011010: data <= 9'h001; 
        10'b0110011011: data <= 9'h001; 
        10'b0110011100: data <= 9'h001; 
        10'b0110011101: data <= 9'h000; 
        10'b0110011110: data <= 9'h1ff; 
        10'b0110011111: data <= 9'h1ff; 
        10'b0110100000: data <= 9'h1ff; 
        10'b0110100001: data <= 9'h000; 
        10'b0110100010: data <= 9'h000; 
        10'b0110100011: data <= 9'h000; 
        10'b0110100100: data <= 9'h000; 
        10'b0110100101: data <= 9'h000; 
        10'b0110100110: data <= 9'h000; 
        10'b0110100111: data <= 9'h000; 
        10'b0110101000: data <= 9'h000; 
        10'b0110101001: data <= 9'h001; 
        10'b0110101010: data <= 9'h001; 
        10'b0110101011: data <= 9'h000; 
        10'b0110101100: data <= 9'h000; 
        10'b0110101101: data <= 9'h1ff; 
        10'b0110101110: data <= 9'h000; 
        10'b0110101111: data <= 9'h000; 
        10'b0110110000: data <= 9'h1ff; 
        10'b0110110001: data <= 9'h000; 
        10'b0110110010: data <= 9'h1ff; 
        10'b0110110011: data <= 9'h002; 
        10'b0110110100: data <= 9'h003; 
        10'b0110110101: data <= 9'h003; 
        10'b0110110110: data <= 9'h001; 
        10'b0110110111: data <= 9'h000; 
        10'b0110111000: data <= 9'h1ff; 
        10'b0110111001: data <= 9'h1fe; 
        10'b0110111010: data <= 9'h1fe; 
        10'b0110111011: data <= 9'h1ff; 
        10'b0110111100: data <= 9'h1ff; 
        10'b0110111101: data <= 9'h000; 
        10'b0110111110: data <= 9'h000; 
        10'b0110111111: data <= 9'h000; 
        10'b0111000000: data <= 9'h000; 
        10'b0111000001: data <= 9'h000; 
        10'b0111000010: data <= 9'h000; 
        10'b0111000011: data <= 9'h000; 
        10'b0111000100: data <= 9'h000; 
        10'b0111000101: data <= 9'h000; 
        10'b0111000110: data <= 9'h1ff; 
        10'b0111000111: data <= 9'h000; 
        10'b0111001000: data <= 9'h001; 
        10'b0111001001: data <= 9'h000; 
        10'b0111001010: data <= 9'h001; 
        10'b0111001011: data <= 9'h001; 
        10'b0111001100: data <= 9'h000; 
        10'b0111001101: data <= 9'h1ff; 
        10'b0111001110: data <= 9'h000; 
        10'b0111001111: data <= 9'h001; 
        10'b0111010000: data <= 9'h002; 
        10'b0111010001: data <= 9'h002; 
        10'b0111010010: data <= 9'h000; 
        10'b0111010011: data <= 9'h1ff; 
        10'b0111010100: data <= 9'h1fe; 
        10'b0111010101: data <= 9'h1fe; 
        10'b0111010110: data <= 9'h1fe; 
        10'b0111010111: data <= 9'h1ff; 
        10'b0111011000: data <= 9'h1ff; 
        10'b0111011001: data <= 9'h000; 
        10'b0111011010: data <= 9'h000; 
        10'b0111011011: data <= 9'h000; 
        10'b0111011100: data <= 9'h000; 
        10'b0111011101: data <= 9'h000; 
        10'b0111011110: data <= 9'h000; 
        10'b0111011111: data <= 9'h000; 
        10'b0111100000: data <= 9'h1ff; 
        10'b0111100001: data <= 9'h1ff; 
        10'b0111100010: data <= 9'h1ff; 
        10'b0111100011: data <= 9'h000; 
        10'b0111100100: data <= 9'h001; 
        10'b0111100101: data <= 9'h001; 
        10'b0111100110: data <= 9'h001; 
        10'b0111100111: data <= 9'h002; 
        10'b0111101000: data <= 9'h001; 
        10'b0111101001: data <= 9'h000; 
        10'b0111101010: data <= 9'h001; 
        10'b0111101011: data <= 9'h002; 
        10'b0111101100: data <= 9'h000; 
        10'b0111101101: data <= 9'h000; 
        10'b0111101110: data <= 9'h1ff; 
        10'b0111101111: data <= 9'h1fe; 
        10'b0111110000: data <= 9'h1fe; 
        10'b0111110001: data <= 9'h1fe; 
        10'b0111110010: data <= 9'h1fe; 
        10'b0111110011: data <= 9'h1ff; 
        10'b0111110100: data <= 9'h1ff; 
        10'b0111110101: data <= 9'h000; 
        10'b0111110110: data <= 9'h000; 
        10'b0111110111: data <= 9'h000; 
        10'b0111111000: data <= 9'h000; 
        10'b0111111001: data <= 9'h000; 
        10'b0111111010: data <= 9'h000; 
        10'b0111111011: data <= 9'h000; 
        10'b0111111100: data <= 9'h1ff; 
        10'b0111111101: data <= 9'h1ff; 
        10'b0111111110: data <= 9'h1ff; 
        10'b0111111111: data <= 9'h1ff; 
        10'b1000000000: data <= 9'h1ff; 
        10'b1000000001: data <= 9'h000; 
        10'b1000000010: data <= 9'h002; 
        10'b1000000011: data <= 9'h001; 
        10'b1000000100: data <= 9'h1ff; 
        10'b1000000101: data <= 9'h1ff; 
        10'b1000000110: data <= 9'h000; 
        10'b1000000111: data <= 9'h001; 
        10'b1000001000: data <= 9'h1ff; 
        10'b1000001001: data <= 9'h1ff; 
        10'b1000001010: data <= 9'h1ff; 
        10'b1000001011: data <= 9'h1ff; 
        10'b1000001100: data <= 9'h1ff; 
        10'b1000001101: data <= 9'h1ff; 
        10'b1000001110: data <= 9'h1ff; 
        10'b1000001111: data <= 9'h1ff; 
        10'b1000010000: data <= 9'h1ff; 
        10'b1000010001: data <= 9'h000; 
        10'b1000010010: data <= 9'h000; 
        10'b1000010011: data <= 9'h000; 
        10'b1000010100: data <= 9'h000; 
        10'b1000010101: data <= 9'h000; 
        10'b1000010110: data <= 9'h000; 
        10'b1000010111: data <= 9'h000; 
        10'b1000011000: data <= 9'h1ff; 
        10'b1000011001: data <= 9'h1ff; 
        10'b1000011010: data <= 9'h1fe; 
        10'b1000011011: data <= 9'h1fe; 
        10'b1000011100: data <= 9'h1fe; 
        10'b1000011101: data <= 9'h1fe; 
        10'b1000011110: data <= 9'h1fe; 
        10'b1000011111: data <= 9'h1fe; 
        10'b1000100000: data <= 9'h1fe; 
        10'b1000100001: data <= 9'h1ff; 
        10'b1000100010: data <= 9'h1ff; 
        10'b1000100011: data <= 9'h1ff; 
        10'b1000100100: data <= 9'h1ff; 
        10'b1000100101: data <= 9'h000; 
        10'b1000100110: data <= 9'h1ff; 
        10'b1000100111: data <= 9'h000; 
        10'b1000101000: data <= 9'h1ff; 
        10'b1000101001: data <= 9'h1ff; 
        10'b1000101010: data <= 9'h1ff; 
        10'b1000101011: data <= 9'h1ff; 
        10'b1000101100: data <= 9'h000; 
        10'b1000101101: data <= 9'h000; 
        10'b1000101110: data <= 9'h000; 
        10'b1000101111: data <= 9'h000; 
        10'b1000110000: data <= 9'h000; 
        10'b1000110001: data <= 9'h000; 
        10'b1000110010: data <= 9'h000; 
        10'b1000110011: data <= 9'h000; 
        10'b1000110100: data <= 9'h1ff; 
        10'b1000110101: data <= 9'h1ff; 
        10'b1000110110: data <= 9'h1ff; 
        10'b1000110111: data <= 9'h1fe; 
        10'b1000111000: data <= 9'h1fd; 
        10'b1000111001: data <= 9'h1fd; 
        10'b1000111010: data <= 9'h1fc; 
        10'b1000111011: data <= 9'h1fd; 
        10'b1000111100: data <= 9'h1fd; 
        10'b1000111101: data <= 9'h1ff; 
        10'b1000111110: data <= 9'h1ff; 
        10'b1000111111: data <= 9'h1ff; 
        10'b1001000000: data <= 9'h1ff; 
        10'b1001000001: data <= 9'h000; 
        10'b1001000010: data <= 9'h1ff; 
        10'b1001000011: data <= 9'h000; 
        10'b1001000100: data <= 9'h1ff; 
        10'b1001000101: data <= 9'h1ff; 
        10'b1001000110: data <= 9'h000; 
        10'b1001000111: data <= 9'h000; 
        10'b1001001000: data <= 9'h000; 
        10'b1001001001: data <= 9'h000; 
        10'b1001001010: data <= 9'h000; 
        10'b1001001011: data <= 9'h000; 
        10'b1001001100: data <= 9'h000; 
        10'b1001001101: data <= 9'h000; 
        10'b1001001110: data <= 9'h000; 
        10'b1001001111: data <= 9'h000; 
        10'b1001010000: data <= 9'h000; 
        10'b1001010001: data <= 9'h1ff; 
        10'b1001010010: data <= 9'h1ff; 
        10'b1001010011: data <= 9'h1fe; 
        10'b1001010100: data <= 9'h1fe; 
        10'b1001010101: data <= 9'h1fd; 
        10'b1001010110: data <= 9'h1fd; 
        10'b1001010111: data <= 9'h1fe; 
        10'b1001011000: data <= 9'h1fe; 
        10'b1001011001: data <= 9'h1fe; 
        10'b1001011010: data <= 9'h1fe; 
        10'b1001011011: data <= 9'h1ff; 
        10'b1001011100: data <= 9'h1ff; 
        10'b1001011101: data <= 9'h1ff; 
        10'b1001011110: data <= 9'h1fe; 
        10'b1001011111: data <= 9'h1ff; 
        10'b1001100000: data <= 9'h000; 
        10'b1001100001: data <= 9'h000; 
        10'b1001100010: data <= 9'h000; 
        10'b1001100011: data <= 9'h000; 
        10'b1001100100: data <= 9'h000; 
        10'b1001100101: data <= 9'h000; 
        10'b1001100110: data <= 9'h000; 
        10'b1001100111: data <= 9'h000; 
        10'b1001101000: data <= 9'h000; 
        10'b1001101001: data <= 9'h000; 
        10'b1001101010: data <= 9'h000; 
        10'b1001101011: data <= 9'h000; 
        10'b1001101100: data <= 9'h000; 
        10'b1001101101: data <= 9'h1ff; 
        10'b1001101110: data <= 9'h1ff; 
        10'b1001101111: data <= 9'h1fe; 
        10'b1001110000: data <= 9'h1ff; 
        10'b1001110001: data <= 9'h1ff; 
        10'b1001110010: data <= 9'h1ff; 
        10'b1001110011: data <= 9'h1ff; 
        10'b1001110100: data <= 9'h1ff; 
        10'b1001110101: data <= 9'h1ff; 
        10'b1001110110: data <= 9'h1ff; 
        10'b1001110111: data <= 9'h1fe; 
        10'b1001111000: data <= 9'h1fe; 
        10'b1001111001: data <= 9'h1fe; 
        10'b1001111010: data <= 9'h1fe; 
        10'b1001111011: data <= 9'h1ff; 
        10'b1001111100: data <= 9'h000; 
        10'b1001111101: data <= 9'h000; 
        10'b1001111110: data <= 9'h000; 
        10'b1001111111: data <= 9'h000; 
        10'b1010000000: data <= 9'h001; 
        10'b1010000001: data <= 9'h000; 
        10'b1010000010: data <= 9'h000; 
        10'b1010000011: data <= 9'h000; 
        10'b1010000100: data <= 9'h000; 
        10'b1010000101: data <= 9'h000; 
        10'b1010000110: data <= 9'h000; 
        10'b1010000111: data <= 9'h000; 
        10'b1010001000: data <= 9'h000; 
        10'b1010001001: data <= 9'h1ff; 
        10'b1010001010: data <= 9'h1ff; 
        10'b1010001011: data <= 9'h1ff; 
        10'b1010001100: data <= 9'h000; 
        10'b1010001101: data <= 9'h000; 
        10'b1010001110: data <= 9'h000; 
        10'b1010001111: data <= 9'h1ff; 
        10'b1010010000: data <= 9'h1ff; 
        10'b1010010001: data <= 9'h1ff; 
        10'b1010010010: data <= 9'h1ff; 
        10'b1010010011: data <= 9'h1fe; 
        10'b1010010100: data <= 9'h1fe; 
        10'b1010010101: data <= 9'h1fe; 
        10'b1010010110: data <= 9'h1ff; 
        10'b1010010111: data <= 9'h000; 
        10'b1010011000: data <= 9'h000; 
        10'b1010011001: data <= 9'h001; 
        10'b1010011010: data <= 9'h001; 
        10'b1010011011: data <= 9'h001; 
        10'b1010011100: data <= 9'h001; 
        10'b1010011101: data <= 9'h000; 
        10'b1010011110: data <= 9'h000; 
        10'b1010011111: data <= 9'h000; 
        10'b1010100000: data <= 9'h000; 
        10'b1010100001: data <= 9'h000; 
        10'b1010100010: data <= 9'h000; 
        10'b1010100011: data <= 9'h000; 
        10'b1010100100: data <= 9'h000; 
        10'b1010100101: data <= 9'h000; 
        10'b1010100110: data <= 9'h000; 
        10'b1010100111: data <= 9'h000; 
        10'b1010101000: data <= 9'h001; 
        10'b1010101001: data <= 9'h000; 
        10'b1010101010: data <= 9'h000; 
        10'b1010101011: data <= 9'h1ff; 
        10'b1010101100: data <= 9'h000; 
        10'b1010101101: data <= 9'h1ff; 
        10'b1010101110: data <= 9'h1ff; 
        10'b1010101111: data <= 9'h1ff; 
        10'b1010110000: data <= 9'h1ff; 
        10'b1010110001: data <= 9'h000; 
        10'b1010110010: data <= 9'h001; 
        10'b1010110011: data <= 9'h001; 
        10'b1010110100: data <= 9'h002; 
        10'b1010110101: data <= 9'h002; 
        10'b1010110110: data <= 9'h001; 
        10'b1010110111: data <= 9'h001; 
        10'b1010111000: data <= 9'h001; 
        10'b1010111001: data <= 9'h000; 
        10'b1010111010: data <= 9'h000; 
        10'b1010111011: data <= 9'h000; 
        10'b1010111100: data <= 9'h000; 
        10'b1010111101: data <= 9'h000; 
        10'b1010111110: data <= 9'h000; 
        10'b1010111111: data <= 9'h000; 
        10'b1011000000: data <= 9'h000; 
        10'b1011000001: data <= 9'h001; 
        10'b1011000010: data <= 9'h000; 
        10'b1011000011: data <= 9'h001; 
        10'b1011000100: data <= 9'h001; 
        10'b1011000101: data <= 9'h001; 
        10'b1011000110: data <= 9'h001; 
        10'b1011000111: data <= 9'h000; 
        10'b1011001000: data <= 9'h001; 
        10'b1011001001: data <= 9'h001; 
        10'b1011001010: data <= 9'h001; 
        10'b1011001011: data <= 9'h001; 
        10'b1011001100: data <= 9'h002; 
        10'b1011001101: data <= 9'h002; 
        10'b1011001110: data <= 9'h002; 
        10'b1011001111: data <= 9'h002; 
        10'b1011010000: data <= 9'h003; 
        10'b1011010001: data <= 9'h002; 
        10'b1011010010: data <= 9'h001; 
        10'b1011010011: data <= 9'h000; 
        10'b1011010100: data <= 9'h000; 
        10'b1011010101: data <= 9'h000; 
        10'b1011010110: data <= 9'h000; 
        10'b1011010111: data <= 9'h000; 
        10'b1011011000: data <= 9'h000; 
        10'b1011011001: data <= 9'h000; 
        10'b1011011010: data <= 9'h000; 
        10'b1011011011: data <= 9'h000; 
        10'b1011011100: data <= 9'h000; 
        10'b1011011101: data <= 9'h000; 
        10'b1011011110: data <= 9'h001; 
        10'b1011011111: data <= 9'h001; 
        10'b1011100000: data <= 9'h001; 
        10'b1011100001: data <= 9'h002; 
        10'b1011100010: data <= 9'h002; 
        10'b1011100011: data <= 9'h002; 
        10'b1011100100: data <= 9'h002; 
        10'b1011100101: data <= 9'h002; 
        10'b1011100110: data <= 9'h003; 
        10'b1011100111: data <= 9'h002; 
        10'b1011101000: data <= 9'h001; 
        10'b1011101001: data <= 9'h001; 
        10'b1011101010: data <= 9'h001; 
        10'b1011101011: data <= 9'h001; 
        10'b1011101100: data <= 9'h001; 
        10'b1011101101: data <= 9'h001; 
        10'b1011101110: data <= 9'h000; 
        10'b1011101111: data <= 9'h000; 
        10'b1011110000: data <= 9'h000; 
        10'b1011110001: data <= 9'h000; 
        10'b1011110010: data <= 9'h000; 
        10'b1011110011: data <= 9'h000; 
        10'b1011110100: data <= 9'h000; 
        10'b1011110101: data <= 9'h000; 
        10'b1011110110: data <= 9'h000; 
        10'b1011110111: data <= 9'h000; 
        10'b1011111000: data <= 9'h000; 
        10'b1011111001: data <= 9'h000; 
        10'b1011111010: data <= 9'h000; 
        10'b1011111011: data <= 9'h000; 
        10'b1011111100: data <= 9'h000; 
        10'b1011111101: data <= 9'h000; 
        10'b1011111110: data <= 9'h000; 
        10'b1011111111: data <= 9'h000; 
        10'b1100000000: data <= 9'h000; 
        10'b1100000001: data <= 9'h000; 
        10'b1100000010: data <= 9'h000; 
        10'b1100000011: data <= 9'h000; 
        10'b1100000100: data <= 9'h000; 
        10'b1100000101: data <= 9'h000; 
        10'b1100000110: data <= 9'h000; 
        10'b1100000111: data <= 9'h000; 
        10'b1100001000: data <= 9'h000; 
        10'b1100001001: data <= 9'h000; 
        10'b1100001010: data <= 9'h000; 
        10'b1100001011: data <= 9'h000; 
        10'b1100001100: data <= 9'h000; 
        10'b1100001101: data <= 9'h000; 
        10'b1100001110: data <= 9'h000; 
        10'b1100001111: data <= 9'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 4) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 10'h001; 
        10'b0000000001: data <= 10'h000; 
        10'b0000000010: data <= 10'h000; 
        10'b0000000011: data <= 10'h000; 
        10'b0000000100: data <= 10'h000; 
        10'b0000000101: data <= 10'h001; 
        10'b0000000110: data <= 10'h000; 
        10'b0000000111: data <= 10'h000; 
        10'b0000001000: data <= 10'h001; 
        10'b0000001001: data <= 10'h000; 
        10'b0000001010: data <= 10'h000; 
        10'b0000001011: data <= 10'h000; 
        10'b0000001100: data <= 10'h001; 
        10'b0000001101: data <= 10'h000; 
        10'b0000001110: data <= 10'h000; 
        10'b0000001111: data <= 10'h000; 
        10'b0000010000: data <= 10'h000; 
        10'b0000010001: data <= 10'h000; 
        10'b0000010010: data <= 10'h001; 
        10'b0000010011: data <= 10'h000; 
        10'b0000010100: data <= 10'h000; 
        10'b0000010101: data <= 10'h000; 
        10'b0000010110: data <= 10'h000; 
        10'b0000010111: data <= 10'h000; 
        10'b0000011000: data <= 10'h001; 
        10'b0000011001: data <= 10'h000; 
        10'b0000011010: data <= 10'h000; 
        10'b0000011011: data <= 10'h000; 
        10'b0000011100: data <= 10'h001; 
        10'b0000011101: data <= 10'h000; 
        10'b0000011110: data <= 10'h000; 
        10'b0000011111: data <= 10'h000; 
        10'b0000100000: data <= 10'h000; 
        10'b0000100001: data <= 10'h000; 
        10'b0000100010: data <= 10'h000; 
        10'b0000100011: data <= 10'h001; 
        10'b0000100100: data <= 10'h000; 
        10'b0000100101: data <= 10'h001; 
        10'b0000100110: data <= 10'h000; 
        10'b0000100111: data <= 10'h000; 
        10'b0000101000: data <= 10'h000; 
        10'b0000101001: data <= 10'h000; 
        10'b0000101010: data <= 10'h000; 
        10'b0000101011: data <= 10'h000; 
        10'b0000101100: data <= 10'h000; 
        10'b0000101101: data <= 10'h000; 
        10'b0000101110: data <= 10'h000; 
        10'b0000101111: data <= 10'h000; 
        10'b0000110000: data <= 10'h001; 
        10'b0000110001: data <= 10'h000; 
        10'b0000110010: data <= 10'h000; 
        10'b0000110011: data <= 10'h000; 
        10'b0000110100: data <= 10'h000; 
        10'b0000110101: data <= 10'h001; 
        10'b0000110110: data <= 10'h000; 
        10'b0000110111: data <= 10'h000; 
        10'b0000111000: data <= 10'h001; 
        10'b0000111001: data <= 10'h001; 
        10'b0000111010: data <= 10'h000; 
        10'b0000111011: data <= 10'h000; 
        10'b0000111100: data <= 10'h001; 
        10'b0000111101: data <= 10'h000; 
        10'b0000111110: data <= 10'h000; 
        10'b0000111111: data <= 10'h000; 
        10'b0001000000: data <= 10'h001; 
        10'b0001000001: data <= 10'h000; 
        10'b0001000010: data <= 10'h000; 
        10'b0001000011: data <= 10'h000; 
        10'b0001000100: data <= 10'h000; 
        10'b0001000101: data <= 10'h001; 
        10'b0001000110: data <= 10'h000; 
        10'b0001000111: data <= 10'h001; 
        10'b0001001000: data <= 10'h000; 
        10'b0001001001: data <= 10'h000; 
        10'b0001001010: data <= 10'h000; 
        10'b0001001011: data <= 10'h000; 
        10'b0001001100: data <= 10'h001; 
        10'b0001001101: data <= 10'h000; 
        10'b0001001110: data <= 10'h000; 
        10'b0001001111: data <= 10'h001; 
        10'b0001010000: data <= 10'h000; 
        10'b0001010001: data <= 10'h000; 
        10'b0001010010: data <= 10'h000; 
        10'b0001010011: data <= 10'h000; 
        10'b0001010100: data <= 10'h001; 
        10'b0001010101: data <= 10'h000; 
        10'b0001010110: data <= 10'h000; 
        10'b0001010111: data <= 10'h000; 
        10'b0001011000: data <= 10'h000; 
        10'b0001011001: data <= 10'h000; 
        10'b0001011010: data <= 10'h001; 
        10'b0001011011: data <= 10'h000; 
        10'b0001011100: data <= 10'h000; 
        10'b0001011101: data <= 10'h001; 
        10'b0001011110: data <= 10'h000; 
        10'b0001011111: data <= 10'h001; 
        10'b0001100000: data <= 10'h000; 
        10'b0001100001: data <= 10'h3ff; 
        10'b0001100010: data <= 10'h000; 
        10'b0001100011: data <= 10'h3ff; 
        10'b0001100100: data <= 10'h000; 
        10'b0001100101: data <= 10'h000; 
        10'b0001100110: data <= 10'h000; 
        10'b0001100111: data <= 10'h000; 
        10'b0001101000: data <= 10'h000; 
        10'b0001101001: data <= 10'h000; 
        10'b0001101010: data <= 10'h001; 
        10'b0001101011: data <= 10'h000; 
        10'b0001101100: data <= 10'h000; 
        10'b0001101101: data <= 10'h001; 
        10'b0001101110: data <= 10'h000; 
        10'b0001101111: data <= 10'h000; 
        10'b0001110000: data <= 10'h000; 
        10'b0001110001: data <= 10'h000; 
        10'b0001110010: data <= 10'h000; 
        10'b0001110011: data <= 10'h000; 
        10'b0001110100: data <= 10'h000; 
        10'b0001110101: data <= 10'h000; 
        10'b0001110110: data <= 10'h000; 
        10'b0001110111: data <= 10'h000; 
        10'b0001111000: data <= 10'h000; 
        10'b0001111001: data <= 10'h000; 
        10'b0001111010: data <= 10'h3ff; 
        10'b0001111011: data <= 10'h3ff; 
        10'b0001111100: data <= 10'h3ff; 
        10'b0001111101: data <= 10'h3fe; 
        10'b0001111110: data <= 10'h3fd; 
        10'b0001111111: data <= 10'h3fc; 
        10'b0010000000: data <= 10'h3fd; 
        10'b0010000001: data <= 10'h3fd; 
        10'b0010000010: data <= 10'h3fe; 
        10'b0010000011: data <= 10'h3ff; 
        10'b0010000100: data <= 10'h000; 
        10'b0010000101: data <= 10'h000; 
        10'b0010000110: data <= 10'h000; 
        10'b0010000111: data <= 10'h001; 
        10'b0010001000: data <= 10'h000; 
        10'b0010001001: data <= 10'h000; 
        10'b0010001010: data <= 10'h000; 
        10'b0010001011: data <= 10'h000; 
        10'b0010001100: data <= 10'h001; 
        10'b0010001101: data <= 10'h000; 
        10'b0010001110: data <= 10'h000; 
        10'b0010001111: data <= 10'h000; 
        10'b0010010000: data <= 10'h000; 
        10'b0010010001: data <= 10'h000; 
        10'b0010010010: data <= 10'h000; 
        10'b0010010011: data <= 10'h000; 
        10'b0010010100: data <= 10'h3ff; 
        10'b0010010101: data <= 10'h3ff; 
        10'b0010010110: data <= 10'h3fe; 
        10'b0010010111: data <= 10'h3fe; 
        10'b0010011000: data <= 10'h3fe; 
        10'b0010011001: data <= 10'h3fd; 
        10'b0010011010: data <= 10'h3fc; 
        10'b0010011011: data <= 10'h3fb; 
        10'b0010011100: data <= 10'h3fa; 
        10'b0010011101: data <= 10'h3fc; 
        10'b0010011110: data <= 10'h3fd; 
        10'b0010011111: data <= 10'h3ff; 
        10'b0010100000: data <= 10'h3ff; 
        10'b0010100001: data <= 10'h3fe; 
        10'b0010100010: data <= 10'h3fe; 
        10'b0010100011: data <= 10'h3ff; 
        10'b0010100100: data <= 10'h000; 
        10'b0010100101: data <= 10'h000; 
        10'b0010100110: data <= 10'h000; 
        10'b0010100111: data <= 10'h000; 
        10'b0010101000: data <= 10'h001; 
        10'b0010101001: data <= 10'h001; 
        10'b0010101010: data <= 10'h000; 
        10'b0010101011: data <= 10'h001; 
        10'b0010101100: data <= 10'h000; 
        10'b0010101101: data <= 10'h3fe; 
        10'b0010101110: data <= 10'h3fe; 
        10'b0010101111: data <= 10'h3fe; 
        10'b0010110000: data <= 10'h3fe; 
        10'b0010110001: data <= 10'h3fd; 
        10'b0010110010: data <= 10'h3fe; 
        10'b0010110011: data <= 10'h3ff; 
        10'b0010110100: data <= 10'h000; 
        10'b0010110101: data <= 10'h003; 
        10'b0010110110: data <= 10'h004; 
        10'b0010110111: data <= 10'h003; 
        10'b0010111000: data <= 10'h002; 
        10'b0010111001: data <= 10'h002; 
        10'b0010111010: data <= 10'h002; 
        10'b0010111011: data <= 10'h000; 
        10'b0010111100: data <= 10'h3ff; 
        10'b0010111101: data <= 10'h3fe; 
        10'b0010111110: data <= 10'h3fd; 
        10'b0010111111: data <= 10'h3fd; 
        10'b0011000000: data <= 10'h3fe; 
        10'b0011000001: data <= 10'h3ff; 
        10'b0011000010: data <= 10'h000; 
        10'b0011000011: data <= 10'h000; 
        10'b0011000100: data <= 10'h001; 
        10'b0011000101: data <= 10'h000; 
        10'b0011000110: data <= 10'h000; 
        10'b0011000111: data <= 10'h000; 
        10'b0011001000: data <= 10'h3fe; 
        10'b0011001001: data <= 10'h3fd; 
        10'b0011001010: data <= 10'h3fd; 
        10'b0011001011: data <= 10'h3fc; 
        10'b0011001100: data <= 10'h3fd; 
        10'b0011001101: data <= 10'h3ff; 
        10'b0011001110: data <= 10'h000; 
        10'b0011001111: data <= 10'h001; 
        10'b0011010000: data <= 10'h004; 
        10'b0011010001: data <= 10'h004; 
        10'b0011010010: data <= 10'h006; 
        10'b0011010011: data <= 10'h006; 
        10'b0011010100: data <= 10'h006; 
        10'b0011010101: data <= 10'h003; 
        10'b0011010110: data <= 10'h002; 
        10'b0011010111: data <= 10'h000; 
        10'b0011011000: data <= 10'h001; 
        10'b0011011001: data <= 10'h001; 
        10'b0011011010: data <= 10'h3fe; 
        10'b0011011011: data <= 10'h3fc; 
        10'b0011011100: data <= 10'h3fe; 
        10'b0011011101: data <= 10'h3ff; 
        10'b0011011110: data <= 10'h3ff; 
        10'b0011011111: data <= 10'h001; 
        10'b0011100000: data <= 10'h001; 
        10'b0011100001: data <= 10'h001; 
        10'b0011100010: data <= 10'h000; 
        10'b0011100011: data <= 10'h000; 
        10'b0011100100: data <= 10'h3fe; 
        10'b0011100101: data <= 10'h3fd; 
        10'b0011100110: data <= 10'h3fd; 
        10'b0011100111: data <= 10'h3fc; 
        10'b0011101000: data <= 10'h3ff; 
        10'b0011101001: data <= 10'h3ff; 
        10'b0011101010: data <= 10'h3ff; 
        10'b0011101011: data <= 10'h3ff; 
        10'b0011101100: data <= 10'h000; 
        10'b0011101101: data <= 10'h002; 
        10'b0011101110: data <= 10'h005; 
        10'b0011101111: data <= 10'h003; 
        10'b0011110000: data <= 10'h003; 
        10'b0011110001: data <= 10'h001; 
        10'b0011110010: data <= 10'h000; 
        10'b0011110011: data <= 10'h000; 
        10'b0011110100: data <= 10'h3ff; 
        10'b0011110101: data <= 10'h000; 
        10'b0011110110: data <= 10'h3ff; 
        10'b0011110111: data <= 10'h3fd; 
        10'b0011111000: data <= 10'h3fd; 
        10'b0011111001: data <= 10'h3ff; 
        10'b0011111010: data <= 10'h3ff; 
        10'b0011111011: data <= 10'h001; 
        10'b0011111100: data <= 10'h000; 
        10'b0011111101: data <= 10'h000; 
        10'b0011111110: data <= 10'h000; 
        10'b0011111111: data <= 10'h3ff; 
        10'b0100000000: data <= 10'h3fd; 
        10'b0100000001: data <= 10'h3fe; 
        10'b0100000010: data <= 10'h3ff; 
        10'b0100000011: data <= 10'h3ff; 
        10'b0100000100: data <= 10'h3ff; 
        10'b0100000101: data <= 10'h000; 
        10'b0100000110: data <= 10'h001; 
        10'b0100000111: data <= 10'h001; 
        10'b0100001000: data <= 10'h000; 
        10'b0100001001: data <= 10'h002; 
        10'b0100001010: data <= 10'h004; 
        10'b0100001011: data <= 10'h003; 
        10'b0100001100: data <= 10'h000; 
        10'b0100001101: data <= 10'h3ff; 
        10'b0100001110: data <= 10'h000; 
        10'b0100001111: data <= 10'h3fe; 
        10'b0100010000: data <= 10'h3ff; 
        10'b0100010001: data <= 10'h3fe; 
        10'b0100010010: data <= 10'h3fe; 
        10'b0100010011: data <= 10'h3fe; 
        10'b0100010100: data <= 10'h3fe; 
        10'b0100010101: data <= 10'h3ff; 
        10'b0100010110: data <= 10'h000; 
        10'b0100010111: data <= 10'h001; 
        10'b0100011000: data <= 10'h000; 
        10'b0100011001: data <= 10'h000; 
        10'b0100011010: data <= 10'h000; 
        10'b0100011011: data <= 10'h000; 
        10'b0100011100: data <= 10'h3fe; 
        10'b0100011101: data <= 10'h3ff; 
        10'b0100011110: data <= 10'h001; 
        10'b0100011111: data <= 10'h001; 
        10'b0100100000: data <= 10'h003; 
        10'b0100100001: data <= 10'h003; 
        10'b0100100010: data <= 10'h002; 
        10'b0100100011: data <= 10'h004; 
        10'b0100100100: data <= 10'h002; 
        10'b0100100101: data <= 10'h000; 
        10'b0100100110: data <= 10'h000; 
        10'b0100100111: data <= 10'h3fe; 
        10'b0100101000: data <= 10'h3ff; 
        10'b0100101001: data <= 10'h000; 
        10'b0100101010: data <= 10'h001; 
        10'b0100101011: data <= 10'h000; 
        10'b0100101100: data <= 10'h001; 
        10'b0100101101: data <= 10'h3ff; 
        10'b0100101110: data <= 10'h3ff; 
        10'b0100101111: data <= 10'h3ff; 
        10'b0100110000: data <= 10'h3fe; 
        10'b0100110001: data <= 10'h000; 
        10'b0100110010: data <= 10'h3ff; 
        10'b0100110011: data <= 10'h000; 
        10'b0100110100: data <= 10'h000; 
        10'b0100110101: data <= 10'h000; 
        10'b0100110110: data <= 10'h000; 
        10'b0100110111: data <= 10'h000; 
        10'b0100111000: data <= 10'h3ff; 
        10'b0100111001: data <= 10'h002; 
        10'b0100111010: data <= 10'h005; 
        10'b0100111011: data <= 10'h003; 
        10'b0100111100: data <= 10'h005; 
        10'b0100111101: data <= 10'h002; 
        10'b0100111110: data <= 10'h002; 
        10'b0100111111: data <= 10'h004; 
        10'b0101000000: data <= 10'h3ff; 
        10'b0101000001: data <= 10'h3ff; 
        10'b0101000010: data <= 10'h3ff; 
        10'b0101000011: data <= 10'h000; 
        10'b0101000100: data <= 10'h001; 
        10'b0101000101: data <= 10'h005; 
        10'b0101000110: data <= 10'h002; 
        10'b0101000111: data <= 10'h002; 
        10'b0101001000: data <= 10'h004; 
        10'b0101001001: data <= 10'h003; 
        10'b0101001010: data <= 10'h002; 
        10'b0101001011: data <= 10'h000; 
        10'b0101001100: data <= 10'h000; 
        10'b0101001101: data <= 10'h3ff; 
        10'b0101001110: data <= 10'h000; 
        10'b0101001111: data <= 10'h000; 
        10'b0101010000: data <= 10'h000; 
        10'b0101010001: data <= 10'h001; 
        10'b0101010010: data <= 10'h000; 
        10'b0101010011: data <= 10'h3ff; 
        10'b0101010100: data <= 10'h002; 
        10'b0101010101: data <= 10'h004; 
        10'b0101010110: data <= 10'h005; 
        10'b0101010111: data <= 10'h003; 
        10'b0101011000: data <= 10'h004; 
        10'b0101011001: data <= 10'h005; 
        10'b0101011010: data <= 10'h003; 
        10'b0101011011: data <= 10'h000; 
        10'b0101011100: data <= 10'h3fd; 
        10'b0101011101: data <= 10'h003; 
        10'b0101011110: data <= 10'h005; 
        10'b0101011111: data <= 10'h004; 
        10'b0101100000: data <= 10'h004; 
        10'b0101100001: data <= 10'h006; 
        10'b0101100010: data <= 10'h006; 
        10'b0101100011: data <= 10'h006; 
        10'b0101100100: data <= 10'h006; 
        10'b0101100101: data <= 10'h004; 
        10'b0101100110: data <= 10'h002; 
        10'b0101100111: data <= 10'h000; 
        10'b0101101000: data <= 10'h3ff; 
        10'b0101101001: data <= 10'h000; 
        10'b0101101010: data <= 10'h000; 
        10'b0101101011: data <= 10'h000; 
        10'b0101101100: data <= 10'h001; 
        10'b0101101101: data <= 10'h000; 
        10'b0101101110: data <= 10'h3ff; 
        10'b0101101111: data <= 10'h000; 
        10'b0101110000: data <= 10'h003; 
        10'b0101110001: data <= 10'h004; 
        10'b0101110010: data <= 10'h004; 
        10'b0101110011: data <= 10'h002; 
        10'b0101110100: data <= 10'h003; 
        10'b0101110101: data <= 10'h002; 
        10'b0101110110: data <= 10'h002; 
        10'b0101110111: data <= 10'h3ff; 
        10'b0101111000: data <= 10'h3fe; 
        10'b0101111001: data <= 10'h004; 
        10'b0101111010: data <= 10'h005; 
        10'b0101111011: data <= 10'h004; 
        10'b0101111100: data <= 10'h005; 
        10'b0101111101: data <= 10'h004; 
        10'b0101111110: data <= 10'h006; 
        10'b0101111111: data <= 10'h006; 
        10'b0110000000: data <= 10'h004; 
        10'b0110000001: data <= 10'h003; 
        10'b0110000010: data <= 10'h000; 
        10'b0110000011: data <= 10'h3fe; 
        10'b0110000100: data <= 10'h3ff; 
        10'b0110000101: data <= 10'h000; 
        10'b0110000110: data <= 10'h000; 
        10'b0110000111: data <= 10'h000; 
        10'b0110001000: data <= 10'h000; 
        10'b0110001001: data <= 10'h000; 
        10'b0110001010: data <= 10'h001; 
        10'b0110001011: data <= 10'h000; 
        10'b0110001100: data <= 10'h001; 
        10'b0110001101: data <= 10'h001; 
        10'b0110001110: data <= 10'h003; 
        10'b0110001111: data <= 10'h002; 
        10'b0110010000: data <= 10'h001; 
        10'b0110010001: data <= 10'h000; 
        10'b0110010010: data <= 10'h000; 
        10'b0110010011: data <= 10'h000; 
        10'b0110010100: data <= 10'h3ff; 
        10'b0110010101: data <= 10'h001; 
        10'b0110010110: data <= 10'h001; 
        10'b0110010111: data <= 10'h003; 
        10'b0110011000: data <= 10'h004; 
        10'b0110011001: data <= 10'h004; 
        10'b0110011010: data <= 10'h003; 
        10'b0110011011: data <= 10'h002; 
        10'b0110011100: data <= 10'h002; 
        10'b0110011101: data <= 10'h000; 
        10'b0110011110: data <= 10'h3fe; 
        10'b0110011111: data <= 10'h3fd; 
        10'b0110100000: data <= 10'h3ff; 
        10'b0110100001: data <= 10'h000; 
        10'b0110100010: data <= 10'h000; 
        10'b0110100011: data <= 10'h000; 
        10'b0110100100: data <= 10'h001; 
        10'b0110100101: data <= 10'h001; 
        10'b0110100110: data <= 10'h000; 
        10'b0110100111: data <= 10'h000; 
        10'b0110101000: data <= 10'h000; 
        10'b0110101001: data <= 10'h001; 
        10'b0110101010: data <= 10'h001; 
        10'b0110101011: data <= 10'h001; 
        10'b0110101100: data <= 10'h001; 
        10'b0110101101: data <= 10'h3fe; 
        10'b0110101110: data <= 10'h3ff; 
        10'b0110101111: data <= 10'h3ff; 
        10'b0110110000: data <= 10'h3ff; 
        10'b0110110001: data <= 10'h3ff; 
        10'b0110110010: data <= 10'h3ff; 
        10'b0110110011: data <= 10'h004; 
        10'b0110110100: data <= 10'h006; 
        10'b0110110101: data <= 10'h005; 
        10'b0110110110: data <= 10'h003; 
        10'b0110110111: data <= 10'h000; 
        10'b0110111000: data <= 10'h3ff; 
        10'b0110111001: data <= 10'h3fd; 
        10'b0110111010: data <= 10'h3fc; 
        10'b0110111011: data <= 10'h3fd; 
        10'b0110111100: data <= 10'h3ff; 
        10'b0110111101: data <= 10'h000; 
        10'b0110111110: data <= 10'h000; 
        10'b0110111111: data <= 10'h000; 
        10'b0111000000: data <= 10'h001; 
        10'b0111000001: data <= 10'h000; 
        10'b0111000010: data <= 10'h000; 
        10'b0111000011: data <= 10'h000; 
        10'b0111000100: data <= 10'h000; 
        10'b0111000101: data <= 10'h000; 
        10'b0111000110: data <= 10'h3ff; 
        10'b0111000111: data <= 10'h001; 
        10'b0111001000: data <= 10'h002; 
        10'b0111001001: data <= 10'h3ff; 
        10'b0111001010: data <= 10'h001; 
        10'b0111001011: data <= 10'h002; 
        10'b0111001100: data <= 10'h000; 
        10'b0111001101: data <= 10'h3fe; 
        10'b0111001110: data <= 10'h000; 
        10'b0111001111: data <= 10'h002; 
        10'b0111010000: data <= 10'h004; 
        10'b0111010001: data <= 10'h004; 
        10'b0111010010: data <= 10'h001; 
        10'b0111010011: data <= 10'h3fe; 
        10'b0111010100: data <= 10'h3fc; 
        10'b0111010101: data <= 10'h3fb; 
        10'b0111010110: data <= 10'h3fd; 
        10'b0111010111: data <= 10'h3fd; 
        10'b0111011000: data <= 10'h3fe; 
        10'b0111011001: data <= 10'h000; 
        10'b0111011010: data <= 10'h000; 
        10'b0111011011: data <= 10'h000; 
        10'b0111011100: data <= 10'h000; 
        10'b0111011101: data <= 10'h000; 
        10'b0111011110: data <= 10'h3ff; 
        10'b0111011111: data <= 10'h3ff; 
        10'b0111100000: data <= 10'h3ff; 
        10'b0111100001: data <= 10'h3fe; 
        10'b0111100010: data <= 10'h3ff; 
        10'b0111100011: data <= 10'h001; 
        10'b0111100100: data <= 10'h001; 
        10'b0111100101: data <= 10'h001; 
        10'b0111100110: data <= 10'h002; 
        10'b0111100111: data <= 10'h003; 
        10'b0111101000: data <= 10'h002; 
        10'b0111101001: data <= 10'h001; 
        10'b0111101010: data <= 10'h001; 
        10'b0111101011: data <= 10'h003; 
        10'b0111101100: data <= 10'h001; 
        10'b0111101101: data <= 10'h3ff; 
        10'b0111101110: data <= 10'h3ff; 
        10'b0111101111: data <= 10'h3fd; 
        10'b0111110000: data <= 10'h3fd; 
        10'b0111110001: data <= 10'h3fd; 
        10'b0111110010: data <= 10'h3fd; 
        10'b0111110011: data <= 10'h3fe; 
        10'b0111110100: data <= 10'h3fe; 
        10'b0111110101: data <= 10'h000; 
        10'b0111110110: data <= 10'h000; 
        10'b0111110111: data <= 10'h000; 
        10'b0111111000: data <= 10'h001; 
        10'b0111111001: data <= 10'h000; 
        10'b0111111010: data <= 10'h000; 
        10'b0111111011: data <= 10'h000; 
        10'b0111111100: data <= 10'h3ff; 
        10'b0111111101: data <= 10'h3fd; 
        10'b0111111110: data <= 10'h3fd; 
        10'b0111111111: data <= 10'h3fd; 
        10'b1000000000: data <= 10'h3ff; 
        10'b1000000001: data <= 10'h000; 
        10'b1000000010: data <= 10'h003; 
        10'b1000000011: data <= 10'h003; 
        10'b1000000100: data <= 10'h3fe; 
        10'b1000000101: data <= 10'h3fe; 
        10'b1000000110: data <= 10'h000; 
        10'b1000000111: data <= 10'h002; 
        10'b1000001000: data <= 10'h3ff; 
        10'b1000001001: data <= 10'h3ff; 
        10'b1000001010: data <= 10'h3fd; 
        10'b1000001011: data <= 10'h3fe; 
        10'b1000001100: data <= 10'h3fe; 
        10'b1000001101: data <= 10'h3fe; 
        10'b1000001110: data <= 10'h3fd; 
        10'b1000001111: data <= 10'h3fd; 
        10'b1000010000: data <= 10'h3fe; 
        10'b1000010001: data <= 10'h000; 
        10'b1000010010: data <= 10'h000; 
        10'b1000010011: data <= 10'h001; 
        10'b1000010100: data <= 10'h000; 
        10'b1000010101: data <= 10'h001; 
        10'b1000010110: data <= 10'h000; 
        10'b1000010111: data <= 10'h3ff; 
        10'b1000011000: data <= 10'h3ff; 
        10'b1000011001: data <= 10'h3fe; 
        10'b1000011010: data <= 10'h3fd; 
        10'b1000011011: data <= 10'h3fd; 
        10'b1000011100: data <= 10'h3fd; 
        10'b1000011101: data <= 10'h3fd; 
        10'b1000011110: data <= 10'h3fc; 
        10'b1000011111: data <= 10'h3fd; 
        10'b1000100000: data <= 10'h3fc; 
        10'b1000100001: data <= 10'h3fd; 
        10'b1000100010: data <= 10'h3fe; 
        10'b1000100011: data <= 10'h3fd; 
        10'b1000100100: data <= 10'h3fe; 
        10'b1000100101: data <= 10'h3ff; 
        10'b1000100110: data <= 10'h3fe; 
        10'b1000100111: data <= 10'h3ff; 
        10'b1000101000: data <= 10'h3ff; 
        10'b1000101001: data <= 10'h3ff; 
        10'b1000101010: data <= 10'h3ff; 
        10'b1000101011: data <= 10'h3ff; 
        10'b1000101100: data <= 10'h3ff; 
        10'b1000101101: data <= 10'h000; 
        10'b1000101110: data <= 10'h000; 
        10'b1000101111: data <= 10'h000; 
        10'b1000110000: data <= 10'h000; 
        10'b1000110001: data <= 10'h000; 
        10'b1000110010: data <= 10'h000; 
        10'b1000110011: data <= 10'h000; 
        10'b1000110100: data <= 10'h3ff; 
        10'b1000110101: data <= 10'h3fe; 
        10'b1000110110: data <= 10'h3fd; 
        10'b1000110111: data <= 10'h3fb; 
        10'b1000111000: data <= 10'h3fb; 
        10'b1000111001: data <= 10'h3fa; 
        10'b1000111010: data <= 10'h3f8; 
        10'b1000111011: data <= 10'h3fa; 
        10'b1000111100: data <= 10'h3fa; 
        10'b1000111101: data <= 10'h3fe; 
        10'b1000111110: data <= 10'h3fd; 
        10'b1000111111: data <= 10'h3ff; 
        10'b1001000000: data <= 10'h3fe; 
        10'b1001000001: data <= 10'h000; 
        10'b1001000010: data <= 10'h3fd; 
        10'b1001000011: data <= 10'h3ff; 
        10'b1001000100: data <= 10'h3ff; 
        10'b1001000101: data <= 10'h3fe; 
        10'b1001000110: data <= 10'h000; 
        10'b1001000111: data <= 10'h3ff; 
        10'b1001001000: data <= 10'h000; 
        10'b1001001001: data <= 10'h001; 
        10'b1001001010: data <= 10'h000; 
        10'b1001001011: data <= 10'h000; 
        10'b1001001100: data <= 10'h000; 
        10'b1001001101: data <= 10'h000; 
        10'b1001001110: data <= 10'h001; 
        10'b1001001111: data <= 10'h3ff; 
        10'b1001010000: data <= 10'h3ff; 
        10'b1001010001: data <= 10'h3fe; 
        10'b1001010010: data <= 10'h3fd; 
        10'b1001010011: data <= 10'h3fc; 
        10'b1001010100: data <= 10'h3fb; 
        10'b1001010101: data <= 10'h3fb; 
        10'b1001010110: data <= 10'h3fb; 
        10'b1001010111: data <= 10'h3fb; 
        10'b1001011000: data <= 10'h3fd; 
        10'b1001011001: data <= 10'h3fd; 
        10'b1001011010: data <= 10'h3fd; 
        10'b1001011011: data <= 10'h3fe; 
        10'b1001011100: data <= 10'h3fe; 
        10'b1001011101: data <= 10'h3fd; 
        10'b1001011110: data <= 10'h3fc; 
        10'b1001011111: data <= 10'h3fe; 
        10'b1001100000: data <= 10'h3ff; 
        10'b1001100001: data <= 10'h000; 
        10'b1001100010: data <= 10'h000; 
        10'b1001100011: data <= 10'h000; 
        10'b1001100100: data <= 10'h000; 
        10'b1001100101: data <= 10'h000; 
        10'b1001100110: data <= 10'h000; 
        10'b1001100111: data <= 10'h000; 
        10'b1001101000: data <= 10'h001; 
        10'b1001101001: data <= 10'h000; 
        10'b1001101010: data <= 10'h000; 
        10'b1001101011: data <= 10'h000; 
        10'b1001101100: data <= 10'h000; 
        10'b1001101101: data <= 10'h3fe; 
        10'b1001101110: data <= 10'h3fe; 
        10'b1001101111: data <= 10'h3fd; 
        10'b1001110000: data <= 10'h3fd; 
        10'b1001110001: data <= 10'h3fd; 
        10'b1001110010: data <= 10'h3fd; 
        10'b1001110011: data <= 10'h3fe; 
        10'b1001110100: data <= 10'h3fe; 
        10'b1001110101: data <= 10'h3fd; 
        10'b1001110110: data <= 10'h3fe; 
        10'b1001110111: data <= 10'h3fd; 
        10'b1001111000: data <= 10'h3fc; 
        10'b1001111001: data <= 10'h3fc; 
        10'b1001111010: data <= 10'h3fd; 
        10'b1001111011: data <= 10'h3fd; 
        10'b1001111100: data <= 10'h3ff; 
        10'b1001111101: data <= 10'h001; 
        10'b1001111110: data <= 10'h001; 
        10'b1001111111: data <= 10'h001; 
        10'b1010000000: data <= 10'h001; 
        10'b1010000001: data <= 10'h000; 
        10'b1010000010: data <= 10'h000; 
        10'b1010000011: data <= 10'h000; 
        10'b1010000100: data <= 10'h001; 
        10'b1010000101: data <= 10'h000; 
        10'b1010000110: data <= 10'h000; 
        10'b1010000111: data <= 10'h000; 
        10'b1010001000: data <= 10'h000; 
        10'b1010001001: data <= 10'h3ff; 
        10'b1010001010: data <= 10'h3fe; 
        10'b1010001011: data <= 10'h3fe; 
        10'b1010001100: data <= 10'h000; 
        10'b1010001101: data <= 10'h3ff; 
        10'b1010001110: data <= 10'h3ff; 
        10'b1010001111: data <= 10'h3fe; 
        10'b1010010000: data <= 10'h3fe; 
        10'b1010010001: data <= 10'h3fd; 
        10'b1010010010: data <= 10'h3fe; 
        10'b1010010011: data <= 10'h3fc; 
        10'b1010010100: data <= 10'h3fc; 
        10'b1010010101: data <= 10'h3fd; 
        10'b1010010110: data <= 10'h3fe; 
        10'b1010010111: data <= 10'h000; 
        10'b1010011000: data <= 10'h001; 
        10'b1010011001: data <= 10'h002; 
        10'b1010011010: data <= 10'h003; 
        10'b1010011011: data <= 10'h002; 
        10'b1010011100: data <= 10'h001; 
        10'b1010011101: data <= 10'h000; 
        10'b1010011110: data <= 10'h001; 
        10'b1010011111: data <= 10'h000; 
        10'b1010100000: data <= 10'h000; 
        10'b1010100001: data <= 10'h000; 
        10'b1010100010: data <= 10'h000; 
        10'b1010100011: data <= 10'h001; 
        10'b1010100100: data <= 10'h000; 
        10'b1010100101: data <= 10'h001; 
        10'b1010100110: data <= 10'h001; 
        10'b1010100111: data <= 10'h001; 
        10'b1010101000: data <= 10'h001; 
        10'b1010101001: data <= 10'h001; 
        10'b1010101010: data <= 10'h000; 
        10'b1010101011: data <= 10'h3ff; 
        10'b1010101100: data <= 10'h000; 
        10'b1010101101: data <= 10'h3fe; 
        10'b1010101110: data <= 10'h3fe; 
        10'b1010101111: data <= 10'h3fd; 
        10'b1010110000: data <= 10'h3ff; 
        10'b1010110001: data <= 10'h001; 
        10'b1010110010: data <= 10'h001; 
        10'b1010110011: data <= 10'h002; 
        10'b1010110100: data <= 10'h003; 
        10'b1010110101: data <= 10'h004; 
        10'b1010110110: data <= 10'h002; 
        10'b1010110111: data <= 10'h001; 
        10'b1010111000: data <= 10'h001; 
        10'b1010111001: data <= 10'h000; 
        10'b1010111010: data <= 10'h000; 
        10'b1010111011: data <= 10'h000; 
        10'b1010111100: data <= 10'h000; 
        10'b1010111101: data <= 10'h001; 
        10'b1010111110: data <= 10'h001; 
        10'b1010111111: data <= 10'h000; 
        10'b1011000000: data <= 10'h000; 
        10'b1011000001: data <= 10'h001; 
        10'b1011000010: data <= 10'h001; 
        10'b1011000011: data <= 10'h003; 
        10'b1011000100: data <= 10'h003; 
        10'b1011000101: data <= 10'h003; 
        10'b1011000110: data <= 10'h002; 
        10'b1011000111: data <= 10'h001; 
        10'b1011001000: data <= 10'h003; 
        10'b1011001001: data <= 10'h002; 
        10'b1011001010: data <= 10'h002; 
        10'b1011001011: data <= 10'h002; 
        10'b1011001100: data <= 10'h004; 
        10'b1011001101: data <= 10'h004; 
        10'b1011001110: data <= 10'h005; 
        10'b1011001111: data <= 10'h005; 
        10'b1011010000: data <= 10'h005; 
        10'b1011010001: data <= 10'h004; 
        10'b1011010010: data <= 10'h001; 
        10'b1011010011: data <= 10'h001; 
        10'b1011010100: data <= 10'h000; 
        10'b1011010101: data <= 10'h000; 
        10'b1011010110: data <= 10'h000; 
        10'b1011010111: data <= 10'h000; 
        10'b1011011000: data <= 10'h000; 
        10'b1011011001: data <= 10'h001; 
        10'b1011011010: data <= 10'h000; 
        10'b1011011011: data <= 10'h000; 
        10'b1011011100: data <= 10'h001; 
        10'b1011011101: data <= 10'h001; 
        10'b1011011110: data <= 10'h001; 
        10'b1011011111: data <= 10'h002; 
        10'b1011100000: data <= 10'h002; 
        10'b1011100001: data <= 10'h003; 
        10'b1011100010: data <= 10'h003; 
        10'b1011100011: data <= 10'h004; 
        10'b1011100100: data <= 10'h004; 
        10'b1011100101: data <= 10'h004; 
        10'b1011100110: data <= 10'h005; 
        10'b1011100111: data <= 10'h003; 
        10'b1011101000: data <= 10'h002; 
        10'b1011101001: data <= 10'h002; 
        10'b1011101010: data <= 10'h003; 
        10'b1011101011: data <= 10'h003; 
        10'b1011101100: data <= 10'h002; 
        10'b1011101101: data <= 10'h001; 
        10'b1011101110: data <= 10'h001; 
        10'b1011101111: data <= 10'h000; 
        10'b1011110000: data <= 10'h000; 
        10'b1011110001: data <= 10'h000; 
        10'b1011110010: data <= 10'h000; 
        10'b1011110011: data <= 10'h000; 
        10'b1011110100: data <= 10'h000; 
        10'b1011110101: data <= 10'h000; 
        10'b1011110110: data <= 10'h000; 
        10'b1011110111: data <= 10'h001; 
        10'b1011111000: data <= 10'h000; 
        10'b1011111001: data <= 10'h000; 
        10'b1011111010: data <= 10'h000; 
        10'b1011111011: data <= 10'h001; 
        10'b1011111100: data <= 10'h001; 
        10'b1011111101: data <= 10'h000; 
        10'b1011111110: data <= 10'h000; 
        10'b1011111111: data <= 10'h000; 
        10'b1100000000: data <= 10'h000; 
        10'b1100000001: data <= 10'h000; 
        10'b1100000010: data <= 10'h000; 
        10'b1100000011: data <= 10'h000; 
        10'b1100000100: data <= 10'h000; 
        10'b1100000101: data <= 10'h000; 
        10'b1100000110: data <= 10'h001; 
        10'b1100000111: data <= 10'h001; 
        10'b1100001000: data <= 10'h000; 
        10'b1100001001: data <= 10'h000; 
        10'b1100001010: data <= 10'h000; 
        10'b1100001011: data <= 10'h001; 
        10'b1100001100: data <= 10'h000; 
        10'b1100001101: data <= 10'h000; 
        10'b1100001110: data <= 10'h000; 
        10'b1100001111: data <= 10'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 5) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 11'h001; 
        10'b0000000001: data <= 11'h001; 
        10'b0000000010: data <= 11'h000; 
        10'b0000000011: data <= 11'h001; 
        10'b0000000100: data <= 11'h001; 
        10'b0000000101: data <= 11'h001; 
        10'b0000000110: data <= 11'h000; 
        10'b0000000111: data <= 11'h000; 
        10'b0000001000: data <= 11'h001; 
        10'b0000001001: data <= 11'h000; 
        10'b0000001010: data <= 11'h000; 
        10'b0000001011: data <= 11'h001; 
        10'b0000001100: data <= 11'h002; 
        10'b0000001101: data <= 11'h001; 
        10'b0000001110: data <= 11'h7ff; 
        10'b0000001111: data <= 11'h000; 
        10'b0000010000: data <= 11'h000; 
        10'b0000010001: data <= 11'h001; 
        10'b0000010010: data <= 11'h001; 
        10'b0000010011: data <= 11'h000; 
        10'b0000010100: data <= 11'h000; 
        10'b0000010101: data <= 11'h000; 
        10'b0000010110: data <= 11'h000; 
        10'b0000010111: data <= 11'h000; 
        10'b0000011000: data <= 11'h001; 
        10'b0000011001: data <= 11'h000; 
        10'b0000011010: data <= 11'h7ff; 
        10'b0000011011: data <= 11'h001; 
        10'b0000011100: data <= 11'h001; 
        10'b0000011101: data <= 11'h001; 
        10'b0000011110: data <= 11'h000; 
        10'b0000011111: data <= 11'h000; 
        10'b0000100000: data <= 11'h7ff; 
        10'b0000100001: data <= 11'h000; 
        10'b0000100010: data <= 11'h000; 
        10'b0000100011: data <= 11'h002; 
        10'b0000100100: data <= 11'h7ff; 
        10'b0000100101: data <= 11'h001; 
        10'b0000100110: data <= 11'h000; 
        10'b0000100111: data <= 11'h001; 
        10'b0000101000: data <= 11'h001; 
        10'b0000101001: data <= 11'h001; 
        10'b0000101010: data <= 11'h000; 
        10'b0000101011: data <= 11'h7ff; 
        10'b0000101100: data <= 11'h000; 
        10'b0000101101: data <= 11'h001; 
        10'b0000101110: data <= 11'h000; 
        10'b0000101111: data <= 11'h000; 
        10'b0000110000: data <= 11'h001; 
        10'b0000110001: data <= 11'h000; 
        10'b0000110010: data <= 11'h000; 
        10'b0000110011: data <= 11'h000; 
        10'b0000110100: data <= 11'h001; 
        10'b0000110101: data <= 11'h001; 
        10'b0000110110: data <= 11'h000; 
        10'b0000110111: data <= 11'h000; 
        10'b0000111000: data <= 11'h001; 
        10'b0000111001: data <= 11'h001; 
        10'b0000111010: data <= 11'h000; 
        10'b0000111011: data <= 11'h001; 
        10'b0000111100: data <= 11'h001; 
        10'b0000111101: data <= 11'h000; 
        10'b0000111110: data <= 11'h000; 
        10'b0000111111: data <= 11'h000; 
        10'b0001000000: data <= 11'h001; 
        10'b0001000001: data <= 11'h000; 
        10'b0001000010: data <= 11'h000; 
        10'b0001000011: data <= 11'h001; 
        10'b0001000100: data <= 11'h001; 
        10'b0001000101: data <= 11'h001; 
        10'b0001000110: data <= 11'h7ff; 
        10'b0001000111: data <= 11'h001; 
        10'b0001001000: data <= 11'h000; 
        10'b0001001001: data <= 11'h000; 
        10'b0001001010: data <= 11'h000; 
        10'b0001001011: data <= 11'h7ff; 
        10'b0001001100: data <= 11'h001; 
        10'b0001001101: data <= 11'h000; 
        10'b0001001110: data <= 11'h000; 
        10'b0001001111: data <= 11'h001; 
        10'b0001010000: data <= 11'h000; 
        10'b0001010001: data <= 11'h000; 
        10'b0001010010: data <= 11'h000; 
        10'b0001010011: data <= 11'h001; 
        10'b0001010100: data <= 11'h002; 
        10'b0001010101: data <= 11'h000; 
        10'b0001010110: data <= 11'h000; 
        10'b0001010111: data <= 11'h000; 
        10'b0001011000: data <= 11'h001; 
        10'b0001011001: data <= 11'h7ff; 
        10'b0001011010: data <= 11'h001; 
        10'b0001011011: data <= 11'h001; 
        10'b0001011100: data <= 11'h000; 
        10'b0001011101: data <= 11'h001; 
        10'b0001011110: data <= 11'h000; 
        10'b0001011111: data <= 11'h001; 
        10'b0001100000: data <= 11'h000; 
        10'b0001100001: data <= 11'h7ff; 
        10'b0001100010: data <= 11'h000; 
        10'b0001100011: data <= 11'h7fe; 
        10'b0001100100: data <= 11'h000; 
        10'b0001100101: data <= 11'h7ff; 
        10'b0001100110: data <= 11'h000; 
        10'b0001100111: data <= 11'h000; 
        10'b0001101000: data <= 11'h000; 
        10'b0001101001: data <= 11'h000; 
        10'b0001101010: data <= 11'h001; 
        10'b0001101011: data <= 11'h000; 
        10'b0001101100: data <= 11'h000; 
        10'b0001101101: data <= 11'h001; 
        10'b0001101110: data <= 11'h001; 
        10'b0001101111: data <= 11'h001; 
        10'b0001110000: data <= 11'h000; 
        10'b0001110001: data <= 11'h000; 
        10'b0001110010: data <= 11'h000; 
        10'b0001110011: data <= 11'h000; 
        10'b0001110100: data <= 11'h7ff; 
        10'b0001110101: data <= 11'h001; 
        10'b0001110110: data <= 11'h001; 
        10'b0001110111: data <= 11'h000; 
        10'b0001111000: data <= 11'h7ff; 
        10'b0001111001: data <= 11'h000; 
        10'b0001111010: data <= 11'h7ff; 
        10'b0001111011: data <= 11'h7fe; 
        10'b0001111100: data <= 11'h7fd; 
        10'b0001111101: data <= 11'h7fb; 
        10'b0001111110: data <= 11'h7fa; 
        10'b0001111111: data <= 11'h7f8; 
        10'b0010000000: data <= 11'h7fa; 
        10'b0010000001: data <= 11'h7fa; 
        10'b0010000010: data <= 11'h7fb; 
        10'b0010000011: data <= 11'h7fe; 
        10'b0010000100: data <= 11'h7ff; 
        10'b0010000101: data <= 11'h7ff; 
        10'b0010000110: data <= 11'h000; 
        10'b0010000111: data <= 11'h001; 
        10'b0010001000: data <= 11'h001; 
        10'b0010001001: data <= 11'h001; 
        10'b0010001010: data <= 11'h000; 
        10'b0010001011: data <= 11'h000; 
        10'b0010001100: data <= 11'h001; 
        10'b0010001101: data <= 11'h001; 
        10'b0010001110: data <= 11'h001; 
        10'b0010001111: data <= 11'h001; 
        10'b0010010000: data <= 11'h001; 
        10'b0010010001: data <= 11'h7ff; 
        10'b0010010010: data <= 11'h7ff; 
        10'b0010010011: data <= 11'h7ff; 
        10'b0010010100: data <= 11'h7fd; 
        10'b0010010101: data <= 11'h7fd; 
        10'b0010010110: data <= 11'h7fd; 
        10'b0010010111: data <= 11'h7fc; 
        10'b0010011000: data <= 11'h7fb; 
        10'b0010011001: data <= 11'h7fa; 
        10'b0010011010: data <= 11'h7f7; 
        10'b0010011011: data <= 11'h7f6; 
        10'b0010011100: data <= 11'h7f4; 
        10'b0010011101: data <= 11'h7f8; 
        10'b0010011110: data <= 11'h7fb; 
        10'b0010011111: data <= 11'h7fe; 
        10'b0010100000: data <= 11'h7fd; 
        10'b0010100001: data <= 11'h7fd; 
        10'b0010100010: data <= 11'h7fd; 
        10'b0010100011: data <= 11'h7fe; 
        10'b0010100100: data <= 11'h7ff; 
        10'b0010100101: data <= 11'h000; 
        10'b0010100110: data <= 11'h000; 
        10'b0010100111: data <= 11'h001; 
        10'b0010101000: data <= 11'h001; 
        10'b0010101001: data <= 11'h001; 
        10'b0010101010: data <= 11'h7ff; 
        10'b0010101011: data <= 11'h001; 
        10'b0010101100: data <= 11'h001; 
        10'b0010101101: data <= 11'h7fd; 
        10'b0010101110: data <= 11'h7fc; 
        10'b0010101111: data <= 11'h7fc; 
        10'b0010110000: data <= 11'h7fb; 
        10'b0010110001: data <= 11'h7fa; 
        10'b0010110010: data <= 11'h7fc; 
        10'b0010110011: data <= 11'h7ff; 
        10'b0010110100: data <= 11'h000; 
        10'b0010110101: data <= 11'h005; 
        10'b0010110110: data <= 11'h008; 
        10'b0010110111: data <= 11'h006; 
        10'b0010111000: data <= 11'h004; 
        10'b0010111001: data <= 11'h004; 
        10'b0010111010: data <= 11'h005; 
        10'b0010111011: data <= 11'h7ff; 
        10'b0010111100: data <= 11'h7ff; 
        10'b0010111101: data <= 11'h7fc; 
        10'b0010111110: data <= 11'h7fa; 
        10'b0010111111: data <= 11'h7fa; 
        10'b0011000000: data <= 11'h7fd; 
        10'b0011000001: data <= 11'h7fe; 
        10'b0011000010: data <= 11'h000; 
        10'b0011000011: data <= 11'h001; 
        10'b0011000100: data <= 11'h002; 
        10'b0011000101: data <= 11'h000; 
        10'b0011000110: data <= 11'h7ff; 
        10'b0011000111: data <= 11'h7ff; 
        10'b0011001000: data <= 11'h7fd; 
        10'b0011001001: data <= 11'h7fb; 
        10'b0011001010: data <= 11'h7fa; 
        10'b0011001011: data <= 11'h7f9; 
        10'b0011001100: data <= 11'h7f9; 
        10'b0011001101: data <= 11'h7fe; 
        10'b0011001110: data <= 11'h000; 
        10'b0011001111: data <= 11'h002; 
        10'b0011010000: data <= 11'h007; 
        10'b0011010001: data <= 11'h009; 
        10'b0011010010: data <= 11'h00c; 
        10'b0011010011: data <= 11'h00c; 
        10'b0011010100: data <= 11'h00d; 
        10'b0011010101: data <= 11'h006; 
        10'b0011010110: data <= 11'h004; 
        10'b0011010111: data <= 11'h000; 
        10'b0011011000: data <= 11'h001; 
        10'b0011011001: data <= 11'h001; 
        10'b0011011010: data <= 11'h7fc; 
        10'b0011011011: data <= 11'h7f8; 
        10'b0011011100: data <= 11'h7fb; 
        10'b0011011101: data <= 11'h7ff; 
        10'b0011011110: data <= 11'h7ff; 
        10'b0011011111: data <= 11'h001; 
        10'b0011100000: data <= 11'h002; 
        10'b0011100001: data <= 11'h002; 
        10'b0011100010: data <= 11'h001; 
        10'b0011100011: data <= 11'h000; 
        10'b0011100100: data <= 11'h7fc; 
        10'b0011100101: data <= 11'h7fb; 
        10'b0011100110: data <= 11'h7fa; 
        10'b0011100111: data <= 11'h7f7; 
        10'b0011101000: data <= 11'h7fe; 
        10'b0011101001: data <= 11'h7ff; 
        10'b0011101010: data <= 11'h7ff; 
        10'b0011101011: data <= 11'h7fd; 
        10'b0011101100: data <= 11'h000; 
        10'b0011101101: data <= 11'h004; 
        10'b0011101110: data <= 11'h00a; 
        10'b0011101111: data <= 11'h006; 
        10'b0011110000: data <= 11'h006; 
        10'b0011110001: data <= 11'h001; 
        10'b0011110010: data <= 11'h000; 
        10'b0011110011: data <= 11'h000; 
        10'b0011110100: data <= 11'h7fe; 
        10'b0011110101: data <= 11'h001; 
        10'b0011110110: data <= 11'h7fe; 
        10'b0011110111: data <= 11'h7fa; 
        10'b0011111000: data <= 11'h7fb; 
        10'b0011111001: data <= 11'h7fd; 
        10'b0011111010: data <= 11'h7ff; 
        10'b0011111011: data <= 11'h001; 
        10'b0011111100: data <= 11'h000; 
        10'b0011111101: data <= 11'h000; 
        10'b0011111110: data <= 11'h000; 
        10'b0011111111: data <= 11'h7fd; 
        10'b0100000000: data <= 11'h7fa; 
        10'b0100000001: data <= 11'h7fc; 
        10'b0100000010: data <= 11'h7ff; 
        10'b0100000011: data <= 11'h7fe; 
        10'b0100000100: data <= 11'h7ff; 
        10'b0100000101: data <= 11'h7ff; 
        10'b0100000110: data <= 11'h003; 
        10'b0100000111: data <= 11'h002; 
        10'b0100001000: data <= 11'h000; 
        10'b0100001001: data <= 11'h004; 
        10'b0100001010: data <= 11'h007; 
        10'b0100001011: data <= 11'h006; 
        10'b0100001100: data <= 11'h000; 
        10'b0100001101: data <= 11'h7fe; 
        10'b0100001110: data <= 11'h000; 
        10'b0100001111: data <= 11'h7fc; 
        10'b0100010000: data <= 11'h7fe; 
        10'b0100010001: data <= 11'h7fc; 
        10'b0100010010: data <= 11'h7fc; 
        10'b0100010011: data <= 11'h7fb; 
        10'b0100010100: data <= 11'h7fd; 
        10'b0100010101: data <= 11'h7ff; 
        10'b0100010110: data <= 11'h7ff; 
        10'b0100010111: data <= 11'h001; 
        10'b0100011000: data <= 11'h000; 
        10'b0100011001: data <= 11'h000; 
        10'b0100011010: data <= 11'h7ff; 
        10'b0100011011: data <= 11'h7ff; 
        10'b0100011100: data <= 11'h7fc; 
        10'b0100011101: data <= 11'h7fe; 
        10'b0100011110: data <= 11'h002; 
        10'b0100011111: data <= 11'h003; 
        10'b0100100000: data <= 11'h006; 
        10'b0100100001: data <= 11'h006; 
        10'b0100100010: data <= 11'h005; 
        10'b0100100011: data <= 11'h007; 
        10'b0100100100: data <= 11'h004; 
        10'b0100100101: data <= 11'h001; 
        10'b0100100110: data <= 11'h001; 
        10'b0100100111: data <= 11'h7fc; 
        10'b0100101000: data <= 11'h7fe; 
        10'b0100101001: data <= 11'h000; 
        10'b0100101010: data <= 11'h003; 
        10'b0100101011: data <= 11'h000; 
        10'b0100101100: data <= 11'h002; 
        10'b0100101101: data <= 11'h7ff; 
        10'b0100101110: data <= 11'h7fd; 
        10'b0100101111: data <= 11'h7fe; 
        10'b0100110000: data <= 11'h7fd; 
        10'b0100110001: data <= 11'h7ff; 
        10'b0100110010: data <= 11'h7ff; 
        10'b0100110011: data <= 11'h001; 
        10'b0100110100: data <= 11'h000; 
        10'b0100110101: data <= 11'h000; 
        10'b0100110110: data <= 11'h7ff; 
        10'b0100110111: data <= 11'h000; 
        10'b0100111000: data <= 11'h7ff; 
        10'b0100111001: data <= 11'h004; 
        10'b0100111010: data <= 11'h009; 
        10'b0100111011: data <= 11'h007; 
        10'b0100111100: data <= 11'h00b; 
        10'b0100111101: data <= 11'h004; 
        10'b0100111110: data <= 11'h004; 
        10'b0100111111: data <= 11'h008; 
        10'b0101000000: data <= 11'h7fe; 
        10'b0101000001: data <= 11'h7fe; 
        10'b0101000010: data <= 11'h7ff; 
        10'b0101000011: data <= 11'h001; 
        10'b0101000100: data <= 11'h003; 
        10'b0101000101: data <= 11'h00a; 
        10'b0101000110: data <= 11'h005; 
        10'b0101000111: data <= 11'h005; 
        10'b0101001000: data <= 11'h008; 
        10'b0101001001: data <= 11'h006; 
        10'b0101001010: data <= 11'h003; 
        10'b0101001011: data <= 11'h001; 
        10'b0101001100: data <= 11'h7ff; 
        10'b0101001101: data <= 11'h7ff; 
        10'b0101001110: data <= 11'h000; 
        10'b0101001111: data <= 11'h000; 
        10'b0101010000: data <= 11'h001; 
        10'b0101010001: data <= 11'h001; 
        10'b0101010010: data <= 11'h7ff; 
        10'b0101010011: data <= 11'h7ff; 
        10'b0101010100: data <= 11'h003; 
        10'b0101010101: data <= 11'h009; 
        10'b0101010110: data <= 11'h00a; 
        10'b0101010111: data <= 11'h006; 
        10'b0101011000: data <= 11'h007; 
        10'b0101011001: data <= 11'h009; 
        10'b0101011010: data <= 11'h006; 
        10'b0101011011: data <= 11'h000; 
        10'b0101011100: data <= 11'h7fa; 
        10'b0101011101: data <= 11'h005; 
        10'b0101011110: data <= 11'h00b; 
        10'b0101011111: data <= 11'h009; 
        10'b0101100000: data <= 11'h007; 
        10'b0101100001: data <= 11'h00b; 
        10'b0101100010: data <= 11'h00b; 
        10'b0101100011: data <= 11'h00c; 
        10'b0101100100: data <= 11'h00c; 
        10'b0101100101: data <= 11'h008; 
        10'b0101100110: data <= 11'h004; 
        10'b0101100111: data <= 11'h000; 
        10'b0101101000: data <= 11'h7fe; 
        10'b0101101001: data <= 11'h000; 
        10'b0101101010: data <= 11'h001; 
        10'b0101101011: data <= 11'h001; 
        10'b0101101100: data <= 11'h002; 
        10'b0101101101: data <= 11'h001; 
        10'b0101101110: data <= 11'h7ff; 
        10'b0101101111: data <= 11'h000; 
        10'b0101110000: data <= 11'h005; 
        10'b0101110001: data <= 11'h008; 
        10'b0101110010: data <= 11'h007; 
        10'b0101110011: data <= 11'h005; 
        10'b0101110100: data <= 11'h006; 
        10'b0101110101: data <= 11'h004; 
        10'b0101110110: data <= 11'h003; 
        10'b0101110111: data <= 11'h7fe; 
        10'b0101111000: data <= 11'h7fd; 
        10'b0101111001: data <= 11'h008; 
        10'b0101111010: data <= 11'h00b; 
        10'b0101111011: data <= 11'h008; 
        10'b0101111100: data <= 11'h009; 
        10'b0101111101: data <= 11'h008; 
        10'b0101111110: data <= 11'h00b; 
        10'b0101111111: data <= 11'h00b; 
        10'b0110000000: data <= 11'h009; 
        10'b0110000001: data <= 11'h005; 
        10'b0110000010: data <= 11'h000; 
        10'b0110000011: data <= 11'h7fc; 
        10'b0110000100: data <= 11'h7fe; 
        10'b0110000101: data <= 11'h7ff; 
        10'b0110000110: data <= 11'h001; 
        10'b0110000111: data <= 11'h001; 
        10'b0110001000: data <= 11'h000; 
        10'b0110001001: data <= 11'h000; 
        10'b0110001010: data <= 11'h001; 
        10'b0110001011: data <= 11'h001; 
        10'b0110001100: data <= 11'h002; 
        10'b0110001101: data <= 11'h002; 
        10'b0110001110: data <= 11'h006; 
        10'b0110001111: data <= 11'h004; 
        10'b0110010000: data <= 11'h002; 
        10'b0110010001: data <= 11'h000; 
        10'b0110010010: data <= 11'h001; 
        10'b0110010011: data <= 11'h000; 
        10'b0110010100: data <= 11'h7fe; 
        10'b0110010101: data <= 11'h003; 
        10'b0110010110: data <= 11'h001; 
        10'b0110010111: data <= 11'h007; 
        10'b0110011000: data <= 11'h007; 
        10'b0110011001: data <= 11'h007; 
        10'b0110011010: data <= 11'h005; 
        10'b0110011011: data <= 11'h003; 
        10'b0110011100: data <= 11'h004; 
        10'b0110011101: data <= 11'h000; 
        10'b0110011110: data <= 11'h7fc; 
        10'b0110011111: data <= 11'h7fa; 
        10'b0110100000: data <= 11'h7fe; 
        10'b0110100001: data <= 11'h000; 
        10'b0110100010: data <= 11'h000; 
        10'b0110100011: data <= 11'h000; 
        10'b0110100100: data <= 11'h001; 
        10'b0110100101: data <= 11'h001; 
        10'b0110100110: data <= 11'h001; 
        10'b0110100111: data <= 11'h7ff; 
        10'b0110101000: data <= 11'h000; 
        10'b0110101001: data <= 11'h003; 
        10'b0110101010: data <= 11'h003; 
        10'b0110101011: data <= 11'h002; 
        10'b0110101100: data <= 11'h002; 
        10'b0110101101: data <= 11'h7fd; 
        10'b0110101110: data <= 11'h7ff; 
        10'b0110101111: data <= 11'h7ff; 
        10'b0110110000: data <= 11'h7fe; 
        10'b0110110001: data <= 11'h7fe; 
        10'b0110110010: data <= 11'h7fe; 
        10'b0110110011: data <= 11'h008; 
        10'b0110110100: data <= 11'h00b; 
        10'b0110110101: data <= 11'h00b; 
        10'b0110110110: data <= 11'h005; 
        10'b0110110111: data <= 11'h001; 
        10'b0110111000: data <= 11'h7fe; 
        10'b0110111001: data <= 11'h7fa; 
        10'b0110111010: data <= 11'h7f8; 
        10'b0110111011: data <= 11'h7fb; 
        10'b0110111100: data <= 11'h7fe; 
        10'b0110111101: data <= 11'h000; 
        10'b0110111110: data <= 11'h001; 
        10'b0110111111: data <= 11'h000; 
        10'b0111000000: data <= 11'h001; 
        10'b0111000001: data <= 11'h000; 
        10'b0111000010: data <= 11'h7ff; 
        10'b0111000011: data <= 11'h000; 
        10'b0111000100: data <= 11'h000; 
        10'b0111000101: data <= 11'h001; 
        10'b0111000110: data <= 11'h7fe; 
        10'b0111000111: data <= 11'h002; 
        10'b0111001000: data <= 11'h005; 
        10'b0111001001: data <= 11'h7ff; 
        10'b0111001010: data <= 11'h003; 
        10'b0111001011: data <= 11'h004; 
        10'b0111001100: data <= 11'h7ff; 
        10'b0111001101: data <= 11'h7fc; 
        10'b0111001110: data <= 11'h7ff; 
        10'b0111001111: data <= 11'h004; 
        10'b0111010000: data <= 11'h008; 
        10'b0111010001: data <= 11'h008; 
        10'b0111010010: data <= 11'h002; 
        10'b0111010011: data <= 11'h7fc; 
        10'b0111010100: data <= 11'h7f9; 
        10'b0111010101: data <= 11'h7f6; 
        10'b0111010110: data <= 11'h7f9; 
        10'b0111010111: data <= 11'h7fa; 
        10'b0111011000: data <= 11'h7fc; 
        10'b0111011001: data <= 11'h000; 
        10'b0111011010: data <= 11'h7ff; 
        10'b0111011011: data <= 11'h001; 
        10'b0111011100: data <= 11'h000; 
        10'b0111011101: data <= 11'h000; 
        10'b0111011110: data <= 11'h7ff; 
        10'b0111011111: data <= 11'h7fe; 
        10'b0111100000: data <= 11'h7fd; 
        10'b0111100001: data <= 11'h7fd; 
        10'b0111100010: data <= 11'h7fd; 
        10'b0111100011: data <= 11'h001; 
        10'b0111100100: data <= 11'h002; 
        10'b0111100101: data <= 11'h003; 
        10'b0111100110: data <= 11'h004; 
        10'b0111100111: data <= 11'h006; 
        10'b0111101000: data <= 11'h004; 
        10'b0111101001: data <= 11'h002; 
        10'b0111101010: data <= 11'h002; 
        10'b0111101011: data <= 11'h006; 
        10'b0111101100: data <= 11'h002; 
        10'b0111101101: data <= 11'h7ff; 
        10'b0111101110: data <= 11'h7fd; 
        10'b0111101111: data <= 11'h7fa; 
        10'b0111110000: data <= 11'h7fa; 
        10'b0111110001: data <= 11'h7f9; 
        10'b0111110010: data <= 11'h7fa; 
        10'b0111110011: data <= 11'h7fb; 
        10'b0111110100: data <= 11'h7fd; 
        10'b0111110101: data <= 11'h000; 
        10'b0111110110: data <= 11'h000; 
        10'b0111110111: data <= 11'h000; 
        10'b0111111000: data <= 11'h001; 
        10'b0111111001: data <= 11'h000; 
        10'b0111111010: data <= 11'h7ff; 
        10'b0111111011: data <= 11'h000; 
        10'b0111111100: data <= 11'h7fe; 
        10'b0111111101: data <= 11'h7fa; 
        10'b0111111110: data <= 11'h7fa; 
        10'b0111111111: data <= 11'h7fa; 
        10'b1000000000: data <= 11'h7fe; 
        10'b1000000001: data <= 11'h001; 
        10'b1000000010: data <= 11'h007; 
        10'b1000000011: data <= 11'h006; 
        10'b1000000100: data <= 11'h7fd; 
        10'b1000000101: data <= 11'h7fd; 
        10'b1000000110: data <= 11'h000; 
        10'b1000000111: data <= 11'h004; 
        10'b1000001000: data <= 11'h7fd; 
        10'b1000001001: data <= 11'h7fd; 
        10'b1000001010: data <= 11'h7fb; 
        10'b1000001011: data <= 11'h7fd; 
        10'b1000001100: data <= 11'h7fd; 
        10'b1000001101: data <= 11'h7fb; 
        10'b1000001110: data <= 11'h7fb; 
        10'b1000001111: data <= 11'h7fb; 
        10'b1000010000: data <= 11'h7fc; 
        10'b1000010001: data <= 11'h7ff; 
        10'b1000010010: data <= 11'h000; 
        10'b1000010011: data <= 11'h001; 
        10'b1000010100: data <= 11'h001; 
        10'b1000010101: data <= 11'h002; 
        10'b1000010110: data <= 11'h000; 
        10'b1000010111: data <= 11'h7ff; 
        10'b1000011000: data <= 11'h7fe; 
        10'b1000011001: data <= 11'h7fc; 
        10'b1000011010: data <= 11'h7fa; 
        10'b1000011011: data <= 11'h7f9; 
        10'b1000011100: data <= 11'h7f9; 
        10'b1000011101: data <= 11'h7f9; 
        10'b1000011110: data <= 11'h7f9; 
        10'b1000011111: data <= 11'h7fa; 
        10'b1000100000: data <= 11'h7f8; 
        10'b1000100001: data <= 11'h7fa; 
        10'b1000100010: data <= 11'h7fb; 
        10'b1000100011: data <= 11'h7fb; 
        10'b1000100100: data <= 11'h7fb; 
        10'b1000100101: data <= 11'h7fe; 
        10'b1000100110: data <= 11'h7fc; 
        10'b1000100111: data <= 11'h7ff; 
        10'b1000101000: data <= 11'h7fe; 
        10'b1000101001: data <= 11'h7fd; 
        10'b1000101010: data <= 11'h7fd; 
        10'b1000101011: data <= 11'h7fe; 
        10'b1000101100: data <= 11'h7fe; 
        10'b1000101101: data <= 11'h000; 
        10'b1000101110: data <= 11'h000; 
        10'b1000101111: data <= 11'h000; 
        10'b1000110000: data <= 11'h000; 
        10'b1000110001: data <= 11'h000; 
        10'b1000110010: data <= 11'h001; 
        10'b1000110011: data <= 11'h000; 
        10'b1000110100: data <= 11'h7fe; 
        10'b1000110101: data <= 11'h7fc; 
        10'b1000110110: data <= 11'h7fa; 
        10'b1000110111: data <= 11'h7f7; 
        10'b1000111000: data <= 11'h7f5; 
        10'b1000111001: data <= 11'h7f4; 
        10'b1000111010: data <= 11'h7f0; 
        10'b1000111011: data <= 11'h7f4; 
        10'b1000111100: data <= 11'h7f4; 
        10'b1000111101: data <= 11'h7fc; 
        10'b1000111110: data <= 11'h7fb; 
        10'b1000111111: data <= 11'h7fd; 
        10'b1001000000: data <= 11'h7fd; 
        10'b1001000001: data <= 11'h7ff; 
        10'b1001000010: data <= 11'h7fb; 
        10'b1001000011: data <= 11'h7fe; 
        10'b1001000100: data <= 11'h7fe; 
        10'b1001000101: data <= 11'h7fd; 
        10'b1001000110: data <= 11'h7ff; 
        10'b1001000111: data <= 11'h7fe; 
        10'b1001001000: data <= 11'h000; 
        10'b1001001001: data <= 11'h001; 
        10'b1001001010: data <= 11'h001; 
        10'b1001001011: data <= 11'h000; 
        10'b1001001100: data <= 11'h000; 
        10'b1001001101: data <= 11'h000; 
        10'b1001001110: data <= 11'h001; 
        10'b1001001111: data <= 11'h7ff; 
        10'b1001010000: data <= 11'h7fe; 
        10'b1001010001: data <= 11'h7fc; 
        10'b1001010010: data <= 11'h7fb; 
        10'b1001010011: data <= 11'h7f8; 
        10'b1001010100: data <= 11'h7f7; 
        10'b1001010101: data <= 11'h7f6; 
        10'b1001010110: data <= 11'h7f5; 
        10'b1001010111: data <= 11'h7f6; 
        10'b1001011000: data <= 11'h7fa; 
        10'b1001011001: data <= 11'h7fa; 
        10'b1001011010: data <= 11'h7fa; 
        10'b1001011011: data <= 11'h7fc; 
        10'b1001011100: data <= 11'h7fc; 
        10'b1001011101: data <= 11'h7fa; 
        10'b1001011110: data <= 11'h7f9; 
        10'b1001011111: data <= 11'h7fd; 
        10'b1001100000: data <= 11'h7fe; 
        10'b1001100001: data <= 11'h7ff; 
        10'b1001100010: data <= 11'h000; 
        10'b1001100011: data <= 11'h000; 
        10'b1001100100: data <= 11'h001; 
        10'b1001100101: data <= 11'h001; 
        10'b1001100110: data <= 11'h000; 
        10'b1001100111: data <= 11'h000; 
        10'b1001101000: data <= 11'h001; 
        10'b1001101001: data <= 11'h000; 
        10'b1001101010: data <= 11'h000; 
        10'b1001101011: data <= 11'h001; 
        10'b1001101100: data <= 11'h7ff; 
        10'b1001101101: data <= 11'h7fd; 
        10'b1001101110: data <= 11'h7fb; 
        10'b1001101111: data <= 11'h7f9; 
        10'b1001110000: data <= 11'h7fb; 
        10'b1001110001: data <= 11'h7fb; 
        10'b1001110010: data <= 11'h7fa; 
        10'b1001110011: data <= 11'h7fc; 
        10'b1001110100: data <= 11'h7fc; 
        10'b1001110101: data <= 11'h7fa; 
        10'b1001110110: data <= 11'h7fb; 
        10'b1001110111: data <= 11'h7f9; 
        10'b1001111000: data <= 11'h7f8; 
        10'b1001111001: data <= 11'h7f9; 
        10'b1001111010: data <= 11'h7fa; 
        10'b1001111011: data <= 11'h7fb; 
        10'b1001111100: data <= 11'h7ff; 
        10'b1001111101: data <= 11'h002; 
        10'b1001111110: data <= 11'h001; 
        10'b1001111111: data <= 11'h001; 
        10'b1010000000: data <= 11'h002; 
        10'b1010000001: data <= 11'h000; 
        10'b1010000010: data <= 11'h000; 
        10'b1010000011: data <= 11'h001; 
        10'b1010000100: data <= 11'h001; 
        10'b1010000101: data <= 11'h001; 
        10'b1010000110: data <= 11'h000; 
        10'b1010000111: data <= 11'h000; 
        10'b1010001000: data <= 11'h7ff; 
        10'b1010001001: data <= 11'h7fd; 
        10'b1010001010: data <= 11'h7fd; 
        10'b1010001011: data <= 11'h7fc; 
        10'b1010001100: data <= 11'h000; 
        10'b1010001101: data <= 11'h7fe; 
        10'b1010001110: data <= 11'h7ff; 
        10'b1010001111: data <= 11'h7fb; 
        10'b1010010000: data <= 11'h7fc; 
        10'b1010010001: data <= 11'h7fb; 
        10'b1010010010: data <= 11'h7fc; 
        10'b1010010011: data <= 11'h7f9; 
        10'b1010010100: data <= 11'h7f8; 
        10'b1010010101: data <= 11'h7f9; 
        10'b1010010110: data <= 11'h7fc; 
        10'b1010010111: data <= 11'h000; 
        10'b1010011000: data <= 11'h002; 
        10'b1010011001: data <= 11'h004; 
        10'b1010011010: data <= 11'h006; 
        10'b1010011011: data <= 11'h005; 
        10'b1010011100: data <= 11'h002; 
        10'b1010011101: data <= 11'h000; 
        10'b1010011110: data <= 11'h002; 
        10'b1010011111: data <= 11'h000; 
        10'b1010100000: data <= 11'h000; 
        10'b1010100001: data <= 11'h7ff; 
        10'b1010100010: data <= 11'h000; 
        10'b1010100011: data <= 11'h001; 
        10'b1010100100: data <= 11'h001; 
        10'b1010100101: data <= 11'h002; 
        10'b1010100110: data <= 11'h001; 
        10'b1010100111: data <= 11'h002; 
        10'b1010101000: data <= 11'h002; 
        10'b1010101001: data <= 11'h001; 
        10'b1010101010: data <= 11'h7ff; 
        10'b1010101011: data <= 11'h7fd; 
        10'b1010101100: data <= 11'h000; 
        10'b1010101101: data <= 11'h7fc; 
        10'b1010101110: data <= 11'h7fb; 
        10'b1010101111: data <= 11'h7fb; 
        10'b1010110000: data <= 11'h7fe; 
        10'b1010110001: data <= 11'h002; 
        10'b1010110010: data <= 11'h003; 
        10'b1010110011: data <= 11'h003; 
        10'b1010110100: data <= 11'h007; 
        10'b1010110101: data <= 11'h007; 
        10'b1010110110: data <= 11'h004; 
        10'b1010110111: data <= 11'h003; 
        10'b1010111000: data <= 11'h002; 
        10'b1010111001: data <= 11'h000; 
        10'b1010111010: data <= 11'h001; 
        10'b1010111011: data <= 11'h000; 
        10'b1010111100: data <= 11'h000; 
        10'b1010111101: data <= 11'h001; 
        10'b1010111110: data <= 11'h001; 
        10'b1010111111: data <= 11'h000; 
        10'b1011000000: data <= 11'h000; 
        10'b1011000001: data <= 11'h002; 
        10'b1011000010: data <= 11'h002; 
        10'b1011000011: data <= 11'h005; 
        10'b1011000100: data <= 11'h005; 
        10'b1011000101: data <= 11'h006; 
        10'b1011000110: data <= 11'h005; 
        10'b1011000111: data <= 11'h002; 
        10'b1011001000: data <= 11'h005; 
        10'b1011001001: data <= 11'h005; 
        10'b1011001010: data <= 11'h004; 
        10'b1011001011: data <= 11'h004; 
        10'b1011001100: data <= 11'h008; 
        10'b1011001101: data <= 11'h008; 
        10'b1011001110: data <= 11'h009; 
        10'b1011001111: data <= 11'h00a; 
        10'b1011010000: data <= 11'h00b; 
        10'b1011010001: data <= 11'h008; 
        10'b1011010010: data <= 11'h003; 
        10'b1011010011: data <= 11'h001; 
        10'b1011010100: data <= 11'h000; 
        10'b1011010101: data <= 11'h000; 
        10'b1011010110: data <= 11'h000; 
        10'b1011010111: data <= 11'h000; 
        10'b1011011000: data <= 11'h000; 
        10'b1011011001: data <= 11'h001; 
        10'b1011011010: data <= 11'h000; 
        10'b1011011011: data <= 11'h000; 
        10'b1011011100: data <= 11'h001; 
        10'b1011011101: data <= 11'h002; 
        10'b1011011110: data <= 11'h003; 
        10'b1011011111: data <= 11'h004; 
        10'b1011100000: data <= 11'h004; 
        10'b1011100001: data <= 11'h006; 
        10'b1011100010: data <= 11'h007; 
        10'b1011100011: data <= 11'h007; 
        10'b1011100100: data <= 11'h009; 
        10'b1011100101: data <= 11'h009; 
        10'b1011100110: data <= 11'h00b; 
        10'b1011100111: data <= 11'h006; 
        10'b1011101000: data <= 11'h004; 
        10'b1011101001: data <= 11'h004; 
        10'b1011101010: data <= 11'h005; 
        10'b1011101011: data <= 11'h006; 
        10'b1011101100: data <= 11'h004; 
        10'b1011101101: data <= 11'h003; 
        10'b1011101110: data <= 11'h001; 
        10'b1011101111: data <= 11'h000; 
        10'b1011110000: data <= 11'h000; 
        10'b1011110001: data <= 11'h000; 
        10'b1011110010: data <= 11'h000; 
        10'b1011110011: data <= 11'h000; 
        10'b1011110100: data <= 11'h000; 
        10'b1011110101: data <= 11'h001; 
        10'b1011110110: data <= 11'h7ff; 
        10'b1011110111: data <= 11'h001; 
        10'b1011111000: data <= 11'h001; 
        10'b1011111001: data <= 11'h000; 
        10'b1011111010: data <= 11'h000; 
        10'b1011111011: data <= 11'h001; 
        10'b1011111100: data <= 11'h001; 
        10'b1011111101: data <= 11'h001; 
        10'b1011111110: data <= 11'h000; 
        10'b1011111111: data <= 11'h000; 
        10'b1100000000: data <= 11'h000; 
        10'b1100000001: data <= 11'h000; 
        10'b1100000010: data <= 11'h000; 
        10'b1100000011: data <= 11'h001; 
        10'b1100000100: data <= 11'h000; 
        10'b1100000101: data <= 11'h001; 
        10'b1100000110: data <= 11'h002; 
        10'b1100000111: data <= 11'h001; 
        10'b1100001000: data <= 11'h001; 
        10'b1100001001: data <= 11'h001; 
        10'b1100001010: data <= 11'h000; 
        10'b1100001011: data <= 11'h002; 
        10'b1100001100: data <= 11'h001; 
        10'b1100001101: data <= 11'h000; 
        10'b1100001110: data <= 11'h000; 
        10'b1100001111: data <= 11'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 6) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 12'h002; 
        10'b0000000001: data <= 12'h002; 
        10'b0000000010: data <= 12'hfff; 
        10'b0000000011: data <= 12'h001; 
        10'b0000000100: data <= 12'h001; 
        10'b0000000101: data <= 12'h002; 
        10'b0000000110: data <= 12'hfff; 
        10'b0000000111: data <= 12'h000; 
        10'b0000001000: data <= 12'h002; 
        10'b0000001001: data <= 12'hfff; 
        10'b0000001010: data <= 12'h000; 
        10'b0000001011: data <= 12'h001; 
        10'b0000001100: data <= 12'h003; 
        10'b0000001101: data <= 12'h002; 
        10'b0000001110: data <= 12'hfff; 
        10'b0000001111: data <= 12'hfff; 
        10'b0000010000: data <= 12'hfff; 
        10'b0000010001: data <= 12'h001; 
        10'b0000010010: data <= 12'h002; 
        10'b0000010011: data <= 12'h000; 
        10'b0000010100: data <= 12'h000; 
        10'b0000010101: data <= 12'h000; 
        10'b0000010110: data <= 12'hfff; 
        10'b0000010111: data <= 12'h000; 
        10'b0000011000: data <= 12'h002; 
        10'b0000011001: data <= 12'h001; 
        10'b0000011010: data <= 12'hfff; 
        10'b0000011011: data <= 12'h001; 
        10'b0000011100: data <= 12'h002; 
        10'b0000011101: data <= 12'h002; 
        10'b0000011110: data <= 12'h001; 
        10'b0000011111: data <= 12'h000; 
        10'b0000100000: data <= 12'hfff; 
        10'b0000100001: data <= 12'hfff; 
        10'b0000100010: data <= 12'h000; 
        10'b0000100011: data <= 12'h003; 
        10'b0000100100: data <= 12'hfff; 
        10'b0000100101: data <= 12'h002; 
        10'b0000100110: data <= 12'h001; 
        10'b0000100111: data <= 12'h002; 
        10'b0000101000: data <= 12'h001; 
        10'b0000101001: data <= 12'h002; 
        10'b0000101010: data <= 12'h000; 
        10'b0000101011: data <= 12'hfff; 
        10'b0000101100: data <= 12'hfff; 
        10'b0000101101: data <= 12'h002; 
        10'b0000101110: data <= 12'h000; 
        10'b0000101111: data <= 12'h001; 
        10'b0000110000: data <= 12'h002; 
        10'b0000110001: data <= 12'h000; 
        10'b0000110010: data <= 12'h000; 
        10'b0000110011: data <= 12'h000; 
        10'b0000110100: data <= 12'h001; 
        10'b0000110101: data <= 12'h003; 
        10'b0000110110: data <= 12'h000; 
        10'b0000110111: data <= 12'h001; 
        10'b0000111000: data <= 12'h003; 
        10'b0000111001: data <= 12'h003; 
        10'b0000111010: data <= 12'h000; 
        10'b0000111011: data <= 12'h002; 
        10'b0000111100: data <= 12'h002; 
        10'b0000111101: data <= 12'h000; 
        10'b0000111110: data <= 12'h000; 
        10'b0000111111: data <= 12'h001; 
        10'b0001000000: data <= 12'h002; 
        10'b0001000001: data <= 12'h000; 
        10'b0001000010: data <= 12'hfff; 
        10'b0001000011: data <= 12'h002; 
        10'b0001000100: data <= 12'h001; 
        10'b0001000101: data <= 12'h002; 
        10'b0001000110: data <= 12'hfff; 
        10'b0001000111: data <= 12'h002; 
        10'b0001001000: data <= 12'hfff; 
        10'b0001001001: data <= 12'hfff; 
        10'b0001001010: data <= 12'h000; 
        10'b0001001011: data <= 12'hfff; 
        10'b0001001100: data <= 12'h003; 
        10'b0001001101: data <= 12'hfff; 
        10'b0001001110: data <= 12'hfff; 
        10'b0001001111: data <= 12'h003; 
        10'b0001010000: data <= 12'h000; 
        10'b0001010001: data <= 12'h000; 
        10'b0001010010: data <= 12'h001; 
        10'b0001010011: data <= 12'h001; 
        10'b0001010100: data <= 12'h003; 
        10'b0001010101: data <= 12'h000; 
        10'b0001010110: data <= 12'h000; 
        10'b0001010111: data <= 12'h001; 
        10'b0001011000: data <= 12'h001; 
        10'b0001011001: data <= 12'hfff; 
        10'b0001011010: data <= 12'h003; 
        10'b0001011011: data <= 12'h001; 
        10'b0001011100: data <= 12'hfff; 
        10'b0001011101: data <= 12'h003; 
        10'b0001011110: data <= 12'h001; 
        10'b0001011111: data <= 12'h002; 
        10'b0001100000: data <= 12'h000; 
        10'b0001100001: data <= 12'hffe; 
        10'b0001100010: data <= 12'h000; 
        10'b0001100011: data <= 12'hffc; 
        10'b0001100100: data <= 12'h000; 
        10'b0001100101: data <= 12'hffe; 
        10'b0001100110: data <= 12'h001; 
        10'b0001100111: data <= 12'h000; 
        10'b0001101000: data <= 12'h001; 
        10'b0001101001: data <= 12'h000; 
        10'b0001101010: data <= 12'h002; 
        10'b0001101011: data <= 12'h000; 
        10'b0001101100: data <= 12'h000; 
        10'b0001101101: data <= 12'h003; 
        10'b0001101110: data <= 12'h001; 
        10'b0001101111: data <= 12'h002; 
        10'b0001110000: data <= 12'h000; 
        10'b0001110001: data <= 12'h001; 
        10'b0001110010: data <= 12'h000; 
        10'b0001110011: data <= 12'hfff; 
        10'b0001110100: data <= 12'hfff; 
        10'b0001110101: data <= 12'h002; 
        10'b0001110110: data <= 12'h001; 
        10'b0001110111: data <= 12'h000; 
        10'b0001111000: data <= 12'hffe; 
        10'b0001111001: data <= 12'h001; 
        10'b0001111010: data <= 12'hffd; 
        10'b0001111011: data <= 12'hffc; 
        10'b0001111100: data <= 12'hffb; 
        10'b0001111101: data <= 12'hff6; 
        10'b0001111110: data <= 12'hff3; 
        10'b0001111111: data <= 12'hfef; 
        10'b0010000000: data <= 12'hff4; 
        10'b0010000001: data <= 12'hff4; 
        10'b0010000010: data <= 12'hff7; 
        10'b0010000011: data <= 12'hffc; 
        10'b0010000100: data <= 12'hffe; 
        10'b0010000101: data <= 12'hfff; 
        10'b0010000110: data <= 12'h000; 
        10'b0010000111: data <= 12'h002; 
        10'b0010001000: data <= 12'h002; 
        10'b0010001001: data <= 12'h002; 
        10'b0010001010: data <= 12'h000; 
        10'b0010001011: data <= 12'h000; 
        10'b0010001100: data <= 12'h002; 
        10'b0010001101: data <= 12'h002; 
        10'b0010001110: data <= 12'h002; 
        10'b0010001111: data <= 12'h001; 
        10'b0010010000: data <= 12'h001; 
        10'b0010010001: data <= 12'hffe; 
        10'b0010010010: data <= 12'hffe; 
        10'b0010010011: data <= 12'hffe; 
        10'b0010010100: data <= 12'hffa; 
        10'b0010010101: data <= 12'hffa; 
        10'b0010010110: data <= 12'hffa; 
        10'b0010010111: data <= 12'hff8; 
        10'b0010011000: data <= 12'hff6; 
        10'b0010011001: data <= 12'hff4; 
        10'b0010011010: data <= 12'hfee; 
        10'b0010011011: data <= 12'hfed; 
        10'b0010011100: data <= 12'hfe8; 
        10'b0010011101: data <= 12'hff0; 
        10'b0010011110: data <= 12'hff6; 
        10'b0010011111: data <= 12'hffb; 
        10'b0010100000: data <= 12'hffb; 
        10'b0010100001: data <= 12'hff9; 
        10'b0010100010: data <= 12'hffa; 
        10'b0010100011: data <= 12'hffc; 
        10'b0010100100: data <= 12'hffe; 
        10'b0010100101: data <= 12'hfff; 
        10'b0010100110: data <= 12'h000; 
        10'b0010100111: data <= 12'h002; 
        10'b0010101000: data <= 12'h002; 
        10'b0010101001: data <= 12'h002; 
        10'b0010101010: data <= 12'hfff; 
        10'b0010101011: data <= 12'h002; 
        10'b0010101100: data <= 12'h001; 
        10'b0010101101: data <= 12'hffa; 
        10'b0010101110: data <= 12'hff9; 
        10'b0010101111: data <= 12'hff7; 
        10'b0010110000: data <= 12'hff6; 
        10'b0010110001: data <= 12'hff4; 
        10'b0010110010: data <= 12'hff7; 
        10'b0010110011: data <= 12'hffd; 
        10'b0010110100: data <= 12'h001; 
        10'b0010110101: data <= 12'h00b; 
        10'b0010110110: data <= 12'h010; 
        10'b0010110111: data <= 12'h00d; 
        10'b0010111000: data <= 12'h009; 
        10'b0010111001: data <= 12'h007; 
        10'b0010111010: data <= 12'h009; 
        10'b0010111011: data <= 12'hffe; 
        10'b0010111100: data <= 12'hffe; 
        10'b0010111101: data <= 12'hff9; 
        10'b0010111110: data <= 12'hff3; 
        10'b0010111111: data <= 12'hff4; 
        10'b0011000000: data <= 12'hff9; 
        10'b0011000001: data <= 12'hffd; 
        10'b0011000010: data <= 12'hfff; 
        10'b0011000011: data <= 12'h001; 
        10'b0011000100: data <= 12'h003; 
        10'b0011000101: data <= 12'h000; 
        10'b0011000110: data <= 12'hfff; 
        10'b0011000111: data <= 12'hfff; 
        10'b0011001000: data <= 12'hff9; 
        10'b0011001001: data <= 12'hff5; 
        10'b0011001010: data <= 12'hff4; 
        10'b0011001011: data <= 12'hff1; 
        10'b0011001100: data <= 12'hff2; 
        10'b0011001101: data <= 12'hffb; 
        10'b0011001110: data <= 12'h000; 
        10'b0011001111: data <= 12'h004; 
        10'b0011010000: data <= 12'h00f; 
        10'b0011010001: data <= 12'h012; 
        10'b0011010010: data <= 12'h018; 
        10'b0011010011: data <= 12'h018; 
        10'b0011010100: data <= 12'h019; 
        10'b0011010101: data <= 12'h00b; 
        10'b0011010110: data <= 12'h009; 
        10'b0011010111: data <= 12'h001; 
        10'b0011011000: data <= 12'h002; 
        10'b0011011001: data <= 12'h003; 
        10'b0011011010: data <= 12'hff7; 
        10'b0011011011: data <= 12'hff1; 
        10'b0011011100: data <= 12'hff7; 
        10'b0011011101: data <= 12'hffe; 
        10'b0011011110: data <= 12'hffe; 
        10'b0011011111: data <= 12'h002; 
        10'b0011100000: data <= 12'h003; 
        10'b0011100001: data <= 12'h003; 
        10'b0011100010: data <= 12'h002; 
        10'b0011100011: data <= 12'hfff; 
        10'b0011100100: data <= 12'hff9; 
        10'b0011100101: data <= 12'hff5; 
        10'b0011100110: data <= 12'hff3; 
        10'b0011100111: data <= 12'hfee; 
        10'b0011101000: data <= 12'hffb; 
        10'b0011101001: data <= 12'hffe; 
        10'b0011101010: data <= 12'hffd; 
        10'b0011101011: data <= 12'hffb; 
        10'b0011101100: data <= 12'h000; 
        10'b0011101101: data <= 12'h007; 
        10'b0011101110: data <= 12'h015; 
        10'b0011101111: data <= 12'h00b; 
        10'b0011110000: data <= 12'h00c; 
        10'b0011110001: data <= 12'h002; 
        10'b0011110010: data <= 12'h001; 
        10'b0011110011: data <= 12'h001; 
        10'b0011110100: data <= 12'hffc; 
        10'b0011110101: data <= 12'h002; 
        10'b0011110110: data <= 12'hffb; 
        10'b0011110111: data <= 12'hff4; 
        10'b0011111000: data <= 12'hff6; 
        10'b0011111001: data <= 12'hffb; 
        10'b0011111010: data <= 12'hffe; 
        10'b0011111011: data <= 12'h003; 
        10'b0011111100: data <= 12'h001; 
        10'b0011111101: data <= 12'h001; 
        10'b0011111110: data <= 12'h000; 
        10'b0011111111: data <= 12'hffb; 
        10'b0100000000: data <= 12'hff5; 
        10'b0100000001: data <= 12'hff7; 
        10'b0100000010: data <= 12'hffe; 
        10'b0100000011: data <= 12'hffb; 
        10'b0100000100: data <= 12'hffd; 
        10'b0100000101: data <= 12'hfff; 
        10'b0100000110: data <= 12'h005; 
        10'b0100000111: data <= 12'h003; 
        10'b0100001000: data <= 12'h001; 
        10'b0100001001: data <= 12'h008; 
        10'b0100001010: data <= 12'h00e; 
        10'b0100001011: data <= 12'h00d; 
        10'b0100001100: data <= 12'h000; 
        10'b0100001101: data <= 12'hffc; 
        10'b0100001110: data <= 12'h000; 
        10'b0100001111: data <= 12'hff8; 
        10'b0100010000: data <= 12'hffd; 
        10'b0100010001: data <= 12'hff8; 
        10'b0100010010: data <= 12'hff7; 
        10'b0100010011: data <= 12'hff7; 
        10'b0100010100: data <= 12'hffa; 
        10'b0100010101: data <= 12'hffd; 
        10'b0100010110: data <= 12'hffe; 
        10'b0100010111: data <= 12'h003; 
        10'b0100011000: data <= 12'h001; 
        10'b0100011001: data <= 12'h000; 
        10'b0100011010: data <= 12'hfff; 
        10'b0100011011: data <= 12'hffe; 
        10'b0100011100: data <= 12'hff7; 
        10'b0100011101: data <= 12'hffb; 
        10'b0100011110: data <= 12'h004; 
        10'b0100011111: data <= 12'h006; 
        10'b0100100000: data <= 12'h00b; 
        10'b0100100001: data <= 12'h00b; 
        10'b0100100010: data <= 12'h00a; 
        10'b0100100011: data <= 12'h00e; 
        10'b0100100100: data <= 12'h007; 
        10'b0100100101: data <= 12'h002; 
        10'b0100100110: data <= 12'h002; 
        10'b0100100111: data <= 12'hff9; 
        10'b0100101000: data <= 12'hffc; 
        10'b0100101001: data <= 12'hfff; 
        10'b0100101010: data <= 12'h005; 
        10'b0100101011: data <= 12'h000; 
        10'b0100101100: data <= 12'h004; 
        10'b0100101101: data <= 12'hffe; 
        10'b0100101110: data <= 12'hffb; 
        10'b0100101111: data <= 12'hffb; 
        10'b0100110000: data <= 12'hffa; 
        10'b0100110001: data <= 12'hffe; 
        10'b0100110010: data <= 12'hffe; 
        10'b0100110011: data <= 12'h001; 
        10'b0100110100: data <= 12'h000; 
        10'b0100110101: data <= 12'h001; 
        10'b0100110110: data <= 12'hfff; 
        10'b0100110111: data <= 12'hfff; 
        10'b0100111000: data <= 12'hffe; 
        10'b0100111001: data <= 12'h008; 
        10'b0100111010: data <= 12'h012; 
        10'b0100111011: data <= 12'h00e; 
        10'b0100111100: data <= 12'h016; 
        10'b0100111101: data <= 12'h009; 
        10'b0100111110: data <= 12'h009; 
        10'b0100111111: data <= 12'h00f; 
        10'b0101000000: data <= 12'hffb; 
        10'b0101000001: data <= 12'hffc; 
        10'b0101000010: data <= 12'hffe; 
        10'b0101000011: data <= 12'h001; 
        10'b0101000100: data <= 12'h006; 
        10'b0101000101: data <= 12'h015; 
        10'b0101000110: data <= 12'h00a; 
        10'b0101000111: data <= 12'h00a; 
        10'b0101001000: data <= 12'h010; 
        10'b0101001001: data <= 12'h00c; 
        10'b0101001010: data <= 12'h007; 
        10'b0101001011: data <= 12'h001; 
        10'b0101001100: data <= 12'hfff; 
        10'b0101001101: data <= 12'hffd; 
        10'b0101001110: data <= 12'h000; 
        10'b0101001111: data <= 12'h000; 
        10'b0101010000: data <= 12'h001; 
        10'b0101010001: data <= 12'h003; 
        10'b0101010010: data <= 12'hffe; 
        10'b0101010011: data <= 12'hffd; 
        10'b0101010100: data <= 12'h007; 
        10'b0101010101: data <= 12'h011; 
        10'b0101010110: data <= 12'h014; 
        10'b0101010111: data <= 12'h00c; 
        10'b0101011000: data <= 12'h00f; 
        10'b0101011001: data <= 12'h012; 
        10'b0101011010: data <= 12'h00c; 
        10'b0101011011: data <= 12'h000; 
        10'b0101011100: data <= 12'hff4; 
        10'b0101011101: data <= 12'h00a; 
        10'b0101011110: data <= 12'h016; 
        10'b0101011111: data <= 12'h011; 
        10'b0101100000: data <= 12'h00f; 
        10'b0101100001: data <= 12'h017; 
        10'b0101100010: data <= 12'h017; 
        10'b0101100011: data <= 12'h018; 
        10'b0101100100: data <= 12'h018; 
        10'b0101100101: data <= 12'h010; 
        10'b0101100110: data <= 12'h008; 
        10'b0101100111: data <= 12'h000; 
        10'b0101101000: data <= 12'hffc; 
        10'b0101101001: data <= 12'h001; 
        10'b0101101010: data <= 12'h001; 
        10'b0101101011: data <= 12'h001; 
        10'b0101101100: data <= 12'h003; 
        10'b0101101101: data <= 12'h002; 
        10'b0101101110: data <= 12'hffd; 
        10'b0101101111: data <= 12'h001; 
        10'b0101110000: data <= 12'h00a; 
        10'b0101110001: data <= 12'h00f; 
        10'b0101110010: data <= 12'h00e; 
        10'b0101110011: data <= 12'h009; 
        10'b0101110100: data <= 12'h00c; 
        10'b0101110101: data <= 12'h008; 
        10'b0101110110: data <= 12'h007; 
        10'b0101110111: data <= 12'hffc; 
        10'b0101111000: data <= 12'hffa; 
        10'b0101111001: data <= 12'h010; 
        10'b0101111010: data <= 12'h016; 
        10'b0101111011: data <= 12'h010; 
        10'b0101111100: data <= 12'h012; 
        10'b0101111101: data <= 12'h010; 
        10'b0101111110: data <= 12'h016; 
        10'b0101111111: data <= 12'h017; 
        10'b0110000000: data <= 12'h012; 
        10'b0110000001: data <= 12'h00a; 
        10'b0110000010: data <= 12'h001; 
        10'b0110000011: data <= 12'hff9; 
        10'b0110000100: data <= 12'hffc; 
        10'b0110000101: data <= 12'hfff; 
        10'b0110000110: data <= 12'h001; 
        10'b0110000111: data <= 12'h001; 
        10'b0110001000: data <= 12'h001; 
        10'b0110001001: data <= 12'h000; 
        10'b0110001010: data <= 12'h002; 
        10'b0110001011: data <= 12'h001; 
        10'b0110001100: data <= 12'h005; 
        10'b0110001101: data <= 12'h004; 
        10'b0110001110: data <= 12'h00c; 
        10'b0110001111: data <= 12'h008; 
        10'b0110010000: data <= 12'h004; 
        10'b0110010001: data <= 12'h000; 
        10'b0110010010: data <= 12'h001; 
        10'b0110010011: data <= 12'hfff; 
        10'b0110010100: data <= 12'hffc; 
        10'b0110010101: data <= 12'h005; 
        10'b0110010110: data <= 12'h003; 
        10'b0110010111: data <= 12'h00e; 
        10'b0110011000: data <= 12'h00f; 
        10'b0110011001: data <= 12'h00f; 
        10'b0110011010: data <= 12'h00a; 
        10'b0110011011: data <= 12'h007; 
        10'b0110011100: data <= 12'h008; 
        10'b0110011101: data <= 12'h000; 
        10'b0110011110: data <= 12'hff8; 
        10'b0110011111: data <= 12'hff4; 
        10'b0110100000: data <= 12'hffb; 
        10'b0110100001: data <= 12'h001; 
        10'b0110100010: data <= 12'h000; 
        10'b0110100011: data <= 12'h001; 
        10'b0110100100: data <= 12'h002; 
        10'b0110100101: data <= 12'h002; 
        10'b0110100110: data <= 12'h001; 
        10'b0110100111: data <= 12'hffe; 
        10'b0110101000: data <= 12'h000; 
        10'b0110101001: data <= 12'h005; 
        10'b0110101010: data <= 12'h005; 
        10'b0110101011: data <= 12'h003; 
        10'b0110101100: data <= 12'h003; 
        10'b0110101101: data <= 12'hffa; 
        10'b0110101110: data <= 12'hffd; 
        10'b0110101111: data <= 12'hffd; 
        10'b0110110000: data <= 12'hffc; 
        10'b0110110001: data <= 12'hffd; 
        10'b0110110010: data <= 12'hffc; 
        10'b0110110011: data <= 12'h00f; 
        10'b0110110100: data <= 12'h016; 
        10'b0110110101: data <= 12'h015; 
        10'b0110110110: data <= 12'h00b; 
        10'b0110110111: data <= 12'h001; 
        10'b0110111000: data <= 12'hffb; 
        10'b0110111001: data <= 12'hff4; 
        10'b0110111010: data <= 12'hff1; 
        10'b0110111011: data <= 12'hff5; 
        10'b0110111100: data <= 12'hffb; 
        10'b0110111101: data <= 12'h000; 
        10'b0110111110: data <= 12'h001; 
        10'b0110111111: data <= 12'h000; 
        10'b0111000000: data <= 12'h003; 
        10'b0111000001: data <= 12'h000; 
        10'b0111000010: data <= 12'hffe; 
        10'b0111000011: data <= 12'h000; 
        10'b0111000100: data <= 12'h000; 
        10'b0111000101: data <= 12'h002; 
        10'b0111000110: data <= 12'hffc; 
        10'b0111000111: data <= 12'h003; 
        10'b0111001000: data <= 12'h009; 
        10'b0111001001: data <= 12'hffe; 
        10'b0111001010: data <= 12'h005; 
        10'b0111001011: data <= 12'h007; 
        10'b0111001100: data <= 12'hfff; 
        10'b0111001101: data <= 12'hff8; 
        10'b0111001110: data <= 12'hfff; 
        10'b0111001111: data <= 12'h008; 
        10'b0111010000: data <= 12'h00f; 
        10'b0111010001: data <= 12'h00f; 
        10'b0111010010: data <= 12'h004; 
        10'b0111010011: data <= 12'hff7; 
        10'b0111010100: data <= 12'hff2; 
        10'b0111010101: data <= 12'hfec; 
        10'b0111010110: data <= 12'hff2; 
        10'b0111010111: data <= 12'hff5; 
        10'b0111011000: data <= 12'hff9; 
        10'b0111011001: data <= 12'h000; 
        10'b0111011010: data <= 12'hffe; 
        10'b0111011011: data <= 12'h001; 
        10'b0111011100: data <= 12'h001; 
        10'b0111011101: data <= 12'hfff; 
        10'b0111011110: data <= 12'hffe; 
        10'b0111011111: data <= 12'hffd; 
        10'b0111100000: data <= 12'hffa; 
        10'b0111100001: data <= 12'hff9; 
        10'b0111100010: data <= 12'hffa; 
        10'b0111100011: data <= 12'h003; 
        10'b0111100100: data <= 12'h005; 
        10'b0111100101: data <= 12'h006; 
        10'b0111100110: data <= 12'h009; 
        10'b0111100111: data <= 12'h00d; 
        10'b0111101000: data <= 12'h008; 
        10'b0111101001: data <= 12'h004; 
        10'b0111101010: data <= 12'h005; 
        10'b0111101011: data <= 12'h00c; 
        10'b0111101100: data <= 12'h004; 
        10'b0111101101: data <= 12'hffd; 
        10'b0111101110: data <= 12'hffa; 
        10'b0111101111: data <= 12'hff3; 
        10'b0111110000: data <= 12'hff4; 
        10'b0111110001: data <= 12'hff3; 
        10'b0111110010: data <= 12'hff3; 
        10'b0111110011: data <= 12'hff7; 
        10'b0111110100: data <= 12'hff9; 
        10'b0111110101: data <= 12'h001; 
        10'b0111110110: data <= 12'h001; 
        10'b0111110111: data <= 12'hfff; 
        10'b0111111000: data <= 12'h002; 
        10'b0111111001: data <= 12'h000; 
        10'b0111111010: data <= 12'hfff; 
        10'b0111111011: data <= 12'hfff; 
        10'b0111111100: data <= 12'hffb; 
        10'b0111111101: data <= 12'hff5; 
        10'b0111111110: data <= 12'hff4; 
        10'b0111111111: data <= 12'hff5; 
        10'b1000000000: data <= 12'hffb; 
        10'b1000000001: data <= 12'h002; 
        10'b1000000010: data <= 12'h00e; 
        10'b1000000011: data <= 12'h00b; 
        10'b1000000100: data <= 12'hff9; 
        10'b1000000101: data <= 12'hff9; 
        10'b1000000110: data <= 12'h000; 
        10'b1000000111: data <= 12'h008; 
        10'b1000001000: data <= 12'hffb; 
        10'b1000001001: data <= 12'hffa; 
        10'b1000001010: data <= 12'hff5; 
        10'b1000001011: data <= 12'hffa; 
        10'b1000001100: data <= 12'hffa; 
        10'b1000001101: data <= 12'hff6; 
        10'b1000001110: data <= 12'hff6; 
        10'b1000001111: data <= 12'hff6; 
        10'b1000010000: data <= 12'hff9; 
        10'b1000010001: data <= 12'hfff; 
        10'b1000010010: data <= 12'h000; 
        10'b1000010011: data <= 12'h002; 
        10'b1000010100: data <= 12'h002; 
        10'b1000010101: data <= 12'h003; 
        10'b1000010110: data <= 12'h001; 
        10'b1000010111: data <= 12'hffd; 
        10'b1000011000: data <= 12'hffb; 
        10'b1000011001: data <= 12'hff8; 
        10'b1000011010: data <= 12'hff3; 
        10'b1000011011: data <= 12'hff3; 
        10'b1000011100: data <= 12'hff2; 
        10'b1000011101: data <= 12'hff3; 
        10'b1000011110: data <= 12'hff1; 
        10'b1000011111: data <= 12'hff3; 
        10'b1000100000: data <= 12'hff0; 
        10'b1000100001: data <= 12'hff5; 
        10'b1000100010: data <= 12'hff6; 
        10'b1000100011: data <= 12'hff5; 
        10'b1000100100: data <= 12'hff7; 
        10'b1000100101: data <= 12'hffd; 
        10'b1000100110: data <= 12'hff9; 
        10'b1000100111: data <= 12'hffe; 
        10'b1000101000: data <= 12'hffb; 
        10'b1000101001: data <= 12'hffa; 
        10'b1000101010: data <= 12'hffb; 
        10'b1000101011: data <= 12'hffb; 
        10'b1000101100: data <= 12'hffd; 
        10'b1000101101: data <= 12'h001; 
        10'b1000101110: data <= 12'hfff; 
        10'b1000101111: data <= 12'h000; 
        10'b1000110000: data <= 12'hfff; 
        10'b1000110001: data <= 12'h000; 
        10'b1000110010: data <= 12'h001; 
        10'b1000110011: data <= 12'h000; 
        10'b1000110100: data <= 12'hffb; 
        10'b1000110101: data <= 12'hff8; 
        10'b1000110110: data <= 12'hff4; 
        10'b1000110111: data <= 12'hfee; 
        10'b1000111000: data <= 12'hfeb; 
        10'b1000111001: data <= 12'hfe8; 
        10'b1000111010: data <= 12'hfe0; 
        10'b1000111011: data <= 12'hfe7; 
        10'b1000111100: data <= 12'hfe8; 
        10'b1000111101: data <= 12'hff8; 
        10'b1000111110: data <= 12'hff5; 
        10'b1000111111: data <= 12'hffb; 
        10'b1001000000: data <= 12'hffa; 
        10'b1001000001: data <= 12'hffe; 
        10'b1001000010: data <= 12'hff5; 
        10'b1001000011: data <= 12'hffd; 
        10'b1001000100: data <= 12'hffc; 
        10'b1001000101: data <= 12'hff9; 
        10'b1001000110: data <= 12'hffe; 
        10'b1001000111: data <= 12'hffd; 
        10'b1001001000: data <= 12'h000; 
        10'b1001001001: data <= 12'h003; 
        10'b1001001010: data <= 12'h002; 
        10'b1001001011: data <= 12'h001; 
        10'b1001001100: data <= 12'h000; 
        10'b1001001101: data <= 12'h000; 
        10'b1001001110: data <= 12'h003; 
        10'b1001001111: data <= 12'hffd; 
        10'b1001010000: data <= 12'hffd; 
        10'b1001010001: data <= 12'hff8; 
        10'b1001010010: data <= 12'hff5; 
        10'b1001010011: data <= 12'hfef; 
        10'b1001010100: data <= 12'hfed; 
        10'b1001010101: data <= 12'hfeb; 
        10'b1001010110: data <= 12'hfea; 
        10'b1001010111: data <= 12'hfec; 
        10'b1001011000: data <= 12'hff3; 
        10'b1001011001: data <= 12'hff4; 
        10'b1001011010: data <= 12'hff3; 
        10'b1001011011: data <= 12'hff9; 
        10'b1001011100: data <= 12'hff8; 
        10'b1001011101: data <= 12'hff4; 
        10'b1001011110: data <= 12'hff2; 
        10'b1001011111: data <= 12'hffa; 
        10'b1001100000: data <= 12'hffd; 
        10'b1001100001: data <= 12'hffe; 
        10'b1001100010: data <= 12'h001; 
        10'b1001100011: data <= 12'h000; 
        10'b1001100100: data <= 12'h001; 
        10'b1001100101: data <= 12'h002; 
        10'b1001100110: data <= 12'h000; 
        10'b1001100111: data <= 12'h000; 
        10'b1001101000: data <= 12'h002; 
        10'b1001101001: data <= 12'h001; 
        10'b1001101010: data <= 12'h001; 
        10'b1001101011: data <= 12'h002; 
        10'b1001101100: data <= 12'hfff; 
        10'b1001101101: data <= 12'hffa; 
        10'b1001101110: data <= 12'hff6; 
        10'b1001101111: data <= 12'hff3; 
        10'b1001110000: data <= 12'hff6; 
        10'b1001110001: data <= 12'hff6; 
        10'b1001110010: data <= 12'hff5; 
        10'b1001110011: data <= 12'hff8; 
        10'b1001110100: data <= 12'hff7; 
        10'b1001110101: data <= 12'hff4; 
        10'b1001110110: data <= 12'hff6; 
        10'b1001110111: data <= 12'hff2; 
        10'b1001111000: data <= 12'hff1; 
        10'b1001111001: data <= 12'hff1; 
        10'b1001111010: data <= 12'hff4; 
        10'b1001111011: data <= 12'hff5; 
        10'b1001111100: data <= 12'hffd; 
        10'b1001111101: data <= 12'h004; 
        10'b1001111110: data <= 12'h002; 
        10'b1001111111: data <= 12'h003; 
        10'b1010000000: data <= 12'h004; 
        10'b1010000001: data <= 12'h001; 
        10'b1010000010: data <= 12'h001; 
        10'b1010000011: data <= 12'h002; 
        10'b1010000100: data <= 12'h002; 
        10'b1010000101: data <= 12'h002; 
        10'b1010000110: data <= 12'h001; 
        10'b1010000111: data <= 12'hfff; 
        10'b1010001000: data <= 12'hffe; 
        10'b1010001001: data <= 12'hffb; 
        10'b1010001010: data <= 12'hffa; 
        10'b1010001011: data <= 12'hff8; 
        10'b1010001100: data <= 12'hfff; 
        10'b1010001101: data <= 12'hffd; 
        10'b1010001110: data <= 12'hffd; 
        10'b1010001111: data <= 12'hff6; 
        10'b1010010000: data <= 12'hff8; 
        10'b1010010001: data <= 12'hff6; 
        10'b1010010010: data <= 12'hff7; 
        10'b1010010011: data <= 12'hff1; 
        10'b1010010100: data <= 12'hff0; 
        10'b1010010101: data <= 12'hff2; 
        10'b1010010110: data <= 12'hff7; 
        10'b1010010111: data <= 12'hfff; 
        10'b1010011000: data <= 12'h003; 
        10'b1010011001: data <= 12'h008; 
        10'b1010011010: data <= 12'h00b; 
        10'b1010011011: data <= 12'h00a; 
        10'b1010011100: data <= 12'h004; 
        10'b1010011101: data <= 12'h000; 
        10'b1010011110: data <= 12'h003; 
        10'b1010011111: data <= 12'h000; 
        10'b1010100000: data <= 12'h000; 
        10'b1010100001: data <= 12'hfff; 
        10'b1010100010: data <= 12'h000; 
        10'b1010100011: data <= 12'h003; 
        10'b1010100100: data <= 12'h002; 
        10'b1010100101: data <= 12'h003; 
        10'b1010100110: data <= 12'h002; 
        10'b1010100111: data <= 12'h003; 
        10'b1010101000: data <= 12'h005; 
        10'b1010101001: data <= 12'h002; 
        10'b1010101010: data <= 12'hffe; 
        10'b1010101011: data <= 12'hffb; 
        10'b1010101100: data <= 12'h000; 
        10'b1010101101: data <= 12'hff8; 
        10'b1010101110: data <= 12'hff6; 
        10'b1010101111: data <= 12'hff6; 
        10'b1010110000: data <= 12'hffb; 
        10'b1010110001: data <= 12'h003; 
        10'b1010110010: data <= 12'h006; 
        10'b1010110011: data <= 12'h006; 
        10'b1010110100: data <= 12'h00e; 
        10'b1010110101: data <= 12'h00f; 
        10'b1010110110: data <= 12'h009; 
        10'b1010110111: data <= 12'h005; 
        10'b1010111000: data <= 12'h004; 
        10'b1010111001: data <= 12'hfff; 
        10'b1010111010: data <= 12'h002; 
        10'b1010111011: data <= 12'h000; 
        10'b1010111100: data <= 12'h001; 
        10'b1010111101: data <= 12'h003; 
        10'b1010111110: data <= 12'h003; 
        10'b1010111111: data <= 12'h000; 
        10'b1011000000: data <= 12'h000; 
        10'b1011000001: data <= 12'h005; 
        10'b1011000010: data <= 12'h003; 
        10'b1011000011: data <= 12'h00a; 
        10'b1011000100: data <= 12'h00b; 
        10'b1011000101: data <= 12'h00b; 
        10'b1011000110: data <= 12'h00a; 
        10'b1011000111: data <= 12'h004; 
        10'b1011001000: data <= 12'h00a; 
        10'b1011001001: data <= 12'h009; 
        10'b1011001010: data <= 12'h009; 
        10'b1011001011: data <= 12'h008; 
        10'b1011001100: data <= 12'h00f; 
        10'b1011001101: data <= 12'h011; 
        10'b1011001110: data <= 12'h012; 
        10'b1011001111: data <= 12'h013; 
        10'b1011010000: data <= 12'h015; 
        10'b1011010001: data <= 12'h00f; 
        10'b1011010010: data <= 12'h006; 
        10'b1011010011: data <= 12'h003; 
        10'b1011010100: data <= 12'h000; 
        10'b1011010101: data <= 12'h000; 
        10'b1011010110: data <= 12'h001; 
        10'b1011010111: data <= 12'h001; 
        10'b1011011000: data <= 12'h000; 
        10'b1011011001: data <= 12'h002; 
        10'b1011011010: data <= 12'h001; 
        10'b1011011011: data <= 12'hfff; 
        10'b1011011100: data <= 12'h002; 
        10'b1011011101: data <= 12'h004; 
        10'b1011011110: data <= 12'h005; 
        10'b1011011111: data <= 12'h007; 
        10'b1011100000: data <= 12'h008; 
        10'b1011100001: data <= 12'h00d; 
        10'b1011100010: data <= 12'h00d; 
        10'b1011100011: data <= 12'h00f; 
        10'b1011100100: data <= 12'h012; 
        10'b1011100101: data <= 12'h012; 
        10'b1011100110: data <= 12'h016; 
        10'b1011100111: data <= 12'h00d; 
        10'b1011101000: data <= 12'h009; 
        10'b1011101001: data <= 12'h007; 
        10'b1011101010: data <= 12'h00b; 
        10'b1011101011: data <= 12'h00c; 
        10'b1011101100: data <= 12'h008; 
        10'b1011101101: data <= 12'h006; 
        10'b1011101110: data <= 12'h002; 
        10'b1011101111: data <= 12'h001; 
        10'b1011110000: data <= 12'h001; 
        10'b1011110001: data <= 12'h001; 
        10'b1011110010: data <= 12'hfff; 
        10'b1011110011: data <= 12'h001; 
        10'b1011110100: data <= 12'hfff; 
        10'b1011110101: data <= 12'h001; 
        10'b1011110110: data <= 12'hfff; 
        10'b1011110111: data <= 12'h003; 
        10'b1011111000: data <= 12'h002; 
        10'b1011111001: data <= 12'h001; 
        10'b1011111010: data <= 12'h000; 
        10'b1011111011: data <= 12'h003; 
        10'b1011111100: data <= 12'h002; 
        10'b1011111101: data <= 12'h002; 
        10'b1011111110: data <= 12'hfff; 
        10'b1011111111: data <= 12'hfff; 
        10'b1100000000: data <= 12'h001; 
        10'b1100000001: data <= 12'hfff; 
        10'b1100000010: data <= 12'h001; 
        10'b1100000011: data <= 12'h002; 
        10'b1100000100: data <= 12'h000; 
        10'b1100000101: data <= 12'h001; 
        10'b1100000110: data <= 12'h003; 
        10'b1100000111: data <= 12'h003; 
        10'b1100001000: data <= 12'h002; 
        10'b1100001001: data <= 12'h001; 
        10'b1100001010: data <= 12'hfff; 
        10'b1100001011: data <= 12'h003; 
        10'b1100001100: data <= 12'h002; 
        10'b1100001101: data <= 12'hfff; 
        10'b1100001110: data <= 12'h000; 
        10'b1100001111: data <= 12'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 7) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 13'h0005; 
        10'b0000000001: data <= 13'h0004; 
        10'b0000000010: data <= 13'h1fff; 
        10'b0000000011: data <= 13'h0003; 
        10'b0000000100: data <= 13'h0003; 
        10'b0000000101: data <= 13'h0004; 
        10'b0000000110: data <= 13'h1ffe; 
        10'b0000000111: data <= 13'h0001; 
        10'b0000001000: data <= 13'h0005; 
        10'b0000001001: data <= 13'h1ffe; 
        10'b0000001010: data <= 13'h1fff; 
        10'b0000001011: data <= 13'h0002; 
        10'b0000001100: data <= 13'h0006; 
        10'b0000001101: data <= 13'h0004; 
        10'b0000001110: data <= 13'h1ffe; 
        10'b0000001111: data <= 13'h1fff; 
        10'b0000010000: data <= 13'h1fff; 
        10'b0000010001: data <= 13'h0002; 
        10'b0000010010: data <= 13'h0004; 
        10'b0000010011: data <= 13'h0000; 
        10'b0000010100: data <= 13'h0000; 
        10'b0000010101: data <= 13'h0000; 
        10'b0000010110: data <= 13'h1ffe; 
        10'b0000010111: data <= 13'h0001; 
        10'b0000011000: data <= 13'h0005; 
        10'b0000011001: data <= 13'h0001; 
        10'b0000011010: data <= 13'h1ffe; 
        10'b0000011011: data <= 13'h0002; 
        10'b0000011100: data <= 13'h0004; 
        10'b0000011101: data <= 13'h0003; 
        10'b0000011110: data <= 13'h0002; 
        10'b0000011111: data <= 13'h1fff; 
        10'b0000100000: data <= 13'h1ffe; 
        10'b0000100001: data <= 13'h1ffe; 
        10'b0000100010: data <= 13'h0000; 
        10'b0000100011: data <= 13'h0006; 
        10'b0000100100: data <= 13'h1ffe; 
        10'b0000100101: data <= 13'h0005; 
        10'b0000100110: data <= 13'h0002; 
        10'b0000100111: data <= 13'h0003; 
        10'b0000101000: data <= 13'h0002; 
        10'b0000101001: data <= 13'h0003; 
        10'b0000101010: data <= 13'h0000; 
        10'b0000101011: data <= 13'h1ffd; 
        10'b0000101100: data <= 13'h1fff; 
        10'b0000101101: data <= 13'h0004; 
        10'b0000101110: data <= 13'h0000; 
        10'b0000101111: data <= 13'h0001; 
        10'b0000110000: data <= 13'h0005; 
        10'b0000110001: data <= 13'h0000; 
        10'b0000110010: data <= 13'h0001; 
        10'b0000110011: data <= 13'h0000; 
        10'b0000110100: data <= 13'h0003; 
        10'b0000110101: data <= 13'h0005; 
        10'b0000110110: data <= 13'h0000; 
        10'b0000110111: data <= 13'h0001; 
        10'b0000111000: data <= 13'h0005; 
        10'b0000111001: data <= 13'h0005; 
        10'b0000111010: data <= 13'h0000; 
        10'b0000111011: data <= 13'h0004; 
        10'b0000111100: data <= 13'h0005; 
        10'b0000111101: data <= 13'h0000; 
        10'b0000111110: data <= 13'h1fff; 
        10'b0000111111: data <= 13'h0002; 
        10'b0001000000: data <= 13'h0005; 
        10'b0001000001: data <= 13'h1fff; 
        10'b0001000010: data <= 13'h1fff; 
        10'b0001000011: data <= 13'h0003; 
        10'b0001000100: data <= 13'h0002; 
        10'b0001000101: data <= 13'h0004; 
        10'b0001000110: data <= 13'h1ffd; 
        10'b0001000111: data <= 13'h0005; 
        10'b0001001000: data <= 13'h1ffe; 
        10'b0001001001: data <= 13'h1ffe; 
        10'b0001001010: data <= 13'h0000; 
        10'b0001001011: data <= 13'h1ffe; 
        10'b0001001100: data <= 13'h0005; 
        10'b0001001101: data <= 13'h1fff; 
        10'b0001001110: data <= 13'h1ffe; 
        10'b0001001111: data <= 13'h0005; 
        10'b0001010000: data <= 13'h0001; 
        10'b0001010001: data <= 13'h0001; 
        10'b0001010010: data <= 13'h0001; 
        10'b0001010011: data <= 13'h0002; 
        10'b0001010100: data <= 13'h0007; 
        10'b0001010101: data <= 13'h0000; 
        10'b0001010110: data <= 13'h1fff; 
        10'b0001010111: data <= 13'h0002; 
        10'b0001011000: data <= 13'h0002; 
        10'b0001011001: data <= 13'h1ffe; 
        10'b0001011010: data <= 13'h0005; 
        10'b0001011011: data <= 13'h0003; 
        10'b0001011100: data <= 13'h1fff; 
        10'b0001011101: data <= 13'h0005; 
        10'b0001011110: data <= 13'h0002; 
        10'b0001011111: data <= 13'h0004; 
        10'b0001100000: data <= 13'h0000; 
        10'b0001100001: data <= 13'h1ffb; 
        10'b0001100010: data <= 13'h0000; 
        10'b0001100011: data <= 13'h1ff9; 
        10'b0001100100: data <= 13'h1fff; 
        10'b0001100101: data <= 13'h1ffc; 
        10'b0001100110: data <= 13'h0001; 
        10'b0001100111: data <= 13'h0001; 
        10'b0001101000: data <= 13'h0002; 
        10'b0001101001: data <= 13'h0000; 
        10'b0001101010: data <= 13'h0004; 
        10'b0001101011: data <= 13'h1fff; 
        10'b0001101100: data <= 13'h1fff; 
        10'b0001101101: data <= 13'h0006; 
        10'b0001101110: data <= 13'h0002; 
        10'b0001101111: data <= 13'h0004; 
        10'b0001110000: data <= 13'h0001; 
        10'b0001110001: data <= 13'h0001; 
        10'b0001110010: data <= 13'h0000; 
        10'b0001110011: data <= 13'h1fff; 
        10'b0001110100: data <= 13'h1ffe; 
        10'b0001110101: data <= 13'h0004; 
        10'b0001110110: data <= 13'h0003; 
        10'b0001110111: data <= 13'h0000; 
        10'b0001111000: data <= 13'h1ffd; 
        10'b0001111001: data <= 13'h0001; 
        10'b0001111010: data <= 13'h1ffb; 
        10'b0001111011: data <= 13'h1ff8; 
        10'b0001111100: data <= 13'h1ff5; 
        10'b0001111101: data <= 13'h1fec; 
        10'b0001111110: data <= 13'h1fe7; 
        10'b0001111111: data <= 13'h1fdf; 
        10'b0010000000: data <= 13'h1fe7; 
        10'b0010000001: data <= 13'h1fe7; 
        10'b0010000010: data <= 13'h1fee; 
        10'b0010000011: data <= 13'h1ff8; 
        10'b0010000100: data <= 13'h1ffc; 
        10'b0010000101: data <= 13'h1ffd; 
        10'b0010000110: data <= 13'h0001; 
        10'b0010000111: data <= 13'h0005; 
        10'b0010001000: data <= 13'h0004; 
        10'b0010001001: data <= 13'h0003; 
        10'b0010001010: data <= 13'h0000; 
        10'b0010001011: data <= 13'h0000; 
        10'b0010001100: data <= 13'h0005; 
        10'b0010001101: data <= 13'h0003; 
        10'b0010001110: data <= 13'h0004; 
        10'b0010001111: data <= 13'h0002; 
        10'b0010010000: data <= 13'h0003; 
        10'b0010010001: data <= 13'h1ffc; 
        10'b0010010010: data <= 13'h1ffd; 
        10'b0010010011: data <= 13'h1ffc; 
        10'b0010010100: data <= 13'h1ff5; 
        10'b0010010101: data <= 13'h1ff5; 
        10'b0010010110: data <= 13'h1ff4; 
        10'b0010010111: data <= 13'h1ff0; 
        10'b0010011000: data <= 13'h1fec; 
        10'b0010011001: data <= 13'h1fe9; 
        10'b0010011010: data <= 13'h1fdc; 
        10'b0010011011: data <= 13'h1fd9; 
        10'b0010011100: data <= 13'h1fcf; 
        10'b0010011101: data <= 13'h1fe0; 
        10'b0010011110: data <= 13'h1fec; 
        10'b0010011111: data <= 13'h1ff6; 
        10'b0010100000: data <= 13'h1ff6; 
        10'b0010100001: data <= 13'h1ff2; 
        10'b0010100010: data <= 13'h1ff3; 
        10'b0010100011: data <= 13'h1ff7; 
        10'b0010100100: data <= 13'h1ffc; 
        10'b0010100101: data <= 13'h1ffe; 
        10'b0010100110: data <= 13'h0001; 
        10'b0010100111: data <= 13'h0003; 
        10'b0010101000: data <= 13'h0004; 
        10'b0010101001: data <= 13'h0004; 
        10'b0010101010: data <= 13'h1ffd; 
        10'b0010101011: data <= 13'h0004; 
        10'b0010101100: data <= 13'h0003; 
        10'b0010101101: data <= 13'h1ff4; 
        10'b0010101110: data <= 13'h1ff1; 
        10'b0010101111: data <= 13'h1fef; 
        10'b0010110000: data <= 13'h1fec; 
        10'b0010110001: data <= 13'h1fe8; 
        10'b0010110010: data <= 13'h1fee; 
        10'b0010110011: data <= 13'h1ffa; 
        10'b0010110100: data <= 13'h0001; 
        10'b0010110101: data <= 13'h0016; 
        10'b0010110110: data <= 13'h0020; 
        10'b0010110111: data <= 13'h001a; 
        10'b0010111000: data <= 13'h0012; 
        10'b0010111001: data <= 13'h000f; 
        10'b0010111010: data <= 13'h0013; 
        10'b0010111011: data <= 13'h1ffd; 
        10'b0010111100: data <= 13'h1ffb; 
        10'b0010111101: data <= 13'h1ff2; 
        10'b0010111110: data <= 13'h1fe6; 
        10'b0010111111: data <= 13'h1fe8; 
        10'b0011000000: data <= 13'h1ff2; 
        10'b0011000001: data <= 13'h1ff9; 
        10'b0011000010: data <= 13'h1fff; 
        10'b0011000011: data <= 13'h0002; 
        10'b0011000100: data <= 13'h0006; 
        10'b0011000101: data <= 13'h0000; 
        10'b0011000110: data <= 13'h1ffe; 
        10'b0011000111: data <= 13'h1ffe; 
        10'b0011001000: data <= 13'h1ff2; 
        10'b0011001001: data <= 13'h1feb; 
        10'b0011001010: data <= 13'h1fe7; 
        10'b0011001011: data <= 13'h1fe3; 
        10'b0011001100: data <= 13'h1fe4; 
        10'b0011001101: data <= 13'h1ff6; 
        10'b0011001110: data <= 13'h1fff; 
        10'b0011001111: data <= 13'h0008; 
        10'b0011010000: data <= 13'h001d; 
        10'b0011010001: data <= 13'h0023; 
        10'b0011010010: data <= 13'h0030; 
        10'b0011010011: data <= 13'h0030; 
        10'b0011010100: data <= 13'h0032; 
        10'b0011010101: data <= 13'h0017; 
        10'b0011010110: data <= 13'h0011; 
        10'b0011010111: data <= 13'h0002; 
        10'b0011011000: data <= 13'h0004; 
        10'b0011011001: data <= 13'h0005; 
        10'b0011011010: data <= 13'h1fef; 
        10'b0011011011: data <= 13'h1fe1; 
        10'b0011011100: data <= 13'h1fee; 
        10'b0011011101: data <= 13'h1ffb; 
        10'b0011011110: data <= 13'h1ffb; 
        10'b0011011111: data <= 13'h0004; 
        10'b0011100000: data <= 13'h0006; 
        10'b0011100001: data <= 13'h0006; 
        10'b0011100010: data <= 13'h0003; 
        10'b0011100011: data <= 13'h1ffe; 
        10'b0011100100: data <= 13'h1ff2; 
        10'b0011100101: data <= 13'h1fea; 
        10'b0011100110: data <= 13'h1fe7; 
        10'b0011100111: data <= 13'h1fdd; 
        10'b0011101000: data <= 13'h1ff7; 
        10'b0011101001: data <= 13'h1ffc; 
        10'b0011101010: data <= 13'h1ffb; 
        10'b0011101011: data <= 13'h1ff6; 
        10'b0011101100: data <= 13'h1fff; 
        10'b0011101101: data <= 13'h000e; 
        10'b0011101110: data <= 13'h0029; 
        10'b0011101111: data <= 13'h0017; 
        10'b0011110000: data <= 13'h0017; 
        10'b0011110001: data <= 13'h0005; 
        10'b0011110010: data <= 13'h0002; 
        10'b0011110011: data <= 13'h0001; 
        10'b0011110100: data <= 13'h1ff8; 
        10'b0011110101: data <= 13'h0004; 
        10'b0011110110: data <= 13'h1ff6; 
        10'b0011110111: data <= 13'h1fe7; 
        10'b0011111000: data <= 13'h1feb; 
        10'b0011111001: data <= 13'h1ff6; 
        10'b0011111010: data <= 13'h1ffc; 
        10'b0011111011: data <= 13'h0006; 
        10'b0011111100: data <= 13'h0002; 
        10'b0011111101: data <= 13'h0001; 
        10'b0011111110: data <= 13'h0000; 
        10'b0011111111: data <= 13'h1ff6; 
        10'b0100000000: data <= 13'h1fea; 
        10'b0100000001: data <= 13'h1fef; 
        10'b0100000010: data <= 13'h1ffb; 
        10'b0100000011: data <= 13'h1ff6; 
        10'b0100000100: data <= 13'h1ffa; 
        10'b0100000101: data <= 13'h1ffd; 
        10'b0100000110: data <= 13'h000b; 
        10'b0100000111: data <= 13'h0006; 
        10'b0100001000: data <= 13'h0002; 
        10'b0100001001: data <= 13'h0011; 
        10'b0100001010: data <= 13'h001c; 
        10'b0100001011: data <= 13'h0019; 
        10'b0100001100: data <= 13'h1fff; 
        10'b0100001101: data <= 13'h1ff9; 
        10'b0100001110: data <= 13'h0000; 
        10'b0100001111: data <= 13'h1ff1; 
        10'b0100010000: data <= 13'h1ffa; 
        10'b0100010001: data <= 13'h1ff0; 
        10'b0100010010: data <= 13'h1fef; 
        10'b0100010011: data <= 13'h1fee; 
        10'b0100010100: data <= 13'h1ff4; 
        10'b0100010101: data <= 13'h1ffb; 
        10'b0100010110: data <= 13'h1ffc; 
        10'b0100010111: data <= 13'h0005; 
        10'b0100011000: data <= 13'h0001; 
        10'b0100011001: data <= 13'h0000; 
        10'b0100011010: data <= 13'h1ffe; 
        10'b0100011011: data <= 13'h1ffc; 
        10'b0100011100: data <= 13'h1fef; 
        10'b0100011101: data <= 13'h1ff7; 
        10'b0100011110: data <= 13'h0008; 
        10'b0100011111: data <= 13'h000b; 
        10'b0100100000: data <= 13'h0016; 
        10'b0100100001: data <= 13'h0016; 
        10'b0100100010: data <= 13'h0013; 
        10'b0100100011: data <= 13'h001d; 
        10'b0100100100: data <= 13'h000f; 
        10'b0100100101: data <= 13'h0003; 
        10'b0100100110: data <= 13'h0004; 
        10'b0100100111: data <= 13'h1ff1; 
        10'b0100101000: data <= 13'h1ff7; 
        10'b0100101001: data <= 13'h1ffe; 
        10'b0100101010: data <= 13'h000a; 
        10'b0100101011: data <= 13'h0000; 
        10'b0100101100: data <= 13'h0008; 
        10'b0100101101: data <= 13'h1ffb; 
        10'b0100101110: data <= 13'h1ff6; 
        10'b0100101111: data <= 13'h1ff7; 
        10'b0100110000: data <= 13'h1ff4; 
        10'b0100110001: data <= 13'h1ffd; 
        10'b0100110010: data <= 13'h1ffb; 
        10'b0100110011: data <= 13'h0003; 
        10'b0100110100: data <= 13'h1fff; 
        10'b0100110101: data <= 13'h0001; 
        10'b0100110110: data <= 13'h1ffd; 
        10'b0100110111: data <= 13'h1ffe; 
        10'b0100111000: data <= 13'h1ffb; 
        10'b0100111001: data <= 13'h0010; 
        10'b0100111010: data <= 13'h0025; 
        10'b0100111011: data <= 13'h001b; 
        10'b0100111100: data <= 13'h002b; 
        10'b0100111101: data <= 13'h0011; 
        10'b0100111110: data <= 13'h0012; 
        10'b0100111111: data <= 13'h001f; 
        10'b0101000000: data <= 13'h1ff6; 
        10'b0101000001: data <= 13'h1ff8; 
        10'b0101000010: data <= 13'h1ffb; 
        10'b0101000011: data <= 13'h0002; 
        10'b0101000100: data <= 13'h000c; 
        10'b0101000101: data <= 13'h002a; 
        10'b0101000110: data <= 13'h0014; 
        10'b0101000111: data <= 13'h0014; 
        10'b0101001000: data <= 13'h0021; 
        10'b0101001001: data <= 13'h0018; 
        10'b0101001010: data <= 13'h000e; 
        10'b0101001011: data <= 13'h0003; 
        10'b0101001100: data <= 13'h1ffe; 
        10'b0101001101: data <= 13'h1ffa; 
        10'b0101001110: data <= 13'h0000; 
        10'b0101001111: data <= 13'h0000; 
        10'b0101010000: data <= 13'h0003; 
        10'b0101010001: data <= 13'h0005; 
        10'b0101010010: data <= 13'h1ffc; 
        10'b0101010011: data <= 13'h1ffa; 
        10'b0101010100: data <= 13'h000d; 
        10'b0101010101: data <= 13'h0023; 
        10'b0101010110: data <= 13'h0028; 
        10'b0101010111: data <= 13'h0018; 
        10'b0101011000: data <= 13'h001e; 
        10'b0101011001: data <= 13'h0025; 
        10'b0101011010: data <= 13'h0017; 
        10'b0101011011: data <= 13'h0000; 
        10'b0101011100: data <= 13'h1fe9; 
        10'b0101011101: data <= 13'h0014; 
        10'b0101011110: data <= 13'h002c; 
        10'b0101011111: data <= 13'h0023; 
        10'b0101100000: data <= 13'h001e; 
        10'b0101100001: data <= 13'h002d; 
        10'b0101100010: data <= 13'h002e; 
        10'b0101100011: data <= 13'h002f; 
        10'b0101100100: data <= 13'h0031; 
        10'b0101100101: data <= 13'h0021; 
        10'b0101100110: data <= 13'h0010; 
        10'b0101100111: data <= 13'h0000; 
        10'b0101101000: data <= 13'h1ff9; 
        10'b0101101001: data <= 13'h0001; 
        10'b0101101010: data <= 13'h0003; 
        10'b0101101011: data <= 13'h0003; 
        10'b0101101100: data <= 13'h0006; 
        10'b0101101101: data <= 13'h0004; 
        10'b0101101110: data <= 13'h1ffb; 
        10'b0101101111: data <= 13'h0002; 
        10'b0101110000: data <= 13'h0014; 
        10'b0101110001: data <= 13'h001f; 
        10'b0101110010: data <= 13'h001d; 
        10'b0101110011: data <= 13'h0013; 
        10'b0101110100: data <= 13'h0018; 
        10'b0101110101: data <= 13'h000f; 
        10'b0101110110: data <= 13'h000e; 
        10'b0101110111: data <= 13'h1ff9; 
        10'b0101111000: data <= 13'h1ff4; 
        10'b0101111001: data <= 13'h0020; 
        10'b0101111010: data <= 13'h002c; 
        10'b0101111011: data <= 13'h0020; 
        10'b0101111100: data <= 13'h0025; 
        10'b0101111101: data <= 13'h0021; 
        10'b0101111110: data <= 13'h002d; 
        10'b0101111111: data <= 13'h002e; 
        10'b0110000000: data <= 13'h0024; 
        10'b0110000001: data <= 13'h0015; 
        10'b0110000010: data <= 13'h0001; 
        10'b0110000011: data <= 13'h1ff2; 
        10'b0110000100: data <= 13'h1ff8; 
        10'b0110000101: data <= 13'h1ffd; 
        10'b0110000110: data <= 13'h0003; 
        10'b0110000111: data <= 13'h0003; 
        10'b0110001000: data <= 13'h0001; 
        10'b0110001001: data <= 13'h0001; 
        10'b0110001010: data <= 13'h0004; 
        10'b0110001011: data <= 13'h0003; 
        10'b0110001100: data <= 13'h0009; 
        10'b0110001101: data <= 13'h0009; 
        10'b0110001110: data <= 13'h0018; 
        10'b0110001111: data <= 13'h0011; 
        10'b0110010000: data <= 13'h0008; 
        10'b0110010001: data <= 13'h0000; 
        10'b0110010010: data <= 13'h0003; 
        10'b0110010011: data <= 13'h1fff; 
        10'b0110010100: data <= 13'h1ff7; 
        10'b0110010101: data <= 13'h000a; 
        10'b0110010110: data <= 13'h0006; 
        10'b0110010111: data <= 13'h001c; 
        10'b0110011000: data <= 13'h001e; 
        10'b0110011001: data <= 13'h001e; 
        10'b0110011010: data <= 13'h0014; 
        10'b0110011011: data <= 13'h000d; 
        10'b0110011100: data <= 13'h0010; 
        10'b0110011101: data <= 13'h0000; 
        10'b0110011110: data <= 13'h1ff0; 
        10'b0110011111: data <= 13'h1fe8; 
        10'b0110100000: data <= 13'h1ff6; 
        10'b0110100001: data <= 13'h0002; 
        10'b0110100010: data <= 13'h0001; 
        10'b0110100011: data <= 13'h0001; 
        10'b0110100100: data <= 13'h0005; 
        10'b0110100101: data <= 13'h0004; 
        10'b0110100110: data <= 13'h0003; 
        10'b0110100111: data <= 13'h1ffd; 
        10'b0110101000: data <= 13'h0001; 
        10'b0110101001: data <= 13'h000b; 
        10'b0110101010: data <= 13'h000a; 
        10'b0110101011: data <= 13'h0007; 
        10'b0110101100: data <= 13'h0007; 
        10'b0110101101: data <= 13'h1ff3; 
        10'b0110101110: data <= 13'h1ffa; 
        10'b0110101111: data <= 13'h1ffa; 
        10'b0110110000: data <= 13'h1ff7; 
        10'b0110110001: data <= 13'h1ff9; 
        10'b0110110010: data <= 13'h1ff8; 
        10'b0110110011: data <= 13'h001f; 
        10'b0110110100: data <= 13'h002d; 
        10'b0110110101: data <= 13'h002b; 
        10'b0110110110: data <= 13'h0015; 
        10'b0110110111: data <= 13'h0002; 
        10'b0110111000: data <= 13'h1ff7; 
        10'b0110111001: data <= 13'h1fe7; 
        10'b0110111010: data <= 13'h1fe1; 
        10'b0110111011: data <= 13'h1fea; 
        10'b0110111100: data <= 13'h1ff6; 
        10'b0110111101: data <= 13'h0000; 
        10'b0110111110: data <= 13'h0003; 
        10'b0110111111: data <= 13'h0000; 
        10'b0111000000: data <= 13'h0005; 
        10'b0111000001: data <= 13'h0000; 
        10'b0111000010: data <= 13'h1ffc; 
        10'b0111000011: data <= 13'h1fff; 
        10'b0111000100: data <= 13'h0000; 
        10'b0111000101: data <= 13'h0003; 
        10'b0111000110: data <= 13'h1ff8; 
        10'b0111000111: data <= 13'h0006; 
        10'b0111001000: data <= 13'h0012; 
        10'b0111001001: data <= 13'h1ffc; 
        10'b0111001010: data <= 13'h000a; 
        10'b0111001011: data <= 13'h000f; 
        10'b0111001100: data <= 13'h1ffe; 
        10'b0111001101: data <= 13'h1fef; 
        10'b0111001110: data <= 13'h1ffd; 
        10'b0111001111: data <= 13'h0011; 
        10'b0111010000: data <= 13'h001f; 
        10'b0111010001: data <= 13'h001e; 
        10'b0111010010: data <= 13'h0008; 
        10'b0111010011: data <= 13'h1fef; 
        10'b0111010100: data <= 13'h1fe3; 
        10'b0111010101: data <= 13'h1fd8; 
        10'b0111010110: data <= 13'h1fe4; 
        10'b0111010111: data <= 13'h1fe9; 
        10'b0111011000: data <= 13'h1ff1; 
        10'b0111011001: data <= 13'h0000; 
        10'b0111011010: data <= 13'h1ffd; 
        10'b0111011011: data <= 13'h0003; 
        10'b0111011100: data <= 13'h0002; 
        10'b0111011101: data <= 13'h1fff; 
        10'b0111011110: data <= 13'h1ffc; 
        10'b0111011111: data <= 13'h1ffa; 
        10'b0111100000: data <= 13'h1ff5; 
        10'b0111100001: data <= 13'h1ff2; 
        10'b0111100010: data <= 13'h1ff5; 
        10'b0111100011: data <= 13'h0005; 
        10'b0111100100: data <= 13'h000a; 
        10'b0111100101: data <= 13'h000b; 
        10'b0111100110: data <= 13'h0011; 
        10'b0111100111: data <= 13'h0019; 
        10'b0111101000: data <= 13'h000f; 
        10'b0111101001: data <= 13'h0007; 
        10'b0111101010: data <= 13'h000a; 
        10'b0111101011: data <= 13'h0019; 
        10'b0111101100: data <= 13'h0007; 
        10'b0111101101: data <= 13'h1ffb; 
        10'b0111101110: data <= 13'h1ff5; 
        10'b0111101111: data <= 13'h1fe7; 
        10'b0111110000: data <= 13'h1fe7; 
        10'b0111110001: data <= 13'h1fe5; 
        10'b0111110010: data <= 13'h1fe7; 
        10'b0111110011: data <= 13'h1fed; 
        10'b0111110100: data <= 13'h1ff2; 
        10'b0111110101: data <= 13'h0001; 
        10'b0111110110: data <= 13'h0001; 
        10'b0111110111: data <= 13'h1fff; 
        10'b0111111000: data <= 13'h0005; 
        10'b0111111001: data <= 13'h0000; 
        10'b0111111010: data <= 13'h1ffd; 
        10'b0111111011: data <= 13'h1fff; 
        10'b0111111100: data <= 13'h1ff6; 
        10'b0111111101: data <= 13'h1fe9; 
        10'b0111111110: data <= 13'h1fe9; 
        10'b0111111111: data <= 13'h1fe9; 
        10'b1000000000: data <= 13'h1ff6; 
        10'b1000000001: data <= 13'h0004; 
        10'b1000000010: data <= 13'h001b; 
        10'b1000000011: data <= 13'h0016; 
        10'b1000000100: data <= 13'h1ff2; 
        10'b1000000101: data <= 13'h1ff2; 
        10'b1000000110: data <= 13'h0001; 
        10'b1000000111: data <= 13'h0010; 
        10'b1000001000: data <= 13'h1ff6; 
        10'b1000001001: data <= 13'h1ff4; 
        10'b1000001010: data <= 13'h1fea; 
        10'b1000001011: data <= 13'h1ff3; 
        10'b1000001100: data <= 13'h1ff4; 
        10'b1000001101: data <= 13'h1fed; 
        10'b1000001110: data <= 13'h1fec; 
        10'b1000001111: data <= 13'h1feb; 
        10'b1000010000: data <= 13'h1ff1; 
        10'b1000010001: data <= 13'h1ffe; 
        10'b1000010010: data <= 13'h0000; 
        10'b1000010011: data <= 13'h0004; 
        10'b1000010100: data <= 13'h0003; 
        10'b1000010101: data <= 13'h0006; 
        10'b1000010110: data <= 13'h0001; 
        10'b1000010111: data <= 13'h1ffb; 
        10'b1000011000: data <= 13'h1ff7; 
        10'b1000011001: data <= 13'h1ff0; 
        10'b1000011010: data <= 13'h1fe7; 
        10'b1000011011: data <= 13'h1fe6; 
        10'b1000011100: data <= 13'h1fe5; 
        10'b1000011101: data <= 13'h1fe5; 
        10'b1000011110: data <= 13'h1fe2; 
        10'b1000011111: data <= 13'h1fe7; 
        10'b1000100000: data <= 13'h1fdf; 
        10'b1000100001: data <= 13'h1fe9; 
        10'b1000100010: data <= 13'h1fed; 
        10'b1000100011: data <= 13'h1fea; 
        10'b1000100100: data <= 13'h1fed; 
        10'b1000100101: data <= 13'h1ffa; 
        10'b1000100110: data <= 13'h1ff2; 
        10'b1000100111: data <= 13'h1ffc; 
        10'b1000101000: data <= 13'h1ff6; 
        10'b1000101001: data <= 13'h1ff5; 
        10'b1000101010: data <= 13'h1ff5; 
        10'b1000101011: data <= 13'h1ff6; 
        10'b1000101100: data <= 13'h1ffa; 
        10'b1000101101: data <= 13'h0002; 
        10'b1000101110: data <= 13'h1ffe; 
        10'b1000101111: data <= 13'h0001; 
        10'b1000110000: data <= 13'h1fff; 
        10'b1000110001: data <= 13'h0001; 
        10'b1000110010: data <= 13'h0003; 
        10'b1000110011: data <= 13'h0000; 
        10'b1000110100: data <= 13'h1ff7; 
        10'b1000110101: data <= 13'h1ff0; 
        10'b1000110110: data <= 13'h1fe8; 
        10'b1000110111: data <= 13'h1fdb; 
        10'b1000111000: data <= 13'h1fd6; 
        10'b1000111001: data <= 13'h1fd1; 
        10'b1000111010: data <= 13'h1fc0; 
        10'b1000111011: data <= 13'h1fcf; 
        10'b1000111100: data <= 13'h1fd0; 
        10'b1000111101: data <= 13'h1ff0; 
        10'b1000111110: data <= 13'h1fea; 
        10'b1000111111: data <= 13'h1ff6; 
        10'b1001000000: data <= 13'h1ff4; 
        10'b1001000001: data <= 13'h1ffd; 
        10'b1001000010: data <= 13'h1feb; 
        10'b1001000011: data <= 13'h1ff9; 
        10'b1001000100: data <= 13'h1ff8; 
        10'b1001000101: data <= 13'h1ff3; 
        10'b1001000110: data <= 13'h1ffc; 
        10'b1001000111: data <= 13'h1ffa; 
        10'b1001001000: data <= 13'h0001; 
        10'b1001001001: data <= 13'h0005; 
        10'b1001001010: data <= 13'h0003; 
        10'b1001001011: data <= 13'h0001; 
        10'b1001001100: data <= 13'h0000; 
        10'b1001001101: data <= 13'h0000; 
        10'b1001001110: data <= 13'h0005; 
        10'b1001001111: data <= 13'h1ffa; 
        10'b1001010000: data <= 13'h1ffa; 
        10'b1001010001: data <= 13'h1ff1; 
        10'b1001010010: data <= 13'h1fea; 
        10'b1001010011: data <= 13'h1fdf; 
        10'b1001010100: data <= 13'h1fda; 
        10'b1001010101: data <= 13'h1fd6; 
        10'b1001010110: data <= 13'h1fd4; 
        10'b1001010111: data <= 13'h1fd9; 
        10'b1001011000: data <= 13'h1fe7; 
        10'b1001011001: data <= 13'h1fe7; 
        10'b1001011010: data <= 13'h1fe7; 
        10'b1001011011: data <= 13'h1ff2; 
        10'b1001011100: data <= 13'h1ff0; 
        10'b1001011101: data <= 13'h1fe9; 
        10'b1001011110: data <= 13'h1fe4; 
        10'b1001011111: data <= 13'h1ff4; 
        10'b1001100000: data <= 13'h1ff9; 
        10'b1001100001: data <= 13'h1ffc; 
        10'b1001100010: data <= 13'h0002; 
        10'b1001100011: data <= 13'h1fff; 
        10'b1001100100: data <= 13'h0002; 
        10'b1001100101: data <= 13'h0003; 
        10'b1001100110: data <= 13'h0000; 
        10'b1001100111: data <= 13'h0000; 
        10'b1001101000: data <= 13'h0004; 
        10'b1001101001: data <= 13'h0001; 
        10'b1001101010: data <= 13'h0001; 
        10'b1001101011: data <= 13'h0004; 
        10'b1001101100: data <= 13'h1ffd; 
        10'b1001101101: data <= 13'h1ff4; 
        10'b1001101110: data <= 13'h1fec; 
        10'b1001101111: data <= 13'h1fe5; 
        10'b1001110000: data <= 13'h1fec; 
        10'b1001110001: data <= 13'h1feb; 
        10'b1001110010: data <= 13'h1fe9; 
        10'b1001110011: data <= 13'h1ff1; 
        10'b1001110100: data <= 13'h1fef; 
        10'b1001110101: data <= 13'h1fe9; 
        10'b1001110110: data <= 13'h1fed; 
        10'b1001110111: data <= 13'h1fe5; 
        10'b1001111000: data <= 13'h1fe2; 
        10'b1001111001: data <= 13'h1fe3; 
        10'b1001111010: data <= 13'h1fe7; 
        10'b1001111011: data <= 13'h1fea; 
        10'b1001111100: data <= 13'h1ffa; 
        10'b1001111101: data <= 13'h0007; 
        10'b1001111110: data <= 13'h0004; 
        10'b1001111111: data <= 13'h0005; 
        10'b1010000000: data <= 13'h0008; 
        10'b1010000001: data <= 13'h0002; 
        10'b1010000010: data <= 13'h0002; 
        10'b1010000011: data <= 13'h0003; 
        10'b1010000100: data <= 13'h0005; 
        10'b1010000101: data <= 13'h0004; 
        10'b1010000110: data <= 13'h0001; 
        10'b1010000111: data <= 13'h1ffe; 
        10'b1010001000: data <= 13'h1ffd; 
        10'b1010001001: data <= 13'h1ff5; 
        10'b1010001010: data <= 13'h1ff4; 
        10'b1010001011: data <= 13'h1ff0; 
        10'b1010001100: data <= 13'h1fff; 
        10'b1010001101: data <= 13'h1ff9; 
        10'b1010001110: data <= 13'h1ffb; 
        10'b1010001111: data <= 13'h1fec; 
        10'b1010010000: data <= 13'h1ff0; 
        10'b1010010001: data <= 13'h1fec; 
        10'b1010010010: data <= 13'h1fef; 
        10'b1010010011: data <= 13'h1fe3; 
        10'b1010010100: data <= 13'h1fe0; 
        10'b1010010101: data <= 13'h1fe4; 
        10'b1010010110: data <= 13'h1fef; 
        10'b1010010111: data <= 13'h1ffe; 
        10'b1010011000: data <= 13'h0007; 
        10'b1010011001: data <= 13'h0010; 
        10'b1010011010: data <= 13'h0017; 
        10'b1010011011: data <= 13'h0013; 
        10'b1010011100: data <= 13'h0009; 
        10'b1010011101: data <= 13'h1fff; 
        10'b1010011110: data <= 13'h0006; 
        10'b1010011111: data <= 13'h1fff; 
        10'b1010100000: data <= 13'h0000; 
        10'b1010100001: data <= 13'h1ffd; 
        10'b1010100010: data <= 13'h1fff; 
        10'b1010100011: data <= 13'h0005; 
        10'b1010100100: data <= 13'h0004; 
        10'b1010100101: data <= 13'h0006; 
        10'b1010100110: data <= 13'h0004; 
        10'b1010100111: data <= 13'h0006; 
        10'b1010101000: data <= 13'h0009; 
        10'b1010101001: data <= 13'h0005; 
        10'b1010101010: data <= 13'h1ffd; 
        10'b1010101011: data <= 13'h1ff6; 
        10'b1010101100: data <= 13'h1fff; 
        10'b1010101101: data <= 13'h1ff0; 
        10'b1010101110: data <= 13'h1fec; 
        10'b1010101111: data <= 13'h1feb; 
        10'b1010110000: data <= 13'h1ff7; 
        10'b1010110001: data <= 13'h0007; 
        10'b1010110010: data <= 13'h000c; 
        10'b1010110011: data <= 13'h000c; 
        10'b1010110100: data <= 13'h001c; 
        10'b1010110101: data <= 13'h001e; 
        10'b1010110110: data <= 13'h0011; 
        10'b1010110111: data <= 13'h000a; 
        10'b1010111000: data <= 13'h0008; 
        10'b1010111001: data <= 13'h1ffe; 
        10'b1010111010: data <= 13'h0004; 
        10'b1010111011: data <= 13'h0000; 
        10'b1010111100: data <= 13'h0001; 
        10'b1010111101: data <= 13'h0005; 
        10'b1010111110: data <= 13'h0005; 
        10'b1010111111: data <= 13'h1fff; 
        10'b1011000000: data <= 13'h0001; 
        10'b1011000001: data <= 13'h0009; 
        10'b1011000010: data <= 13'h0007; 
        10'b1011000011: data <= 13'h0014; 
        10'b1011000100: data <= 13'h0016; 
        10'b1011000101: data <= 13'h0016; 
        10'b1011000110: data <= 13'h0013; 
        10'b1011000111: data <= 13'h0008; 
        10'b1011001000: data <= 13'h0014; 
        10'b1011001001: data <= 13'h0012; 
        10'b1011001010: data <= 13'h0011; 
        10'b1011001011: data <= 13'h0010; 
        10'b1011001100: data <= 13'h001f; 
        10'b1011001101: data <= 13'h0021; 
        10'b1011001110: data <= 13'h0024; 
        10'b1011001111: data <= 13'h0026; 
        10'b1011010000: data <= 13'h002a; 
        10'b1011010001: data <= 13'h001e; 
        10'b1011010010: data <= 13'h000c; 
        10'b1011010011: data <= 13'h0006; 
        10'b1011010100: data <= 13'h1fff; 
        10'b1011010101: data <= 13'h0000; 
        10'b1011010110: data <= 13'h0002; 
        10'b1011010111: data <= 13'h0001; 
        10'b1011011000: data <= 13'h0000; 
        10'b1011011001: data <= 13'h0005; 
        10'b1011011010: data <= 13'h0001; 
        10'b1011011011: data <= 13'h1ffe; 
        10'b1011011100: data <= 13'h0005; 
        10'b1011011101: data <= 13'h0008; 
        10'b1011011110: data <= 13'h000b; 
        10'b1011011111: data <= 13'h000f; 
        10'b1011100000: data <= 13'h0011; 
        10'b1011100001: data <= 13'h001a; 
        10'b1011100010: data <= 13'h001a; 
        10'b1011100011: data <= 13'h001e; 
        10'b1011100100: data <= 13'h0023; 
        10'b1011100101: data <= 13'h0023; 
        10'b1011100110: data <= 13'h002b; 
        10'b1011100111: data <= 13'h0019; 
        10'b1011101000: data <= 13'h0011; 
        10'b1011101001: data <= 13'h000e; 
        10'b1011101010: data <= 13'h0015; 
        10'b1011101011: data <= 13'h0017; 
        10'b1011101100: data <= 13'h0011; 
        10'b1011101101: data <= 13'h000c; 
        10'b1011101110: data <= 13'h0005; 
        10'b1011101111: data <= 13'h0002; 
        10'b1011110000: data <= 13'h0001; 
        10'b1011110001: data <= 13'h0002; 
        10'b1011110010: data <= 13'h1ffe; 
        10'b1011110011: data <= 13'h0001; 
        10'b1011110100: data <= 13'h1fff; 
        10'b1011110101: data <= 13'h0002; 
        10'b1011110110: data <= 13'h1ffe; 
        10'b1011110111: data <= 13'h0006; 
        10'b1011111000: data <= 13'h0003; 
        10'b1011111001: data <= 13'h0002; 
        10'b1011111010: data <= 13'h1fff; 
        10'b1011111011: data <= 13'h0006; 
        10'b1011111100: data <= 13'h0005; 
        10'b1011111101: data <= 13'h0003; 
        10'b1011111110: data <= 13'h1fff; 
        10'b1011111111: data <= 13'h1fff; 
        10'b1100000000: data <= 13'h0001; 
        10'b1100000001: data <= 13'h1fff; 
        10'b1100000010: data <= 13'h0001; 
        10'b1100000011: data <= 13'h0004; 
        10'b1100000100: data <= 13'h0000; 
        10'b1100000101: data <= 13'h0002; 
        10'b1100000110: data <= 13'h0007; 
        10'b1100000111: data <= 13'h0006; 
        10'b1100001000: data <= 13'h0003; 
        10'b1100001001: data <= 13'h0002; 
        10'b1100001010: data <= 13'h1ffe; 
        10'b1100001011: data <= 13'h0006; 
        10'b1100001100: data <= 13'h0004; 
        10'b1100001101: data <= 13'h1fff; 
        10'b1100001110: data <= 13'h0000; 
        10'b1100001111: data <= 13'h1fff; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 8) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 14'h0009; 
        10'b0000000001: data <= 14'h0008; 
        10'b0000000010: data <= 14'h3ffe; 
        10'b0000000011: data <= 14'h0006; 
        10'b0000000100: data <= 14'h0005; 
        10'b0000000101: data <= 14'h0008; 
        10'b0000000110: data <= 14'h3ffd; 
        10'b0000000111: data <= 14'h0002; 
        10'b0000001000: data <= 14'h000a; 
        10'b0000001001: data <= 14'h3ffc; 
        10'b0000001010: data <= 14'h3fff; 
        10'b0000001011: data <= 14'h0004; 
        10'b0000001100: data <= 14'h000c; 
        10'b0000001101: data <= 14'h0008; 
        10'b0000001110: data <= 14'h3ffb; 
        10'b0000001111: data <= 14'h3ffe; 
        10'b0000010000: data <= 14'h3ffd; 
        10'b0000010001: data <= 14'h0005; 
        10'b0000010010: data <= 14'h0009; 
        10'b0000010011: data <= 14'h0001; 
        10'b0000010100: data <= 14'h0001; 
        10'b0000010101: data <= 14'h3fff; 
        10'b0000010110: data <= 14'h3ffc; 
        10'b0000010111: data <= 14'h0001; 
        10'b0000011000: data <= 14'h000a; 
        10'b0000011001: data <= 14'h0003; 
        10'b0000011010: data <= 14'h3ffc; 
        10'b0000011011: data <= 14'h0005; 
        10'b0000011100: data <= 14'h0008; 
        10'b0000011101: data <= 14'h0007; 
        10'b0000011110: data <= 14'h0003; 
        10'b0000011111: data <= 14'h3ffe; 
        10'b0000100000: data <= 14'h3ffb; 
        10'b0000100001: data <= 14'h3ffc; 
        10'b0000100010: data <= 14'h3fff; 
        10'b0000100011: data <= 14'h000c; 
        10'b0000100100: data <= 14'h3ffb; 
        10'b0000100101: data <= 14'h000a; 
        10'b0000100110: data <= 14'h0004; 
        10'b0000100111: data <= 14'h0006; 
        10'b0000101000: data <= 14'h0005; 
        10'b0000101001: data <= 14'h0007; 
        10'b0000101010: data <= 14'h0000; 
        10'b0000101011: data <= 14'h3ffb; 
        10'b0000101100: data <= 14'h3ffd; 
        10'b0000101101: data <= 14'h0007; 
        10'b0000101110: data <= 14'h0000; 
        10'b0000101111: data <= 14'h0002; 
        10'b0000110000: data <= 14'h0009; 
        10'b0000110001: data <= 14'h3fff; 
        10'b0000110010: data <= 14'h0002; 
        10'b0000110011: data <= 14'h0001; 
        10'b0000110100: data <= 14'h0005; 
        10'b0000110101: data <= 14'h000a; 
        10'b0000110110: data <= 14'h0000; 
        10'b0000110111: data <= 14'h0002; 
        10'b0000111000: data <= 14'h000b; 
        10'b0000111001: data <= 14'h000b; 
        10'b0000111010: data <= 14'h0001; 
        10'b0000111011: data <= 14'h0007; 
        10'b0000111100: data <= 14'h0009; 
        10'b0000111101: data <= 14'h0000; 
        10'b0000111110: data <= 14'h3fff; 
        10'b0000111111: data <= 14'h0003; 
        10'b0001000000: data <= 14'h0009; 
        10'b0001000001: data <= 14'h3fff; 
        10'b0001000010: data <= 14'h3ffd; 
        10'b0001000011: data <= 14'h0007; 
        10'b0001000100: data <= 14'h0004; 
        10'b0001000101: data <= 14'h0009; 
        10'b0001000110: data <= 14'h3ffb; 
        10'b0001000111: data <= 14'h0009; 
        10'b0001001000: data <= 14'h3ffd; 
        10'b0001001001: data <= 14'h3ffc; 
        10'b0001001010: data <= 14'h0001; 
        10'b0001001011: data <= 14'h3ffc; 
        10'b0001001100: data <= 14'h000b; 
        10'b0001001101: data <= 14'h3ffd; 
        10'b0001001110: data <= 14'h3ffc; 
        10'b0001001111: data <= 14'h000a; 
        10'b0001010000: data <= 14'h0002; 
        10'b0001010001: data <= 14'h0002; 
        10'b0001010010: data <= 14'h0002; 
        10'b0001010011: data <= 14'h0005; 
        10'b0001010100: data <= 14'h000d; 
        10'b0001010101: data <= 14'h0000; 
        10'b0001010110: data <= 14'h3fff; 
        10'b0001010111: data <= 14'h0004; 
        10'b0001011000: data <= 14'h0004; 
        10'b0001011001: data <= 14'h3ffc; 
        10'b0001011010: data <= 14'h000b; 
        10'b0001011011: data <= 14'h0006; 
        10'b0001011100: data <= 14'h3ffe; 
        10'b0001011101: data <= 14'h000b; 
        10'b0001011110: data <= 14'h0003; 
        10'b0001011111: data <= 14'h0009; 
        10'b0001100000: data <= 14'h3fff; 
        10'b0001100001: data <= 14'h3ff6; 
        10'b0001100010: data <= 14'h3fff; 
        10'b0001100011: data <= 14'h3ff1; 
        10'b0001100100: data <= 14'h3ffe; 
        10'b0001100101: data <= 14'h3ff8; 
        10'b0001100110: data <= 14'h0003; 
        10'b0001100111: data <= 14'h0002; 
        10'b0001101000: data <= 14'h0003; 
        10'b0001101001: data <= 14'h3fff; 
        10'b0001101010: data <= 14'h0008; 
        10'b0001101011: data <= 14'h3fff; 
        10'b0001101100: data <= 14'h3fff; 
        10'b0001101101: data <= 14'h000c; 
        10'b0001101110: data <= 14'h0004; 
        10'b0001101111: data <= 14'h0007; 
        10'b0001110000: data <= 14'h0001; 
        10'b0001110001: data <= 14'h0002; 
        10'b0001110010: data <= 14'h0001; 
        10'b0001110011: data <= 14'h3ffd; 
        10'b0001110100: data <= 14'h3ffc; 
        10'b0001110101: data <= 14'h0008; 
        10'b0001110110: data <= 14'h0005; 
        10'b0001110111: data <= 14'h3fff; 
        10'b0001111000: data <= 14'h3ff9; 
        10'b0001111001: data <= 14'h0003; 
        10'b0001111010: data <= 14'h3ff5; 
        10'b0001111011: data <= 14'h3ff1; 
        10'b0001111100: data <= 14'h3fea; 
        10'b0001111101: data <= 14'h3fd9; 
        10'b0001111110: data <= 14'h3fce; 
        10'b0001111111: data <= 14'h3fbd; 
        10'b0010000000: data <= 14'h3fcf; 
        10'b0010000001: data <= 14'h3fce; 
        10'b0010000010: data <= 14'h3fdb; 
        10'b0010000011: data <= 14'h3ff0; 
        10'b0010000100: data <= 14'h3ff8; 
        10'b0010000101: data <= 14'h3ffb; 
        10'b0010000110: data <= 14'h0002; 
        10'b0010000111: data <= 14'h0009; 
        10'b0010001000: data <= 14'h0007; 
        10'b0010001001: data <= 14'h0007; 
        10'b0010001010: data <= 14'h0000; 
        10'b0010001011: data <= 14'h0000; 
        10'b0010001100: data <= 14'h0009; 
        10'b0010001101: data <= 14'h0006; 
        10'b0010001110: data <= 14'h0008; 
        10'b0010001111: data <= 14'h0005; 
        10'b0010010000: data <= 14'h0006; 
        10'b0010010001: data <= 14'h3ff9; 
        10'b0010010010: data <= 14'h3ffa; 
        10'b0010010011: data <= 14'h3ff9; 
        10'b0010010100: data <= 14'h3fe9; 
        10'b0010010101: data <= 14'h3fea; 
        10'b0010010110: data <= 14'h3fe8; 
        10'b0010010111: data <= 14'h3fe0; 
        10'b0010011000: data <= 14'h3fd8; 
        10'b0010011001: data <= 14'h3fd1; 
        10'b0010011010: data <= 14'h3fb8; 
        10'b0010011011: data <= 14'h3fb3; 
        10'b0010011100: data <= 14'h3f9e; 
        10'b0010011101: data <= 14'h3fc0; 
        10'b0010011110: data <= 14'h3fd7; 
        10'b0010011111: data <= 14'h3fec; 
        10'b0010100000: data <= 14'h3feb; 
        10'b0010100001: data <= 14'h3fe5; 
        10'b0010100010: data <= 14'h3fe7; 
        10'b0010100011: data <= 14'h3fee; 
        10'b0010100100: data <= 14'h3ff9; 
        10'b0010100101: data <= 14'h3ffd; 
        10'b0010100110: data <= 14'h0001; 
        10'b0010100111: data <= 14'h0006; 
        10'b0010101000: data <= 14'h0008; 
        10'b0010101001: data <= 14'h0008; 
        10'b0010101010: data <= 14'h3ffb; 
        10'b0010101011: data <= 14'h0008; 
        10'b0010101100: data <= 14'h0005; 
        10'b0010101101: data <= 14'h3fe8; 
        10'b0010101110: data <= 14'h3fe3; 
        10'b0010101111: data <= 14'h3fdd; 
        10'b0010110000: data <= 14'h3fd9; 
        10'b0010110001: data <= 14'h3fd0; 
        10'b0010110010: data <= 14'h3fdd; 
        10'b0010110011: data <= 14'h3ff5; 
        10'b0010110100: data <= 14'h0003; 
        10'b0010110101: data <= 14'h002b; 
        10'b0010110110: data <= 14'h0041; 
        10'b0010110111: data <= 14'h0033; 
        10'b0010111000: data <= 14'h0024; 
        10'b0010111001: data <= 14'h001e; 
        10'b0010111010: data <= 14'h0026; 
        10'b0010111011: data <= 14'h3ffa; 
        10'b0010111100: data <= 14'h3ff7; 
        10'b0010111101: data <= 14'h3fe3; 
        10'b0010111110: data <= 14'h3fcc; 
        10'b0010111111: data <= 14'h3fd0; 
        10'b0011000000: data <= 14'h3fe4; 
        10'b0011000001: data <= 14'h3ff3; 
        10'b0011000010: data <= 14'h3ffe; 
        10'b0011000011: data <= 14'h0004; 
        10'b0011000100: data <= 14'h000c; 
        10'b0011000101: data <= 14'h0000; 
        10'b0011000110: data <= 14'h3ffc; 
        10'b0011000111: data <= 14'h3ffc; 
        10'b0011001000: data <= 14'h3fe4; 
        10'b0011001001: data <= 14'h3fd6; 
        10'b0011001010: data <= 14'h3fcf; 
        10'b0011001011: data <= 14'h3fc5; 
        10'b0011001100: data <= 14'h3fc8; 
        10'b0011001101: data <= 14'h3fec; 
        10'b0011001110: data <= 14'h3ffe; 
        10'b0011001111: data <= 14'h000f; 
        10'b0011010000: data <= 14'h003b; 
        10'b0011010001: data <= 14'h0046; 
        10'b0011010010: data <= 14'h0060; 
        10'b0011010011: data <= 14'h0060; 
        10'b0011010100: data <= 14'h0064; 
        10'b0011010101: data <= 14'h002e; 
        10'b0011010110: data <= 14'h0022; 
        10'b0011010111: data <= 14'h0004; 
        10'b0011011000: data <= 14'h0009; 
        10'b0011011001: data <= 14'h000a; 
        10'b0011011010: data <= 14'h3fdd; 
        10'b0011011011: data <= 14'h3fc2; 
        10'b0011011100: data <= 14'h3fdb; 
        10'b0011011101: data <= 14'h3ff7; 
        10'b0011011110: data <= 14'h3ff7; 
        10'b0011011111: data <= 14'h0008; 
        10'b0011100000: data <= 14'h000c; 
        10'b0011100001: data <= 14'h000c; 
        10'b0011100010: data <= 14'h0006; 
        10'b0011100011: data <= 14'h3ffc; 
        10'b0011100100: data <= 14'h3fe3; 
        10'b0011100101: data <= 14'h3fd4; 
        10'b0011100110: data <= 14'h3fcd; 
        10'b0011100111: data <= 14'h3fb9; 
        10'b0011101000: data <= 14'h3fed; 
        10'b0011101001: data <= 14'h3ff7; 
        10'b0011101010: data <= 14'h3ff6; 
        10'b0011101011: data <= 14'h3fec; 
        10'b0011101100: data <= 14'h3ffe; 
        10'b0011101101: data <= 14'h001c; 
        10'b0011101110: data <= 14'h0052; 
        10'b0011101111: data <= 14'h002d; 
        10'b0011110000: data <= 14'h002e; 
        10'b0011110001: data <= 14'h0009; 
        10'b0011110010: data <= 14'h0004; 
        10'b0011110011: data <= 14'h0002; 
        10'b0011110100: data <= 14'h3ff1; 
        10'b0011110101: data <= 14'h0008; 
        10'b0011110110: data <= 14'h3fed; 
        10'b0011110111: data <= 14'h3fcf; 
        10'b0011111000: data <= 14'h3fd6; 
        10'b0011111001: data <= 14'h3fec; 
        10'b0011111010: data <= 14'h3ff7; 
        10'b0011111011: data <= 14'h000b; 
        10'b0011111100: data <= 14'h0004; 
        10'b0011111101: data <= 14'h0002; 
        10'b0011111110: data <= 14'h0001; 
        10'b0011111111: data <= 14'h3feb; 
        10'b0100000000: data <= 14'h3fd3; 
        10'b0100000001: data <= 14'h3fde; 
        10'b0100000010: data <= 14'h3ff6; 
        10'b0100000011: data <= 14'h3fec; 
        10'b0100000100: data <= 14'h3ff4; 
        10'b0100000101: data <= 14'h3ffb; 
        10'b0100000110: data <= 14'h0015; 
        10'b0100000111: data <= 14'h000d; 
        10'b0100001000: data <= 14'h0004; 
        10'b0100001001: data <= 14'h0022; 
        10'b0100001010: data <= 14'h0039; 
        10'b0100001011: data <= 14'h0033; 
        10'b0100001100: data <= 14'h3ffe; 
        10'b0100001101: data <= 14'h3ff1; 
        10'b0100001110: data <= 14'h0001; 
        10'b0100001111: data <= 14'h3fe2; 
        10'b0100010000: data <= 14'h3ff3; 
        10'b0100010001: data <= 14'h3fe0; 
        10'b0100010010: data <= 14'h3fde; 
        10'b0100010011: data <= 14'h3fdc; 
        10'b0100010100: data <= 14'h3fe7; 
        10'b0100010101: data <= 14'h3ff5; 
        10'b0100010110: data <= 14'h3ff8; 
        10'b0100010111: data <= 14'h000a; 
        10'b0100011000: data <= 14'h0002; 
        10'b0100011001: data <= 14'h0000; 
        10'b0100011010: data <= 14'h3ffb; 
        10'b0100011011: data <= 14'h3ff8; 
        10'b0100011100: data <= 14'h3fdd; 
        10'b0100011101: data <= 14'h3fee; 
        10'b0100011110: data <= 14'h0011; 
        10'b0100011111: data <= 14'h0016; 
        10'b0100100000: data <= 14'h002d; 
        10'b0100100001: data <= 14'h002c; 
        10'b0100100010: data <= 14'h0026; 
        10'b0100100011: data <= 14'h003a; 
        10'b0100100100: data <= 14'h001d; 
        10'b0100100101: data <= 14'h0007; 
        10'b0100100110: data <= 14'h0007; 
        10'b0100100111: data <= 14'h3fe3; 
        10'b0100101000: data <= 14'h3fef; 
        10'b0100101001: data <= 14'h3ffd; 
        10'b0100101010: data <= 14'h0014; 
        10'b0100101011: data <= 14'h0000; 
        10'b0100101100: data <= 14'h0010; 
        10'b0100101101: data <= 14'h3ff6; 
        10'b0100101110: data <= 14'h3fec; 
        10'b0100101111: data <= 14'h3fed; 
        10'b0100110000: data <= 14'h3fe8; 
        10'b0100110001: data <= 14'h3ff9; 
        10'b0100110010: data <= 14'h3ff7; 
        10'b0100110011: data <= 14'h0006; 
        10'b0100110100: data <= 14'h3ffe; 
        10'b0100110101: data <= 14'h0002; 
        10'b0100110110: data <= 14'h3ffb; 
        10'b0100110111: data <= 14'h3ffd; 
        10'b0100111000: data <= 14'h3ff7; 
        10'b0100111001: data <= 14'h0020; 
        10'b0100111010: data <= 14'h004a; 
        10'b0100111011: data <= 14'h0037; 
        10'b0100111100: data <= 14'h0056; 
        10'b0100111101: data <= 14'h0023; 
        10'b0100111110: data <= 14'h0024; 
        10'b0100111111: data <= 14'h003e; 
        10'b0101000000: data <= 14'h3fec; 
        10'b0101000001: data <= 14'h3fef; 
        10'b0101000010: data <= 14'h3ff7; 
        10'b0101000011: data <= 14'h0004; 
        10'b0101000100: data <= 14'h0018; 
        10'b0101000101: data <= 14'h0053; 
        10'b0101000110: data <= 14'h0027; 
        10'b0101000111: data <= 14'h0028; 
        10'b0101001000: data <= 14'h0041; 
        10'b0101001001: data <= 14'h002f; 
        10'b0101001010: data <= 14'h001c; 
        10'b0101001011: data <= 14'h0006; 
        10'b0101001100: data <= 14'h3ffb; 
        10'b0101001101: data <= 14'h3ff5; 
        10'b0101001110: data <= 14'h0000; 
        10'b0101001111: data <= 14'h0000; 
        10'b0101010000: data <= 14'h0005; 
        10'b0101010001: data <= 14'h000b; 
        10'b0101010010: data <= 14'h3ff9; 
        10'b0101010011: data <= 14'h3ff4; 
        10'b0101010100: data <= 14'h001b; 
        10'b0101010101: data <= 14'h0046; 
        10'b0101010110: data <= 14'h0051; 
        10'b0101010111: data <= 14'h0030; 
        10'b0101011000: data <= 14'h003c; 
        10'b0101011001: data <= 14'h0049; 
        10'b0101011010: data <= 14'h002f; 
        10'b0101011011: data <= 14'h0001; 
        10'b0101011100: data <= 14'h3fd1; 
        10'b0101011101: data <= 14'h0029; 
        10'b0101011110: data <= 14'h0058; 
        10'b0101011111: data <= 14'h0045; 
        10'b0101100000: data <= 14'h003b; 
        10'b0101100001: data <= 14'h005b; 
        10'b0101100010: data <= 14'h005b; 
        10'b0101100011: data <= 14'h005f; 
        10'b0101100100: data <= 14'h0062; 
        10'b0101100101: data <= 14'h0041; 
        10'b0101100110: data <= 14'h001f; 
        10'b0101100111: data <= 14'h0001; 
        10'b0101101000: data <= 14'h3ff1; 
        10'b0101101001: data <= 14'h0002; 
        10'b0101101010: data <= 14'h0005; 
        10'b0101101011: data <= 14'h0006; 
        10'b0101101100: data <= 14'h000c; 
        10'b0101101101: data <= 14'h0007; 
        10'b0101101110: data <= 14'h3ff6; 
        10'b0101101111: data <= 14'h0004; 
        10'b0101110000: data <= 14'h0029; 
        10'b0101110001: data <= 14'h003d; 
        10'b0101110010: data <= 14'h003a; 
        10'b0101110011: data <= 14'h0026; 
        10'b0101110100: data <= 14'h002f; 
        10'b0101110101: data <= 14'h001e; 
        10'b0101110110: data <= 14'h001c; 
        10'b0101110111: data <= 14'h3ff2; 
        10'b0101111000: data <= 14'h3fe7; 
        10'b0101111001: data <= 14'h0040; 
        10'b0101111010: data <= 14'h0058; 
        10'b0101111011: data <= 14'h003f; 
        10'b0101111100: data <= 14'h0049; 
        10'b0101111101: data <= 14'h0042; 
        10'b0101111110: data <= 14'h005a; 
        10'b0101111111: data <= 14'h005b; 
        10'b0110000000: data <= 14'h0047; 
        10'b0110000001: data <= 14'h002a; 
        10'b0110000010: data <= 14'h0002; 
        10'b0110000011: data <= 14'h3fe4; 
        10'b0110000100: data <= 14'h3fef; 
        10'b0110000101: data <= 14'h3ffb; 
        10'b0110000110: data <= 14'h0005; 
        10'b0110000111: data <= 14'h0005; 
        10'b0110001000: data <= 14'h0002; 
        10'b0110001001: data <= 14'h0001; 
        10'b0110001010: data <= 14'h0008; 
        10'b0110001011: data <= 14'h0005; 
        10'b0110001100: data <= 14'h0013; 
        10'b0110001101: data <= 14'h0012; 
        10'b0110001110: data <= 14'h0030; 
        10'b0110001111: data <= 14'h0021; 
        10'b0110010000: data <= 14'h0010; 
        10'b0110010001: data <= 14'h0000; 
        10'b0110010010: data <= 14'h0006; 
        10'b0110010011: data <= 14'h3ffd; 
        10'b0110010100: data <= 14'h3fee; 
        10'b0110010101: data <= 14'h0015; 
        10'b0110010110: data <= 14'h000c; 
        10'b0110010111: data <= 14'h0038; 
        10'b0110011000: data <= 14'h003b; 
        10'b0110011001: data <= 14'h003b; 
        10'b0110011010: data <= 14'h0028; 
        10'b0110011011: data <= 14'h001a; 
        10'b0110011100: data <= 14'h0020; 
        10'b0110011101: data <= 14'h0001; 
        10'b0110011110: data <= 14'h3fdf; 
        10'b0110011111: data <= 14'h3fd0; 
        10'b0110100000: data <= 14'h3fec; 
        10'b0110100001: data <= 14'h0003; 
        10'b0110100010: data <= 14'h0002; 
        10'b0110100011: data <= 14'h0002; 
        10'b0110100100: data <= 14'h0009; 
        10'b0110100101: data <= 14'h0008; 
        10'b0110100110: data <= 14'h0006; 
        10'b0110100111: data <= 14'h3ff9; 
        10'b0110101000: data <= 14'h0001; 
        10'b0110101001: data <= 14'h0015; 
        10'b0110101010: data <= 14'h0014; 
        10'b0110101011: data <= 14'h000d; 
        10'b0110101100: data <= 14'h000e; 
        10'b0110101101: data <= 14'h3fe7; 
        10'b0110101110: data <= 14'h3ff4; 
        10'b0110101111: data <= 14'h3ff4; 
        10'b0110110000: data <= 14'h3fee; 
        10'b0110110001: data <= 14'h3ff2; 
        10'b0110110010: data <= 14'h3ff0; 
        10'b0110110011: data <= 14'h003d; 
        10'b0110110100: data <= 14'h005a; 
        10'b0110110101: data <= 14'h0056; 
        10'b0110110110: data <= 14'h002b; 
        10'b0110110111: data <= 14'h0004; 
        10'b0110111000: data <= 14'h3fed; 
        10'b0110111001: data <= 14'h3fcf; 
        10'b0110111010: data <= 14'h3fc3; 
        10'b0110111011: data <= 14'h3fd4; 
        10'b0110111100: data <= 14'h3fec; 
        10'b0110111101: data <= 14'h0000; 
        10'b0110111110: data <= 14'h0005; 
        10'b0110111111: data <= 14'h3fff; 
        10'b0111000000: data <= 14'h000b; 
        10'b0111000001: data <= 14'h0001; 
        10'b0111000010: data <= 14'h3ff8; 
        10'b0111000011: data <= 14'h3ffe; 
        10'b0111000100: data <= 14'h0001; 
        10'b0111000101: data <= 14'h0006; 
        10'b0111000110: data <= 14'h3ff0; 
        10'b0111000111: data <= 14'h000d; 
        10'b0111001000: data <= 14'h0025; 
        10'b0111001001: data <= 14'h3ff7; 
        10'b0111001010: data <= 14'h0015; 
        10'b0111001011: data <= 14'h001e; 
        10'b0111001100: data <= 14'h3ffc; 
        10'b0111001101: data <= 14'h3fde; 
        10'b0111001110: data <= 14'h3ffa; 
        10'b0111001111: data <= 14'h0022; 
        10'b0111010000: data <= 14'h003d; 
        10'b0111010001: data <= 14'h003d; 
        10'b0111010010: data <= 14'h000f; 
        10'b0111010011: data <= 14'h3fdd; 
        10'b0111010100: data <= 14'h3fc7; 
        10'b0111010101: data <= 14'h3fb1; 
        10'b0111010110: data <= 14'h3fc8; 
        10'b0111010111: data <= 14'h3fd3; 
        10'b0111011000: data <= 14'h3fe2; 
        10'b0111011001: data <= 14'h0001; 
        10'b0111011010: data <= 14'h3ff9; 
        10'b0111011011: data <= 14'h0006; 
        10'b0111011100: data <= 14'h0003; 
        10'b0111011101: data <= 14'h3ffe; 
        10'b0111011110: data <= 14'h3ff8; 
        10'b0111011111: data <= 14'h3ff4; 
        10'b0111100000: data <= 14'h3fe9; 
        10'b0111100001: data <= 14'h3fe5; 
        10'b0111100010: data <= 14'h3fe9; 
        10'b0111100011: data <= 14'h000a; 
        10'b0111100100: data <= 14'h0014; 
        10'b0111100101: data <= 14'h0017; 
        10'b0111100110: data <= 14'h0022; 
        10'b0111100111: data <= 14'h0032; 
        10'b0111101000: data <= 14'h001f; 
        10'b0111101001: data <= 14'h000e; 
        10'b0111101010: data <= 14'h0013; 
        10'b0111101011: data <= 14'h0032; 
        10'b0111101100: data <= 14'h000f; 
        10'b0111101101: data <= 14'h3ff6; 
        10'b0111101110: data <= 14'h3fea; 
        10'b0111101111: data <= 14'h3fcd; 
        10'b0111110000: data <= 14'h3fce; 
        10'b0111110001: data <= 14'h3fca; 
        10'b0111110010: data <= 14'h3fcd; 
        10'b0111110011: data <= 14'h3fdb; 
        10'b0111110100: data <= 14'h3fe5; 
        10'b0111110101: data <= 14'h0003; 
        10'b0111110110: data <= 14'h0003; 
        10'b0111110111: data <= 14'h3ffe; 
        10'b0111111000: data <= 14'h000a; 
        10'b0111111001: data <= 14'h0000; 
        10'b0111111010: data <= 14'h3ffa; 
        10'b0111111011: data <= 14'h3ffe; 
        10'b0111111100: data <= 14'h3fec; 
        10'b0111111101: data <= 14'h3fd3; 
        10'b0111111110: data <= 14'h3fd2; 
        10'b0111111111: data <= 14'h3fd3; 
        10'b1000000000: data <= 14'h3fed; 
        10'b1000000001: data <= 14'h0008; 
        10'b1000000010: data <= 14'h0037; 
        10'b1000000011: data <= 14'h002c; 
        10'b1000000100: data <= 14'h3fe5; 
        10'b1000000101: data <= 14'h3fe5; 
        10'b1000000110: data <= 14'h0002; 
        10'b1000000111: data <= 14'h0021; 
        10'b1000001000: data <= 14'h3fec; 
        10'b1000001001: data <= 14'h3fe9; 
        10'b1000001010: data <= 14'h3fd5; 
        10'b1000001011: data <= 14'h3fe6; 
        10'b1000001100: data <= 14'h3fe8; 
        10'b1000001101: data <= 14'h3fda; 
        10'b1000001110: data <= 14'h3fd8; 
        10'b1000001111: data <= 14'h3fd6; 
        10'b1000010000: data <= 14'h3fe2; 
        10'b1000010001: data <= 14'h3ffb; 
        10'b1000010010: data <= 14'h0001; 
        10'b1000010011: data <= 14'h0009; 
        10'b1000010100: data <= 14'h0006; 
        10'b1000010101: data <= 14'h000d; 
        10'b1000010110: data <= 14'h0002; 
        10'b1000010111: data <= 14'h3ff5; 
        10'b1000011000: data <= 14'h3fee; 
        10'b1000011001: data <= 14'h3fe0; 
        10'b1000011010: data <= 14'h3fcd; 
        10'b1000011011: data <= 14'h3fcc; 
        10'b1000011100: data <= 14'h3fca; 
        10'b1000011101: data <= 14'h3fca; 
        10'b1000011110: data <= 14'h3fc4; 
        10'b1000011111: data <= 14'h3fcd; 
        10'b1000100000: data <= 14'h3fbe; 
        10'b1000100001: data <= 14'h3fd2; 
        10'b1000100010: data <= 14'h3fd9; 
        10'b1000100011: data <= 14'h3fd4; 
        10'b1000100100: data <= 14'h3fda; 
        10'b1000100101: data <= 14'h3ff4; 
        10'b1000100110: data <= 14'h3fe3; 
        10'b1000100111: data <= 14'h3ff8; 
        10'b1000101000: data <= 14'h3fed; 
        10'b1000101001: data <= 14'h3fe9; 
        10'b1000101010: data <= 14'h3fea; 
        10'b1000101011: data <= 14'h3fed; 
        10'b1000101100: data <= 14'h3ff4; 
        10'b1000101101: data <= 14'h0003; 
        10'b1000101110: data <= 14'h3ffc; 
        10'b1000101111: data <= 14'h0001; 
        10'b1000110000: data <= 14'h3ffe; 
        10'b1000110001: data <= 14'h0002; 
        10'b1000110010: data <= 14'h0005; 
        10'b1000110011: data <= 14'h0000; 
        10'b1000110100: data <= 14'h3fed; 
        10'b1000110101: data <= 14'h3fe1; 
        10'b1000110110: data <= 14'h3fd1; 
        10'b1000110111: data <= 14'h3fb6; 
        10'b1000111000: data <= 14'h3fac; 
        10'b1000111001: data <= 14'h3fa1; 
        10'b1000111010: data <= 14'h3f80; 
        10'b1000111011: data <= 14'h3f9e; 
        10'b1000111100: data <= 14'h3fa0; 
        10'b1000111101: data <= 14'h3fe1; 
        10'b1000111110: data <= 14'h3fd4; 
        10'b1000111111: data <= 14'h3feb; 
        10'b1001000000: data <= 14'h3fe7; 
        10'b1001000001: data <= 14'h3ff9; 
        10'b1001000010: data <= 14'h3fd6; 
        10'b1001000011: data <= 14'h3ff2; 
        10'b1001000100: data <= 14'h3fef; 
        10'b1001000101: data <= 14'h3fe5; 
        10'b1001000110: data <= 14'h3ff8; 
        10'b1001000111: data <= 14'h3ff3; 
        10'b1001001000: data <= 14'h0001; 
        10'b1001001001: data <= 14'h000b; 
        10'b1001001010: data <= 14'h0006; 
        10'b1001001011: data <= 14'h0002; 
        10'b1001001100: data <= 14'h0001; 
        10'b1001001101: data <= 14'h0000; 
        10'b1001001110: data <= 14'h000b; 
        10'b1001001111: data <= 14'h3ff5; 
        10'b1001010000: data <= 14'h3ff3; 
        10'b1001010001: data <= 14'h3fe1; 
        10'b1001010010: data <= 14'h3fd5; 
        10'b1001010011: data <= 14'h3fbd; 
        10'b1001010100: data <= 14'h3fb4; 
        10'b1001010101: data <= 14'h3fad; 
        10'b1001010110: data <= 14'h3fa9; 
        10'b1001010111: data <= 14'h3fb1; 
        10'b1001011000: data <= 14'h3fce; 
        10'b1001011001: data <= 14'h3fcf; 
        10'b1001011010: data <= 14'h3fce; 
        10'b1001011011: data <= 14'h3fe3; 
        10'b1001011100: data <= 14'h3fe1; 
        10'b1001011101: data <= 14'h3fd1; 
        10'b1001011110: data <= 14'h3fc7; 
        10'b1001011111: data <= 14'h3fe8; 
        10'b1001100000: data <= 14'h3ff3; 
        10'b1001100001: data <= 14'h3ff8; 
        10'b1001100010: data <= 14'h0004; 
        10'b1001100011: data <= 14'h3fff; 
        10'b1001100100: data <= 14'h0005; 
        10'b1001100101: data <= 14'h0007; 
        10'b1001100110: data <= 14'h0000; 
        10'b1001100111: data <= 14'h0001; 
        10'b1001101000: data <= 14'h0008; 
        10'b1001101001: data <= 14'h0002; 
        10'b1001101010: data <= 14'h0002; 
        10'b1001101011: data <= 14'h0008; 
        10'b1001101100: data <= 14'h3ffb; 
        10'b1001101101: data <= 14'h3fe7; 
        10'b1001101110: data <= 14'h3fd8; 
        10'b1001101111: data <= 14'h3fca; 
        10'b1001110000: data <= 14'h3fd8; 
        10'b1001110001: data <= 14'h3fd6; 
        10'b1001110010: data <= 14'h3fd2; 
        10'b1001110011: data <= 14'h3fe1; 
        10'b1001110100: data <= 14'h3fdd; 
        10'b1001110101: data <= 14'h3fd2; 
        10'b1001110110: data <= 14'h3fd9; 
        10'b1001110111: data <= 14'h3fca; 
        10'b1001111000: data <= 14'h3fc4; 
        10'b1001111001: data <= 14'h3fc5; 
        10'b1001111010: data <= 14'h3fcf; 
        10'b1001111011: data <= 14'h3fd4; 
        10'b1001111100: data <= 14'h3ff4; 
        10'b1001111101: data <= 14'h000f; 
        10'b1001111110: data <= 14'h0008; 
        10'b1001111111: data <= 14'h000a; 
        10'b1010000000: data <= 14'h0011; 
        10'b1010000001: data <= 14'h0003; 
        10'b1010000010: data <= 14'h0004; 
        10'b1010000011: data <= 14'h0006; 
        10'b1010000100: data <= 14'h000a; 
        10'b1010000101: data <= 14'h0008; 
        10'b1010000110: data <= 14'h0003; 
        10'b1010000111: data <= 14'h3ffc; 
        10'b1010001000: data <= 14'h3ff9; 
        10'b1010001001: data <= 14'h3feb; 
        10'b1010001010: data <= 14'h3fe7; 
        10'b1010001011: data <= 14'h3fdf; 
        10'b1010001100: data <= 14'h3ffe; 
        10'b1010001101: data <= 14'h3ff3; 
        10'b1010001110: data <= 14'h3ff5; 
        10'b1010001111: data <= 14'h3fd8; 
        10'b1010010000: data <= 14'h3fe0; 
        10'b1010010001: data <= 14'h3fd7; 
        10'b1010010010: data <= 14'h3fde; 
        10'b1010010011: data <= 14'h3fc5; 
        10'b1010010100: data <= 14'h3fc1; 
        10'b1010010101: data <= 14'h3fc8; 
        10'b1010010110: data <= 14'h3fdd; 
        10'b1010010111: data <= 14'h3ffd; 
        10'b1010011000: data <= 14'h000e; 
        10'b1010011001: data <= 14'h0020; 
        10'b1010011010: data <= 14'h002e; 
        10'b1010011011: data <= 14'h0026; 
        10'b1010011100: data <= 14'h0012; 
        10'b1010011101: data <= 14'h3fff; 
        10'b1010011110: data <= 14'h000d; 
        10'b1010011111: data <= 14'h3fff; 
        10'b1010100000: data <= 14'h0000; 
        10'b1010100001: data <= 14'h3ffb; 
        10'b1010100010: data <= 14'h3fff; 
        10'b1010100011: data <= 14'h000b; 
        10'b1010100100: data <= 14'h0008; 
        10'b1010100101: data <= 14'h000c; 
        10'b1010100110: data <= 14'h0009; 
        10'b1010100111: data <= 14'h000d; 
        10'b1010101000: data <= 14'h0012; 
        10'b1010101001: data <= 14'h000a; 
        10'b1010101010: data <= 14'h3ffa; 
        10'b1010101011: data <= 14'h3fec; 
        10'b1010101100: data <= 14'h3fff; 
        10'b1010101101: data <= 14'h3fe1; 
        10'b1010101110: data <= 14'h3fd9; 
        10'b1010101111: data <= 14'h3fd6; 
        10'b1010110000: data <= 14'h3fed; 
        10'b1010110001: data <= 14'h000e; 
        10'b1010110010: data <= 14'h0017; 
        10'b1010110011: data <= 14'h0018; 
        10'b1010110100: data <= 14'h0037; 
        10'b1010110101: data <= 14'h003b; 
        10'b1010110110: data <= 14'h0022; 
        10'b1010110111: data <= 14'h0015; 
        10'b1010111000: data <= 14'h0010; 
        10'b1010111001: data <= 14'h3ffd; 
        10'b1010111010: data <= 14'h0007; 
        10'b1010111011: data <= 14'h0000; 
        10'b1010111100: data <= 14'h0003; 
        10'b1010111101: data <= 14'h000b; 
        10'b1010111110: data <= 14'h000b; 
        10'b1010111111: data <= 14'h3fff; 
        10'b1011000000: data <= 14'h0001; 
        10'b1011000001: data <= 14'h0012; 
        10'b1011000010: data <= 14'h000e; 
        10'b1011000011: data <= 14'h0028; 
        10'b1011000100: data <= 14'h002c; 
        10'b1011000101: data <= 14'h002d; 
        10'b1011000110: data <= 14'h0027; 
        10'b1011000111: data <= 14'h000f; 
        10'b1011001000: data <= 14'h0029; 
        10'b1011001001: data <= 14'h0024; 
        10'b1011001010: data <= 14'h0023; 
        10'b1011001011: data <= 14'h0021; 
        10'b1011001100: data <= 14'h003d; 
        10'b1011001101: data <= 14'h0042; 
        10'b1011001110: data <= 14'h0049; 
        10'b1011001111: data <= 14'h004c; 
        10'b1011010000: data <= 14'h0055; 
        10'b1011010001: data <= 14'h003c; 
        10'b1011010010: data <= 14'h0018; 
        10'b1011010011: data <= 14'h000b; 
        10'b1011010100: data <= 14'h3fff; 
        10'b1011010101: data <= 14'h3fff; 
        10'b1011010110: data <= 14'h0003; 
        10'b1011010111: data <= 14'h0003; 
        10'b1011011000: data <= 14'h0000; 
        10'b1011011001: data <= 14'h000a; 
        10'b1011011010: data <= 14'h0003; 
        10'b1011011011: data <= 14'h3ffc; 
        10'b1011011100: data <= 14'h000a; 
        10'b1011011101: data <= 14'h000f; 
        10'b1011011110: data <= 14'h0015; 
        10'b1011011111: data <= 14'h001e; 
        10'b1011100000: data <= 14'h0022; 
        10'b1011100001: data <= 14'h0033; 
        10'b1011100010: data <= 14'h0035; 
        10'b1011100011: data <= 14'h003b; 
        10'b1011100100: data <= 14'h0046; 
        10'b1011100101: data <= 14'h0047; 
        10'b1011100110: data <= 14'h0057; 
        10'b1011100111: data <= 14'h0032; 
        10'b1011101000: data <= 14'h0022; 
        10'b1011101001: data <= 14'h001d; 
        10'b1011101010: data <= 14'h002b; 
        10'b1011101011: data <= 14'h002e; 
        10'b1011101100: data <= 14'h0021; 
        10'b1011101101: data <= 14'h0017; 
        10'b1011101110: data <= 14'h000a; 
        10'b1011101111: data <= 14'h0003; 
        10'b1011110000: data <= 14'h0002; 
        10'b1011110001: data <= 14'h0004; 
        10'b1011110010: data <= 14'h3ffc; 
        10'b1011110011: data <= 14'h0002; 
        10'b1011110100: data <= 14'h3ffe; 
        10'b1011110101: data <= 14'h0004; 
        10'b1011110110: data <= 14'h3ffc; 
        10'b1011110111: data <= 14'h000c; 
        10'b1011111000: data <= 14'h0007; 
        10'b1011111001: data <= 14'h0004; 
        10'b1011111010: data <= 14'h3ffe; 
        10'b1011111011: data <= 14'h000b; 
        10'b1011111100: data <= 14'h000a; 
        10'b1011111101: data <= 14'h0007; 
        10'b1011111110: data <= 14'h3ffe; 
        10'b1011111111: data <= 14'h3ffe; 
        10'b1100000000: data <= 14'h0002; 
        10'b1100000001: data <= 14'h3ffe; 
        10'b1100000010: data <= 14'h0002; 
        10'b1100000011: data <= 14'h0007; 
        10'b1100000100: data <= 14'h0001; 
        10'b1100000101: data <= 14'h0004; 
        10'b1100000110: data <= 14'h000d; 
        10'b1100000111: data <= 14'h000c; 
        10'b1100001000: data <= 14'h0007; 
        10'b1100001001: data <= 14'h0004; 
        10'b1100001010: data <= 14'h3ffd; 
        10'b1100001011: data <= 14'h000d; 
        10'b1100001100: data <= 14'h0007; 
        10'b1100001101: data <= 14'h3ffe; 
        10'b1100001110: data <= 14'h0001; 
        10'b1100001111: data <= 14'h3fff; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 9) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 15'h0012; 
        10'b0000000001: data <= 15'h0010; 
        10'b0000000010: data <= 15'h7ffb; 
        10'b0000000011: data <= 15'h000b; 
        10'b0000000100: data <= 15'h000a; 
        10'b0000000101: data <= 15'h0011; 
        10'b0000000110: data <= 15'h7ffa; 
        10'b0000000111: data <= 15'h0003; 
        10'b0000001000: data <= 15'h0013; 
        10'b0000001001: data <= 15'h7ff8; 
        10'b0000001010: data <= 15'h7ffe; 
        10'b0000001011: data <= 15'h0008; 
        10'b0000001100: data <= 15'h0018; 
        10'b0000001101: data <= 15'h0010; 
        10'b0000001110: data <= 15'h7ff6; 
        10'b0000001111: data <= 15'h7ffb; 
        10'b0000010000: data <= 15'h7ffb; 
        10'b0000010001: data <= 15'h0009; 
        10'b0000010010: data <= 15'h0011; 
        10'b0000010011: data <= 15'h0001; 
        10'b0000010100: data <= 15'h0002; 
        10'b0000010101: data <= 15'h7fff; 
        10'b0000010110: data <= 15'h7ff8; 
        10'b0000010111: data <= 15'h0003; 
        10'b0000011000: data <= 15'h0014; 
        10'b0000011001: data <= 15'h0006; 
        10'b0000011010: data <= 15'h7ff7; 
        10'b0000011011: data <= 15'h000a; 
        10'b0000011100: data <= 15'h0010; 
        10'b0000011101: data <= 15'h000e; 
        10'b0000011110: data <= 15'h0007; 
        10'b0000011111: data <= 15'h7ffc; 
        10'b0000100000: data <= 15'h7ff7; 
        10'b0000100001: data <= 15'h7ff8; 
        10'b0000100010: data <= 15'h7ffe; 
        10'b0000100011: data <= 15'h0018; 
        10'b0000100100: data <= 15'h7ff7; 
        10'b0000100101: data <= 15'h0014; 
        10'b0000100110: data <= 15'h0008; 
        10'b0000100111: data <= 15'h000c; 
        10'b0000101000: data <= 15'h0009; 
        10'b0000101001: data <= 15'h000e; 
        10'b0000101010: data <= 15'h0000; 
        10'b0000101011: data <= 15'h7ff5; 
        10'b0000101100: data <= 15'h7ffb; 
        10'b0000101101: data <= 15'h000f; 
        10'b0000101110: data <= 15'h7fff; 
        10'b0000101111: data <= 15'h0004; 
        10'b0000110000: data <= 15'h0013; 
        10'b0000110001: data <= 15'h7fff; 
        10'b0000110010: data <= 15'h0003; 
        10'b0000110011: data <= 15'h0002; 
        10'b0000110100: data <= 15'h000a; 
        10'b0000110101: data <= 15'h0014; 
        10'b0000110110: data <= 15'h0000; 
        10'b0000110111: data <= 15'h0004; 
        10'b0000111000: data <= 15'h0015; 
        10'b0000111001: data <= 15'h0016; 
        10'b0000111010: data <= 15'h0002; 
        10'b0000111011: data <= 15'h000f; 
        10'b0000111100: data <= 15'h0012; 
        10'b0000111101: data <= 15'h7fff; 
        10'b0000111110: data <= 15'h7ffe; 
        10'b0000111111: data <= 15'h0007; 
        10'b0001000000: data <= 15'h0012; 
        10'b0001000001: data <= 15'h7ffd; 
        10'b0001000010: data <= 15'h7ffa; 
        10'b0001000011: data <= 15'h000e; 
        10'b0001000100: data <= 15'h0008; 
        10'b0001000101: data <= 15'h0011; 
        10'b0001000110: data <= 15'h7ff6; 
        10'b0001000111: data <= 15'h0012; 
        10'b0001001000: data <= 15'h7ff9; 
        10'b0001001001: data <= 15'h7ff9; 
        10'b0001001010: data <= 15'h0002; 
        10'b0001001011: data <= 15'h7ff7; 
        10'b0001001100: data <= 15'h0015; 
        10'b0001001101: data <= 15'h7ffa; 
        10'b0001001110: data <= 15'h7ff8; 
        10'b0001001111: data <= 15'h0015; 
        10'b0001010000: data <= 15'h0004; 
        10'b0001010001: data <= 15'h0004; 
        10'b0001010010: data <= 15'h0005; 
        10'b0001010011: data <= 15'h0009; 
        10'b0001010100: data <= 15'h001a; 
        10'b0001010101: data <= 15'h0001; 
        10'b0001010110: data <= 15'h7ffe; 
        10'b0001010111: data <= 15'h0008; 
        10'b0001011000: data <= 15'h0008; 
        10'b0001011001: data <= 15'h7ff7; 
        10'b0001011010: data <= 15'h0015; 
        10'b0001011011: data <= 15'h000c; 
        10'b0001011100: data <= 15'h7ffc; 
        10'b0001011101: data <= 15'h0016; 
        10'b0001011110: data <= 15'h0007; 
        10'b0001011111: data <= 15'h0011; 
        10'b0001100000: data <= 15'h7ffe; 
        10'b0001100001: data <= 15'h7fed; 
        10'b0001100010: data <= 15'h7ffe; 
        10'b0001100011: data <= 15'h7fe2; 
        10'b0001100100: data <= 15'h7ffc; 
        10'b0001100101: data <= 15'h7ff1; 
        10'b0001100110: data <= 15'h0005; 
        10'b0001100111: data <= 15'h0003; 
        10'b0001101000: data <= 15'h0007; 
        10'b0001101001: data <= 15'h7ffe; 
        10'b0001101010: data <= 15'h0011; 
        10'b0001101011: data <= 15'h7ffe; 
        10'b0001101100: data <= 15'h7ffd; 
        10'b0001101101: data <= 15'h0017; 
        10'b0001101110: data <= 15'h0009; 
        10'b0001101111: data <= 15'h000f; 
        10'b0001110000: data <= 15'h0003; 
        10'b0001110001: data <= 15'h0005; 
        10'b0001110010: data <= 15'h0001; 
        10'b0001110011: data <= 15'h7ffb; 
        10'b0001110100: data <= 15'h7ff8; 
        10'b0001110101: data <= 15'h000f; 
        10'b0001110110: data <= 15'h000a; 
        10'b0001110111: data <= 15'h7ffe; 
        10'b0001111000: data <= 15'h7ff3; 
        10'b0001111001: data <= 15'h0005; 
        10'b0001111010: data <= 15'h7fea; 
        10'b0001111011: data <= 15'h7fe1; 
        10'b0001111100: data <= 15'h7fd5; 
        10'b0001111101: data <= 15'h7fb1; 
        10'b0001111110: data <= 15'h7f9c; 
        10'b0001111111: data <= 15'h7f7a; 
        10'b0010000000: data <= 15'h7f9d; 
        10'b0010000001: data <= 15'h7f9d; 
        10'b0010000010: data <= 15'h7fb6; 
        10'b0010000011: data <= 15'h7fe0; 
        10'b0010000100: data <= 15'h7ff1; 
        10'b0010000101: data <= 15'h7ff5; 
        10'b0010000110: data <= 15'h0004; 
        10'b0010000111: data <= 15'h0013; 
        10'b0010001000: data <= 15'h000f; 
        10'b0010001001: data <= 15'h000e; 
        10'b0010001010: data <= 15'h0000; 
        10'b0010001011: data <= 15'h0001; 
        10'b0010001100: data <= 15'h0012; 
        10'b0010001101: data <= 15'h000d; 
        10'b0010001110: data <= 15'h000f; 
        10'b0010001111: data <= 15'h000a; 
        10'b0010010000: data <= 15'h000b; 
        10'b0010010001: data <= 15'h7ff2; 
        10'b0010010010: data <= 15'h7ff3; 
        10'b0010010011: data <= 15'h7ff2; 
        10'b0010010100: data <= 15'h7fd3; 
        10'b0010010101: data <= 15'h7fd3; 
        10'b0010010110: data <= 15'h7fd0; 
        10'b0010010111: data <= 15'h7fc1; 
        10'b0010011000: data <= 15'h7fb1; 
        10'b0010011001: data <= 15'h7fa2; 
        10'b0010011010: data <= 15'h7f71; 
        10'b0010011011: data <= 15'h7f65; 
        10'b0010011100: data <= 15'h7f3c; 
        10'b0010011101: data <= 15'h7f7f; 
        10'b0010011110: data <= 15'h7faf; 
        10'b0010011111: data <= 15'h7fd9; 
        10'b0010100000: data <= 15'h7fd6; 
        10'b0010100001: data <= 15'h7fca; 
        10'b0010100010: data <= 15'h7fce; 
        10'b0010100011: data <= 15'h7fdc; 
        10'b0010100100: data <= 15'h7ff2; 
        10'b0010100101: data <= 15'h7ff9; 
        10'b0010100110: data <= 15'h0002; 
        10'b0010100111: data <= 15'h000d; 
        10'b0010101000: data <= 15'h0010; 
        10'b0010101001: data <= 15'h0011; 
        10'b0010101010: data <= 15'h7ff6; 
        10'b0010101011: data <= 15'h0011; 
        10'b0010101100: data <= 15'h000b; 
        10'b0010101101: data <= 15'h7fd0; 
        10'b0010101110: data <= 15'h7fc5; 
        10'b0010101111: data <= 15'h7fbb; 
        10'b0010110000: data <= 15'h7fb2; 
        10'b0010110001: data <= 15'h7fa0; 
        10'b0010110010: data <= 15'h7fba; 
        10'b0010110011: data <= 15'h7fe9; 
        10'b0010110100: data <= 15'h0006; 
        10'b0010110101: data <= 15'h0057; 
        10'b0010110110: data <= 15'h0081; 
        10'b0010110111: data <= 15'h0067; 
        10'b0010111000: data <= 15'h0048; 
        10'b0010111001: data <= 15'h003c; 
        10'b0010111010: data <= 15'h004c; 
        10'b0010111011: data <= 15'h7ff3; 
        10'b0010111100: data <= 15'h7fee; 
        10'b0010111101: data <= 15'h7fc6; 
        10'b0010111110: data <= 15'h7f99; 
        10'b0010111111: data <= 15'h7fa0; 
        10'b0011000000: data <= 15'h7fc9; 
        10'b0011000001: data <= 15'h7fe5; 
        10'b0011000010: data <= 15'h7ffc; 
        10'b0011000011: data <= 15'h0009; 
        10'b0011000100: data <= 15'h0019; 
        10'b0011000101: data <= 15'h7fff; 
        10'b0011000110: data <= 15'h7ff8; 
        10'b0011000111: data <= 15'h7ff7; 
        10'b0011001000: data <= 15'h7fc9; 
        10'b0011001001: data <= 15'h7fac; 
        10'b0011001010: data <= 15'h7f9d; 
        10'b0011001011: data <= 15'h7f8a; 
        10'b0011001100: data <= 15'h7f91; 
        10'b0011001101: data <= 15'h7fd9; 
        10'b0011001110: data <= 15'h7ffd; 
        10'b0011001111: data <= 15'h001f; 
        10'b0011010000: data <= 15'h0075; 
        10'b0011010001: data <= 15'h008c; 
        10'b0011010010: data <= 15'h00c0; 
        10'b0011010011: data <= 15'h00c1; 
        10'b0011010100: data <= 15'h00c9; 
        10'b0011010101: data <= 15'h005b; 
        10'b0011010110: data <= 15'h0045; 
        10'b0011010111: data <= 15'h0007; 
        10'b0011011000: data <= 15'h0012; 
        10'b0011011001: data <= 15'h0014; 
        10'b0011011010: data <= 15'h7fbb; 
        10'b0011011011: data <= 15'h7f84; 
        10'b0011011100: data <= 15'h7fb7; 
        10'b0011011101: data <= 15'h7fee; 
        10'b0011011110: data <= 15'h7fed; 
        10'b0011011111: data <= 15'h0010; 
        10'b0011100000: data <= 15'h0018; 
        10'b0011100001: data <= 15'h0018; 
        10'b0011100010: data <= 15'h000c; 
        10'b0011100011: data <= 15'h7ff9; 
        10'b0011100100: data <= 15'h7fc6; 
        10'b0011100101: data <= 15'h7fa9; 
        10'b0011100110: data <= 15'h7f9b; 
        10'b0011100111: data <= 15'h7f72; 
        10'b0011101000: data <= 15'h7fdb; 
        10'b0011101001: data <= 15'h7fef; 
        10'b0011101010: data <= 15'h7fec; 
        10'b0011101011: data <= 15'h7fd8; 
        10'b0011101100: data <= 15'h7ffd; 
        10'b0011101101: data <= 15'h0038; 
        10'b0011101110: data <= 15'h00a5; 
        10'b0011101111: data <= 15'h005b; 
        10'b0011110000: data <= 15'h005c; 
        10'b0011110001: data <= 15'h0013; 
        10'b0011110010: data <= 15'h0007; 
        10'b0011110011: data <= 15'h0005; 
        10'b0011110100: data <= 15'h7fe2; 
        10'b0011110101: data <= 15'h0010; 
        10'b0011110110: data <= 15'h7fd9; 
        10'b0011110111: data <= 15'h7f9d; 
        10'b0011111000: data <= 15'h7fad; 
        10'b0011111001: data <= 15'h7fd8; 
        10'b0011111010: data <= 15'h7fef; 
        10'b0011111011: data <= 15'h0017; 
        10'b0011111100: data <= 15'h0007; 
        10'b0011111101: data <= 15'h0004; 
        10'b0011111110: data <= 15'h0002; 
        10'b0011111111: data <= 15'h7fd7; 
        10'b0100000000: data <= 15'h7fa6; 
        10'b0100000001: data <= 15'h7fbb; 
        10'b0100000010: data <= 15'h7fed; 
        10'b0100000011: data <= 15'h7fd9; 
        10'b0100000100: data <= 15'h7fe9; 
        10'b0100000101: data <= 15'h7ff5; 
        10'b0100000110: data <= 15'h002a; 
        10'b0100000111: data <= 15'h0019; 
        10'b0100001000: data <= 15'h0007; 
        10'b0100001001: data <= 15'h0044; 
        10'b0100001010: data <= 15'h0072; 
        10'b0100001011: data <= 15'h0065; 
        10'b0100001100: data <= 15'h7ffc; 
        10'b0100001101: data <= 15'h7fe3; 
        10'b0100001110: data <= 15'h0001; 
        10'b0100001111: data <= 15'h7fc3; 
        10'b0100010000: data <= 15'h7fe6; 
        10'b0100010001: data <= 15'h7fc0; 
        10'b0100010010: data <= 15'h7fbc; 
        10'b0100010011: data <= 15'h7fb7; 
        10'b0100010100: data <= 15'h7fcf; 
        10'b0100010101: data <= 15'h7fea; 
        10'b0100010110: data <= 15'h7ff0; 
        10'b0100010111: data <= 15'h0014; 
        10'b0100011000: data <= 15'h0004; 
        10'b0100011001: data <= 15'h7fff; 
        10'b0100011010: data <= 15'h7ff6; 
        10'b0100011011: data <= 15'h7ff0; 
        10'b0100011100: data <= 15'h7fbb; 
        10'b0100011101: data <= 15'h7fdc; 
        10'b0100011110: data <= 15'h0022; 
        10'b0100011111: data <= 15'h002c; 
        10'b0100100000: data <= 15'h005a; 
        10'b0100100001: data <= 15'h0059; 
        10'b0100100010: data <= 15'h004d; 
        10'b0100100011: data <= 15'h0073; 
        10'b0100100100: data <= 15'h003a; 
        10'b0100100101: data <= 15'h000e; 
        10'b0100100110: data <= 15'h000f; 
        10'b0100100111: data <= 15'h7fc6; 
        10'b0100101000: data <= 15'h7fdd; 
        10'b0100101001: data <= 15'h7ff9; 
        10'b0100101010: data <= 15'h0029; 
        10'b0100101011: data <= 15'h7fff; 
        10'b0100101100: data <= 15'h0021; 
        10'b0100101101: data <= 15'h7fec; 
        10'b0100101110: data <= 15'h7fd8; 
        10'b0100101111: data <= 15'h7fda; 
        10'b0100110000: data <= 15'h7fd0; 
        10'b0100110001: data <= 15'h7ff2; 
        10'b0100110010: data <= 15'h7fee; 
        10'b0100110011: data <= 15'h000b; 
        10'b0100110100: data <= 15'h7ffc; 
        10'b0100110101: data <= 15'h0005; 
        10'b0100110110: data <= 15'h7ff6; 
        10'b0100110111: data <= 15'h7ff9; 
        10'b0100111000: data <= 15'h7fed; 
        10'b0100111001: data <= 15'h0040; 
        10'b0100111010: data <= 15'h0093; 
        10'b0100111011: data <= 15'h006e; 
        10'b0100111100: data <= 15'h00ad; 
        10'b0100111101: data <= 15'h0045; 
        10'b0100111110: data <= 15'h0048; 
        10'b0100111111: data <= 15'h007b; 
        10'b0101000000: data <= 15'h7fd9; 
        10'b0101000001: data <= 15'h7fdf; 
        10'b0101000010: data <= 15'h7fee; 
        10'b0101000011: data <= 15'h0009; 
        10'b0101000100: data <= 15'h0030; 
        10'b0101000101: data <= 15'h00a7; 
        10'b0101000110: data <= 15'h004f; 
        10'b0101000111: data <= 15'h0050; 
        10'b0101001000: data <= 15'h0083; 
        10'b0101001001: data <= 15'h005f; 
        10'b0101001010: data <= 15'h0037; 
        10'b0101001011: data <= 15'h000b; 
        10'b0101001100: data <= 15'h7ff7; 
        10'b0101001101: data <= 15'h7fe9; 
        10'b0101001110: data <= 15'h7fff; 
        10'b0101001111: data <= 15'h0000; 
        10'b0101010000: data <= 15'h000a; 
        10'b0101010001: data <= 15'h0015; 
        10'b0101010010: data <= 15'h7ff1; 
        10'b0101010011: data <= 15'h7fe8; 
        10'b0101010100: data <= 15'h0036; 
        10'b0101010101: data <= 15'h008c; 
        10'b0101010110: data <= 15'h00a1; 
        10'b0101010111: data <= 15'h0060; 
        10'b0101011000: data <= 15'h0078; 
        10'b0101011001: data <= 15'h0092; 
        10'b0101011010: data <= 15'h005d; 
        10'b0101011011: data <= 15'h0001; 
        10'b0101011100: data <= 15'h7fa2; 
        10'b0101011101: data <= 15'h0051; 
        10'b0101011110: data <= 15'h00af; 
        10'b0101011111: data <= 15'h008b; 
        10'b0101100000: data <= 15'h0077; 
        10'b0101100001: data <= 15'h00b5; 
        10'b0101100010: data <= 15'h00b7; 
        10'b0101100011: data <= 15'h00be; 
        10'b0101100100: data <= 15'h00c3; 
        10'b0101100101: data <= 15'h0082; 
        10'b0101100110: data <= 15'h003f; 
        10'b0101100111: data <= 15'h0002; 
        10'b0101101000: data <= 15'h7fe3; 
        10'b0101101001: data <= 15'h0005; 
        10'b0101101010: data <= 15'h000b; 
        10'b0101101011: data <= 15'h000b; 
        10'b0101101100: data <= 15'h0018; 
        10'b0101101101: data <= 15'h000f; 
        10'b0101101110: data <= 15'h7fec; 
        10'b0101101111: data <= 15'h0008; 
        10'b0101110000: data <= 15'h0051; 
        10'b0101110001: data <= 15'h007a; 
        10'b0101110010: data <= 15'h0073; 
        10'b0101110011: data <= 15'h004c; 
        10'b0101110100: data <= 15'h005f; 
        10'b0101110101: data <= 15'h003d; 
        10'b0101110110: data <= 15'h0037; 
        10'b0101110111: data <= 15'h7fe4; 
        10'b0101111000: data <= 15'h7fcf; 
        10'b0101111001: data <= 15'h0080; 
        10'b0101111010: data <= 15'h00af; 
        10'b0101111011: data <= 15'h007f; 
        10'b0101111100: data <= 15'h0092; 
        10'b0101111101: data <= 15'h0083; 
        10'b0101111110: data <= 15'h00b4; 
        10'b0101111111: data <= 15'h00b7; 
        10'b0110000000: data <= 15'h008f; 
        10'b0110000001: data <= 15'h0054; 
        10'b0110000010: data <= 15'h0005; 
        10'b0110000011: data <= 15'h7fc7; 
        10'b0110000100: data <= 15'h7fdf; 
        10'b0110000101: data <= 15'h7ff6; 
        10'b0110000110: data <= 15'h000b; 
        10'b0110000111: data <= 15'h000b; 
        10'b0110001000: data <= 15'h0005; 
        10'b0110001001: data <= 15'h0002; 
        10'b0110001010: data <= 15'h0011; 
        10'b0110001011: data <= 15'h000b; 
        10'b0110001100: data <= 15'h0025; 
        10'b0110001101: data <= 15'h0023; 
        10'b0110001110: data <= 15'h005f; 
        10'b0110001111: data <= 15'h0043; 
        10'b0110010000: data <= 15'h0020; 
        10'b0110010001: data <= 15'h0000; 
        10'b0110010010: data <= 15'h000c; 
        10'b0110010011: data <= 15'h7ffa; 
        10'b0110010100: data <= 15'h7fdc; 
        10'b0110010101: data <= 15'h0029; 
        10'b0110010110: data <= 15'h0018; 
        10'b0110010111: data <= 15'h0070; 
        10'b0110011000: data <= 15'h0077; 
        10'b0110011001: data <= 15'h0077; 
        10'b0110011010: data <= 15'h0051; 
        10'b0110011011: data <= 15'h0034; 
        10'b0110011100: data <= 15'h0041; 
        10'b0110011101: data <= 15'h0001; 
        10'b0110011110: data <= 15'h7fbe; 
        10'b0110011111: data <= 15'h7fa1; 
        10'b0110100000: data <= 15'h7fd9; 
        10'b0110100001: data <= 15'h0007; 
        10'b0110100010: data <= 15'h0004; 
        10'b0110100011: data <= 15'h0004; 
        10'b0110100100: data <= 15'h0012; 
        10'b0110100101: data <= 15'h0011; 
        10'b0110100110: data <= 15'h000b; 
        10'b0110100111: data <= 15'h7ff3; 
        10'b0110101000: data <= 15'h0003; 
        10'b0110101001: data <= 15'h002a; 
        10'b0110101010: data <= 15'h0029; 
        10'b0110101011: data <= 15'h001b; 
        10'b0110101100: data <= 15'h001b; 
        10'b0110101101: data <= 15'h7fce; 
        10'b0110101110: data <= 15'h7fe9; 
        10'b0110101111: data <= 15'h7fe8; 
        10'b0110110000: data <= 15'h7fdd; 
        10'b0110110001: data <= 15'h7fe5; 
        10'b0110110010: data <= 15'h7fdf; 
        10'b0110110011: data <= 15'h007a; 
        10'b0110110100: data <= 15'h00b3; 
        10'b0110110101: data <= 15'h00ac; 
        10'b0110110110: data <= 15'h0056; 
        10'b0110110111: data <= 15'h0008; 
        10'b0110111000: data <= 15'h7fdb; 
        10'b0110111001: data <= 15'h7f9e; 
        10'b0110111010: data <= 15'h7f85; 
        10'b0110111011: data <= 15'h7fa8; 
        10'b0110111100: data <= 15'h7fd9; 
        10'b0110111101: data <= 15'h0001; 
        10'b0110111110: data <= 15'h000a; 
        10'b0110111111: data <= 15'h7fff; 
        10'b0111000000: data <= 15'h0015; 
        10'b0111000001: data <= 15'h0002; 
        10'b0111000010: data <= 15'h7ff1; 
        10'b0111000011: data <= 15'h7ffc; 
        10'b0111000100: data <= 15'h0001; 
        10'b0111000101: data <= 15'h000d; 
        10'b0111000110: data <= 15'h7fdf; 
        10'b0111000111: data <= 15'h001a; 
        10'b0111001000: data <= 15'h004a; 
        10'b0111001001: data <= 15'h7fef; 
        10'b0111001010: data <= 15'h002a; 
        10'b0111001011: data <= 15'h003b; 
        10'b0111001100: data <= 15'h7ff8; 
        10'b0111001101: data <= 15'h7fbd; 
        10'b0111001110: data <= 15'h7ff5; 
        10'b0111001111: data <= 15'h0044; 
        10'b0111010000: data <= 15'h007a; 
        10'b0111010001: data <= 15'h0079; 
        10'b0111010010: data <= 15'h001e; 
        10'b0111010011: data <= 15'h7fbb; 
        10'b0111010100: data <= 15'h7f8d; 
        10'b0111010101: data <= 15'h7f62; 
        10'b0111010110: data <= 15'h7f91; 
        10'b0111010111: data <= 15'h7fa6; 
        10'b0111011000: data <= 15'h7fc4; 
        10'b0111011001: data <= 15'h0002; 
        10'b0111011010: data <= 15'h7ff3; 
        10'b0111011011: data <= 15'h000b; 
        10'b0111011100: data <= 15'h0007; 
        10'b0111011101: data <= 15'h7ffb; 
        10'b0111011110: data <= 15'h7ff0; 
        10'b0111011111: data <= 15'h7fe8; 
        10'b0111100000: data <= 15'h7fd3; 
        10'b0111100001: data <= 15'h7fc9; 
        10'b0111100010: data <= 15'h7fd3; 
        10'b0111100011: data <= 15'h0014; 
        10'b0111100100: data <= 15'h0028; 
        10'b0111100101: data <= 15'h002d; 
        10'b0111100110: data <= 15'h0045; 
        10'b0111100111: data <= 15'h0064; 
        10'b0111101000: data <= 15'h003d; 
        10'b0111101001: data <= 15'h001c; 
        10'b0111101010: data <= 15'h0027; 
        10'b0111101011: data <= 15'h0064; 
        10'b0111101100: data <= 15'h001e; 
        10'b0111101101: data <= 15'h7fec; 
        10'b0111101110: data <= 15'h7fd4; 
        10'b0111101111: data <= 15'h7f9b; 
        10'b0111110000: data <= 15'h7f9c; 
        10'b0111110001: data <= 15'h7f94; 
        10'b0111110010: data <= 15'h7f9b; 
        10'b0111110011: data <= 15'h7fb6; 
        10'b0111110100: data <= 15'h7fca; 
        10'b0111110101: data <= 15'h0005; 
        10'b0111110110: data <= 15'h0006; 
        10'b0111110111: data <= 15'h7ffb; 
        10'b0111111000: data <= 15'h0013; 
        10'b0111111001: data <= 15'h0000; 
        10'b0111111010: data <= 15'h7ff5; 
        10'b0111111011: data <= 15'h7ffb; 
        10'b0111111100: data <= 15'h7fd8; 
        10'b0111111101: data <= 15'h7fa5; 
        10'b0111111110: data <= 15'h7fa3; 
        10'b0111111111: data <= 15'h7fa5; 
        10'b1000000000: data <= 15'h7fda; 
        10'b1000000001: data <= 15'h000f; 
        10'b1000000010: data <= 15'h006e; 
        10'b1000000011: data <= 15'h0059; 
        10'b1000000100: data <= 15'h7fca; 
        10'b1000000101: data <= 15'h7fc9; 
        10'b1000000110: data <= 15'h0003; 
        10'b1000000111: data <= 15'h0042; 
        10'b1000001000: data <= 15'h7fd8; 
        10'b1000001001: data <= 15'h7fd2; 
        10'b1000001010: data <= 15'h7faa; 
        10'b1000001011: data <= 15'h7fcc; 
        10'b1000001100: data <= 15'h7fcf; 
        10'b1000001101: data <= 15'h7fb4; 
        10'b1000001110: data <= 15'h7fb0; 
        10'b1000001111: data <= 15'h7fac; 
        10'b1000010000: data <= 15'h7fc5; 
        10'b1000010001: data <= 15'h7ff7; 
        10'b1000010010: data <= 15'h0001; 
        10'b1000010011: data <= 15'h0012; 
        10'b1000010100: data <= 15'h000d; 
        10'b1000010101: data <= 15'h0019; 
        10'b1000010110: data <= 15'h0004; 
        10'b1000010111: data <= 15'h7fea; 
        10'b1000011000: data <= 15'h7fdc; 
        10'b1000011001: data <= 15'h7fc0; 
        10'b1000011010: data <= 15'h7f9a; 
        10'b1000011011: data <= 15'h7f98; 
        10'b1000011100: data <= 15'h7f94; 
        10'b1000011101: data <= 15'h7f95; 
        10'b1000011110: data <= 15'h7f88; 
        10'b1000011111: data <= 15'h7f9b; 
        10'b1000100000: data <= 15'h7f7d; 
        10'b1000100001: data <= 15'h7fa4; 
        10'b1000100010: data <= 15'h7fb3; 
        10'b1000100011: data <= 15'h7fa8; 
        10'b1000100100: data <= 15'h7fb4; 
        10'b1000100101: data <= 15'h7fe7; 
        10'b1000100110: data <= 15'h7fc6; 
        10'b1000100111: data <= 15'h7ff0; 
        10'b1000101000: data <= 15'h7fd9; 
        10'b1000101001: data <= 15'h7fd2; 
        10'b1000101010: data <= 15'h7fd5; 
        10'b1000101011: data <= 15'h7fda; 
        10'b1000101100: data <= 15'h7fe8; 
        10'b1000101101: data <= 15'h0007; 
        10'b1000101110: data <= 15'h7ff8; 
        10'b1000101111: data <= 15'h0003; 
        10'b1000110000: data <= 15'h7ffb; 
        10'b1000110001: data <= 15'h0004; 
        10'b1000110010: data <= 15'h000b; 
        10'b1000110011: data <= 15'h0001; 
        10'b1000110100: data <= 15'h7fda; 
        10'b1000110101: data <= 15'h7fc2; 
        10'b1000110110: data <= 15'h7fa2; 
        10'b1000110111: data <= 15'h7f6c; 
        10'b1000111000: data <= 15'h7f57; 
        10'b1000111001: data <= 15'h7f42; 
        10'b1000111010: data <= 15'h7eff; 
        10'b1000111011: data <= 15'h7f3c; 
        10'b1000111100: data <= 15'h7f41; 
        10'b1000111101: data <= 15'h7fc1; 
        10'b1000111110: data <= 15'h7fa8; 
        10'b1000111111: data <= 15'h7fd7; 
        10'b1001000000: data <= 15'h7fcf; 
        10'b1001000001: data <= 15'h7ff3; 
        10'b1001000010: data <= 15'h7fac; 
        10'b1001000011: data <= 15'h7fe4; 
        10'b1001000100: data <= 15'h7fdf; 
        10'b1001000101: data <= 15'h7fca; 
        10'b1001000110: data <= 15'h7ff1; 
        10'b1001000111: data <= 15'h7fe6; 
        10'b1001001000: data <= 15'h0003; 
        10'b1001001001: data <= 15'h0015; 
        10'b1001001010: data <= 15'h000d; 
        10'b1001001011: data <= 15'h0004; 
        10'b1001001100: data <= 15'h0002; 
        10'b1001001101: data <= 15'h0000; 
        10'b1001001110: data <= 15'h0015; 
        10'b1001001111: data <= 15'h7fe9; 
        10'b1001010000: data <= 15'h7fe7; 
        10'b1001010001: data <= 15'h7fc3; 
        10'b1001010010: data <= 15'h7faa; 
        10'b1001010011: data <= 15'h7f7b; 
        10'b1001010100: data <= 15'h7f68; 
        10'b1001010101: data <= 15'h7f59; 
        10'b1001010110: data <= 15'h7f51; 
        10'b1001010111: data <= 15'h7f63; 
        10'b1001011000: data <= 15'h7f9c; 
        10'b1001011001: data <= 15'h7f9d; 
        10'b1001011010: data <= 15'h7f9c; 
        10'b1001011011: data <= 15'h7fc6; 
        10'b1001011100: data <= 15'h7fc2; 
        10'b1001011101: data <= 15'h7fa2; 
        10'b1001011110: data <= 15'h7f8f; 
        10'b1001011111: data <= 15'h7fd0; 
        10'b1001100000: data <= 15'h7fe5; 
        10'b1001100001: data <= 15'h7ff1; 
        10'b1001100010: data <= 15'h0008; 
        10'b1001100011: data <= 15'h7ffe; 
        10'b1001100100: data <= 15'h000a; 
        10'b1001100101: data <= 15'h000d; 
        10'b1001100110: data <= 15'h0001; 
        10'b1001100111: data <= 15'h0002; 
        10'b1001101000: data <= 15'h0010; 
        10'b1001101001: data <= 15'h0004; 
        10'b1001101010: data <= 15'h0005; 
        10'b1001101011: data <= 15'h0010; 
        10'b1001101100: data <= 15'h7ff6; 
        10'b1001101101: data <= 15'h7fcf; 
        10'b1001101110: data <= 15'h7fb1; 
        10'b1001101111: data <= 15'h7f94; 
        10'b1001110000: data <= 15'h7fb0; 
        10'b1001110001: data <= 15'h7fac; 
        10'b1001110010: data <= 15'h7fa5; 
        10'b1001110011: data <= 15'h7fc2; 
        10'b1001110100: data <= 15'h7fbb; 
        10'b1001110101: data <= 15'h7fa4; 
        10'b1001110110: data <= 15'h7fb2; 
        10'b1001110111: data <= 15'h7f93; 
        10'b1001111000: data <= 15'h7f88; 
        10'b1001111001: data <= 15'h7f8a; 
        10'b1001111010: data <= 15'h7f9e; 
        10'b1001111011: data <= 15'h7fa9; 
        10'b1001111100: data <= 15'h7fe8; 
        10'b1001111101: data <= 15'h001d; 
        10'b1001111110: data <= 15'h0010; 
        10'b1001111111: data <= 15'h0014; 
        10'b1010000000: data <= 15'h0021; 
        10'b1010000001: data <= 15'h0007; 
        10'b1010000010: data <= 15'h0008; 
        10'b1010000011: data <= 15'h000c; 
        10'b1010000100: data <= 15'h0013; 
        10'b1010000101: data <= 15'h000f; 
        10'b1010000110: data <= 15'h0006; 
        10'b1010000111: data <= 15'h7ff8; 
        10'b1010001000: data <= 15'h7ff2; 
        10'b1010001001: data <= 15'h7fd5; 
        10'b1010001010: data <= 15'h7fcf; 
        10'b1010001011: data <= 15'h7fbf; 
        10'b1010001100: data <= 15'h7ffb; 
        10'b1010001101: data <= 15'h7fe6; 
        10'b1010001110: data <= 15'h7feb; 
        10'b1010001111: data <= 15'h7fb1; 
        10'b1010010000: data <= 15'h7fbf; 
        10'b1010010001: data <= 15'h7faf; 
        10'b1010010010: data <= 15'h7fbb; 
        10'b1010010011: data <= 15'h7f8a; 
        10'b1010010100: data <= 15'h7f81; 
        10'b1010010101: data <= 15'h7f90; 
        10'b1010010110: data <= 15'h7fba; 
        10'b1010010111: data <= 15'h7ff9; 
        10'b1010011000: data <= 15'h001b; 
        10'b1010011001: data <= 15'h003f; 
        10'b1010011010: data <= 15'h005b; 
        10'b1010011011: data <= 15'h004c; 
        10'b1010011100: data <= 15'h0024; 
        10'b1010011101: data <= 15'h7ffe; 
        10'b1010011110: data <= 15'h001a; 
        10'b1010011111: data <= 15'h7ffd; 
        10'b1010100000: data <= 15'h0000; 
        10'b1010100001: data <= 15'h7ff6; 
        10'b1010100010: data <= 15'h7ffd; 
        10'b1010100011: data <= 15'h0016; 
        10'b1010100100: data <= 15'h0010; 
        10'b1010100101: data <= 15'h0018; 
        10'b1010100110: data <= 15'h0012; 
        10'b1010100111: data <= 15'h001a; 
        10'b1010101000: data <= 15'h0024; 
        10'b1010101001: data <= 15'h0014; 
        10'b1010101010: data <= 15'h7ff3; 
        10'b1010101011: data <= 15'h7fd7; 
        10'b1010101100: data <= 15'h7ffd; 
        10'b1010101101: data <= 15'h7fc2; 
        10'b1010101110: data <= 15'h7fb1; 
        10'b1010101111: data <= 15'h7fad; 
        10'b1010110000: data <= 15'h7fda; 
        10'b1010110001: data <= 15'h001b; 
        10'b1010110010: data <= 15'h002f; 
        10'b1010110011: data <= 15'h0030; 
        10'b1010110100: data <= 15'h006e; 
        10'b1010110101: data <= 15'h0077; 
        10'b1010110110: data <= 15'h0044; 
        10'b1010110111: data <= 15'h002a; 
        10'b1010111000: data <= 15'h0021; 
        10'b1010111001: data <= 15'h7ffa; 
        10'b1010111010: data <= 15'h000f; 
        10'b1010111011: data <= 15'h7fff; 
        10'b1010111100: data <= 15'h0005; 
        10'b1010111101: data <= 15'h0015; 
        10'b1010111110: data <= 15'h0015; 
        10'b1010111111: data <= 15'h7ffe; 
        10'b1011000000: data <= 15'h0002; 
        10'b1011000001: data <= 15'h0025; 
        10'b1011000010: data <= 15'h001c; 
        10'b1011000011: data <= 15'h0050; 
        10'b1011000100: data <= 15'h0058; 
        10'b1011000101: data <= 15'h0059; 
        10'b1011000110: data <= 15'h004d; 
        10'b1011000111: data <= 15'h001f; 
        10'b1011001000: data <= 15'h0051; 
        10'b1011001001: data <= 15'h0049; 
        10'b1011001010: data <= 15'h0046; 
        10'b1011001011: data <= 15'h0041; 
        10'b1011001100: data <= 15'h007a; 
        10'b1011001101: data <= 15'h0085; 
        10'b1011001110: data <= 15'h0092; 
        10'b1011001111: data <= 15'h0098; 
        10'b1011010000: data <= 15'h00aa; 
        10'b1011010001: data <= 15'h0079; 
        10'b1011010010: data <= 15'h002f; 
        10'b1011010011: data <= 15'h0016; 
        10'b1011010100: data <= 15'h7ffd; 
        10'b1011010101: data <= 15'h7ffe; 
        10'b1011010110: data <= 15'h0006; 
        10'b1011010111: data <= 15'h0005; 
        10'b1011011000: data <= 15'h0001; 
        10'b1011011001: data <= 15'h0014; 
        10'b1011011010: data <= 15'h0005; 
        10'b1011011011: data <= 15'h7ff9; 
        10'b1011011100: data <= 15'h0014; 
        10'b1011011101: data <= 15'h001e; 
        10'b1011011110: data <= 15'h002b; 
        10'b1011011111: data <= 15'h003b; 
        10'b1011100000: data <= 15'h0043; 
        10'b1011100001: data <= 15'h0066; 
        10'b1011100010: data <= 15'h006a; 
        10'b1011100011: data <= 15'h0077; 
        10'b1011100100: data <= 15'h008c; 
        10'b1011100101: data <= 15'h008e; 
        10'b1011100110: data <= 15'h00ad; 
        10'b1011100111: data <= 15'h0064; 
        10'b1011101000: data <= 15'h0045; 
        10'b1011101001: data <= 15'h003a; 
        10'b1011101010: data <= 15'h0055; 
        10'b1011101011: data <= 15'h005c; 
        10'b1011101100: data <= 15'h0043; 
        10'b1011101101: data <= 15'h002f; 
        10'b1011101110: data <= 15'h0013; 
        10'b1011101111: data <= 15'h0007; 
        10'b1011110000: data <= 15'h0004; 
        10'b1011110001: data <= 15'h0008; 
        10'b1011110010: data <= 15'h7ff9; 
        10'b1011110011: data <= 15'h0004; 
        10'b1011110100: data <= 15'h7ffb; 
        10'b1011110101: data <= 15'h0009; 
        10'b1011110110: data <= 15'h7ff8; 
        10'b1011110111: data <= 15'h0018; 
        10'b1011111000: data <= 15'h000e; 
        10'b1011111001: data <= 15'h0008; 
        10'b1011111010: data <= 15'h7ffd; 
        10'b1011111011: data <= 15'h0017; 
        10'b1011111100: data <= 15'h0013; 
        10'b1011111101: data <= 15'h000d; 
        10'b1011111110: data <= 15'h7ffc; 
        10'b1011111111: data <= 15'h7ffb; 
        10'b1100000000: data <= 15'h0005; 
        10'b1100000001: data <= 15'h7ffc; 
        10'b1100000010: data <= 15'h0005; 
        10'b1100000011: data <= 15'h000f; 
        10'b1100000100: data <= 15'h0001; 
        10'b1100000101: data <= 15'h0008; 
        10'b1100000110: data <= 15'h001a; 
        10'b1100000111: data <= 15'h0017; 
        10'b1100001000: data <= 15'h000d; 
        10'b1100001001: data <= 15'h0008; 
        10'b1100001010: data <= 15'h7ff9; 
        10'b1100001011: data <= 15'h001a; 
        10'b1100001100: data <= 15'h000e; 
        10'b1100001101: data <= 15'h7ffb; 
        10'b1100001110: data <= 15'h0002; 
        10'b1100001111: data <= 15'h7ffd; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 10) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 16'h0024; 
        10'b0000000001: data <= 16'h0020; 
        10'b0000000010: data <= 16'hfff6; 
        10'b0000000011: data <= 16'h0016; 
        10'b0000000100: data <= 16'h0014; 
        10'b0000000101: data <= 16'h0021; 
        10'b0000000110: data <= 16'hfff4; 
        10'b0000000111: data <= 16'h0006; 
        10'b0000001000: data <= 16'h0026; 
        10'b0000001001: data <= 16'hfff0; 
        10'b0000001010: data <= 16'hfffb; 
        10'b0000001011: data <= 16'h0011; 
        10'b0000001100: data <= 16'h0030; 
        10'b0000001101: data <= 16'h001f; 
        10'b0000001110: data <= 16'hffec; 
        10'b0000001111: data <= 16'hfff7; 
        10'b0000010000: data <= 16'hfff6; 
        10'b0000010001: data <= 16'h0013; 
        10'b0000010010: data <= 16'h0023; 
        10'b0000010011: data <= 16'h0003; 
        10'b0000010100: data <= 16'h0003; 
        10'b0000010101: data <= 16'hfffd; 
        10'b0000010110: data <= 16'hfff1; 
        10'b0000010111: data <= 16'h0005; 
        10'b0000011000: data <= 16'h0027; 
        10'b0000011001: data <= 16'h000c; 
        10'b0000011010: data <= 16'hffee; 
        10'b0000011011: data <= 16'h0013; 
        10'b0000011100: data <= 16'h0020; 
        10'b0000011101: data <= 16'h001b; 
        10'b0000011110: data <= 16'h000d; 
        10'b0000011111: data <= 16'hfff8; 
        10'b0000100000: data <= 16'hffed; 
        10'b0000100001: data <= 16'hfff1; 
        10'b0000100010: data <= 16'hfffd; 
        10'b0000100011: data <= 16'h0031; 
        10'b0000100100: data <= 16'hffee; 
        10'b0000100101: data <= 16'h0027; 
        10'b0000100110: data <= 16'h000f; 
        10'b0000100111: data <= 16'h0018; 
        10'b0000101000: data <= 16'h0013; 
        10'b0000101001: data <= 16'h001c; 
        10'b0000101010: data <= 16'h0001; 
        10'b0000101011: data <= 16'hffeb; 
        10'b0000101100: data <= 16'hfff5; 
        10'b0000101101: data <= 16'h001e; 
        10'b0000101110: data <= 16'hffff; 
        10'b0000101111: data <= 16'h0009; 
        10'b0000110000: data <= 16'h0026; 
        10'b0000110001: data <= 16'hfffd; 
        10'b0000110010: data <= 16'h0007; 
        10'b0000110011: data <= 16'h0003; 
        10'b0000110100: data <= 16'h0015; 
        10'b0000110101: data <= 16'h0029; 
        10'b0000110110: data <= 16'h0000; 
        10'b0000110111: data <= 16'h0009; 
        10'b0000111000: data <= 16'h002b; 
        10'b0000111001: data <= 16'h002c; 
        10'b0000111010: data <= 16'h0003; 
        10'b0000111011: data <= 16'h001e; 
        10'b0000111100: data <= 16'h0024; 
        10'b0000111101: data <= 16'hfffe; 
        10'b0000111110: data <= 16'hfffc; 
        10'b0000111111: data <= 16'h000d; 
        10'b0001000000: data <= 16'h0024; 
        10'b0001000001: data <= 16'hfffb; 
        10'b0001000010: data <= 16'hfff5; 
        10'b0001000011: data <= 16'h001c; 
        10'b0001000100: data <= 16'h0010; 
        10'b0001000101: data <= 16'h0023; 
        10'b0001000110: data <= 16'hffeb; 
        10'b0001000111: data <= 16'h0025; 
        10'b0001001000: data <= 16'hfff3; 
        10'b0001001001: data <= 16'hfff2; 
        10'b0001001010: data <= 16'h0003; 
        10'b0001001011: data <= 16'hffee; 
        10'b0001001100: data <= 16'h002a; 
        10'b0001001101: data <= 16'hfff5; 
        10'b0001001110: data <= 16'hfff1; 
        10'b0001001111: data <= 16'h002a; 
        10'b0001010000: data <= 16'h0008; 
        10'b0001010001: data <= 16'h0007; 
        10'b0001010010: data <= 16'h0009; 
        10'b0001010011: data <= 16'h0013; 
        10'b0001010100: data <= 16'h0034; 
        10'b0001010101: data <= 16'h0002; 
        10'b0001010110: data <= 16'hfffb; 
        10'b0001010111: data <= 16'h000f; 
        10'b0001011000: data <= 16'h0010; 
        10'b0001011001: data <= 16'hffef; 
        10'b0001011010: data <= 16'h002b; 
        10'b0001011011: data <= 16'h0017; 
        10'b0001011100: data <= 16'hfff8; 
        10'b0001011101: data <= 16'h002b; 
        10'b0001011110: data <= 16'h000e; 
        10'b0001011111: data <= 16'h0022; 
        10'b0001100000: data <= 16'hfffc; 
        10'b0001100001: data <= 16'hffd9; 
        10'b0001100010: data <= 16'hfffc; 
        10'b0001100011: data <= 16'hffc5; 
        10'b0001100100: data <= 16'hfff9; 
        10'b0001100101: data <= 16'hffe1; 
        10'b0001100110: data <= 16'h000a; 
        10'b0001100111: data <= 16'h0006; 
        10'b0001101000: data <= 16'h000d; 
        10'b0001101001: data <= 16'hfffd; 
        10'b0001101010: data <= 16'h0022; 
        10'b0001101011: data <= 16'hfffc; 
        10'b0001101100: data <= 16'hfffb; 
        10'b0001101101: data <= 16'h002f; 
        10'b0001101110: data <= 16'h0011; 
        10'b0001101111: data <= 16'h001e; 
        10'b0001110000: data <= 16'h0006; 
        10'b0001110001: data <= 16'h000a; 
        10'b0001110010: data <= 16'h0002; 
        10'b0001110011: data <= 16'hfff6; 
        10'b0001110100: data <= 16'hffef; 
        10'b0001110101: data <= 16'h001e; 
        10'b0001110110: data <= 16'h0015; 
        10'b0001110111: data <= 16'hfffc; 
        10'b0001111000: data <= 16'hffe5; 
        10'b0001111001: data <= 16'h000a; 
        10'b0001111010: data <= 16'hffd4; 
        10'b0001111011: data <= 16'hffc2; 
        10'b0001111100: data <= 16'hffa9; 
        10'b0001111101: data <= 16'hff63; 
        10'b0001111110: data <= 16'hff38; 
        10'b0001111111: data <= 16'hfef4; 
        10'b0010000000: data <= 16'hff3a; 
        10'b0010000001: data <= 16'hff39; 
        10'b0010000010: data <= 16'hff6c; 
        10'b0010000011: data <= 16'hffbf; 
        10'b0010000100: data <= 16'hffe2; 
        10'b0010000101: data <= 16'hffea; 
        10'b0010000110: data <= 16'h0007; 
        10'b0010000111: data <= 16'h0025; 
        10'b0010001000: data <= 16'h001d; 
        10'b0010001001: data <= 16'h001b; 
        10'b0010001010: data <= 16'h0000; 
        10'b0010001011: data <= 16'h0001; 
        10'b0010001100: data <= 16'h0024; 
        10'b0010001101: data <= 16'h001a; 
        10'b0010001110: data <= 16'h001e; 
        10'b0010001111: data <= 16'h0013; 
        10'b0010010000: data <= 16'h0017; 
        10'b0010010001: data <= 16'hffe3; 
        10'b0010010010: data <= 16'hffe7; 
        10'b0010010011: data <= 16'hffe4; 
        10'b0010010100: data <= 16'hffa5; 
        10'b0010010101: data <= 16'hffa7; 
        10'b0010010110: data <= 16'hffa0; 
        10'b0010010111: data <= 16'hff81; 
        10'b0010011000: data <= 16'hff61; 
        10'b0010011001: data <= 16'hff44; 
        10'b0010011010: data <= 16'hfee1; 
        10'b0010011011: data <= 16'hfeca; 
        10'b0010011100: data <= 16'hfe79; 
        10'b0010011101: data <= 16'hfefe; 
        10'b0010011110: data <= 16'hff5d; 
        10'b0010011111: data <= 16'hffb1; 
        10'b0010100000: data <= 16'hffad; 
        10'b0010100001: data <= 16'hff94; 
        10'b0010100010: data <= 16'hff9b; 
        10'b0010100011: data <= 16'hffb8; 
        10'b0010100100: data <= 16'hffe3; 
        10'b0010100101: data <= 16'hfff3; 
        10'b0010100110: data <= 16'h0004; 
        10'b0010100111: data <= 16'h0019; 
        10'b0010101000: data <= 16'h0021; 
        10'b0010101001: data <= 16'h0021; 
        10'b0010101010: data <= 16'hffeb; 
        10'b0010101011: data <= 16'h0022; 
        10'b0010101100: data <= 16'h0015; 
        10'b0010101101: data <= 16'hff9f; 
        10'b0010101110: data <= 16'hff8a; 
        10'b0010101111: data <= 16'hff75; 
        10'b0010110000: data <= 16'hff64; 
        10'b0010110001: data <= 16'hff40; 
        10'b0010110010: data <= 16'hff73; 
        10'b0010110011: data <= 16'hffd3; 
        10'b0010110100: data <= 16'h000b; 
        10'b0010110101: data <= 16'h00ad; 
        10'b0010110110: data <= 16'h0102; 
        10'b0010110111: data <= 16'h00cd; 
        10'b0010111000: data <= 16'h0090; 
        10'b0010111001: data <= 16'h0078; 
        10'b0010111010: data <= 16'h0098; 
        10'b0010111011: data <= 16'hffe6; 
        10'b0010111100: data <= 16'hffdb; 
        10'b0010111101: data <= 16'hff8d; 
        10'b0010111110: data <= 16'hff31; 
        10'b0010111111: data <= 16'hff3f; 
        10'b0011000000: data <= 16'hff92; 
        10'b0011000001: data <= 16'hffca; 
        10'b0011000010: data <= 16'hfff8; 
        10'b0011000011: data <= 16'h0011; 
        10'b0011000100: data <= 16'h0032; 
        10'b0011000101: data <= 16'hfffe; 
        10'b0011000110: data <= 16'hfff0; 
        10'b0011000111: data <= 16'hffee; 
        10'b0011001000: data <= 16'hff91; 
        10'b0011001001: data <= 16'hff58; 
        10'b0011001010: data <= 16'hff3a; 
        10'b0011001011: data <= 16'hff14; 
        10'b0011001100: data <= 16'hff21; 
        10'b0011001101: data <= 16'hffb1; 
        10'b0011001110: data <= 16'hfffa; 
        10'b0011001111: data <= 16'h003d; 
        10'b0011010000: data <= 16'h00eb; 
        10'b0011010001: data <= 16'h0118; 
        10'b0011010010: data <= 16'h0180; 
        10'b0011010011: data <= 16'h0182; 
        10'b0011010100: data <= 16'h0192; 
        10'b0011010101: data <= 16'h00b6; 
        10'b0011010110: data <= 16'h0089; 
        10'b0011010111: data <= 16'h000f; 
        10'b0011011000: data <= 16'h0024; 
        10'b0011011001: data <= 16'h0028; 
        10'b0011011010: data <= 16'hff76; 
        10'b0011011011: data <= 16'hff08; 
        10'b0011011100: data <= 16'hff6e; 
        10'b0011011101: data <= 16'hffdc; 
        10'b0011011110: data <= 16'hffdb; 
        10'b0011011111: data <= 16'h0021; 
        10'b0011100000: data <= 16'h0030; 
        10'b0011100001: data <= 16'h0031; 
        10'b0011100010: data <= 16'h0019; 
        10'b0011100011: data <= 16'hfff1; 
        10'b0011100100: data <= 16'hff8d; 
        10'b0011100101: data <= 16'hff52; 
        10'b0011100110: data <= 16'hff35; 
        10'b0011100111: data <= 16'hfee4; 
        10'b0011101000: data <= 16'hffb5; 
        10'b0011101001: data <= 16'hffdd; 
        10'b0011101010: data <= 16'hffd8; 
        10'b0011101011: data <= 16'hffaf; 
        10'b0011101100: data <= 16'hfffa; 
        10'b0011101101: data <= 16'h0070; 
        10'b0011101110: data <= 16'h0149; 
        10'b0011101111: data <= 16'h00b6; 
        10'b0011110000: data <= 16'h00b9; 
        10'b0011110001: data <= 16'h0026; 
        10'b0011110010: data <= 16'h000f; 
        10'b0011110011: data <= 16'h000a; 
        10'b0011110100: data <= 16'hffc3; 
        10'b0011110101: data <= 16'h0020; 
        10'b0011110110: data <= 16'hffb2; 
        10'b0011110111: data <= 16'hff3a; 
        10'b0011111000: data <= 16'hff59; 
        10'b0011111001: data <= 16'hffb0; 
        10'b0011111010: data <= 16'hffdd; 
        10'b0011111011: data <= 16'h002d; 
        10'b0011111100: data <= 16'h000f; 
        10'b0011111101: data <= 16'h0009; 
        10'b0011111110: data <= 16'h0003; 
        10'b0011111111: data <= 16'hffae; 
        10'b0100000000: data <= 16'hff4d; 
        10'b0100000001: data <= 16'hff76; 
        10'b0100000010: data <= 16'hffd9; 
        10'b0100000011: data <= 16'hffb1; 
        10'b0100000100: data <= 16'hffd1; 
        10'b0100000101: data <= 16'hffeb; 
        10'b0100000110: data <= 16'h0054; 
        10'b0100000111: data <= 16'h0033; 
        10'b0100001000: data <= 16'h000f; 
        10'b0100001001: data <= 16'h0088; 
        10'b0100001010: data <= 16'h00e4; 
        10'b0100001011: data <= 16'h00cb; 
        10'b0100001100: data <= 16'hfff8; 
        10'b0100001101: data <= 16'hffc6; 
        10'b0100001110: data <= 16'h0002; 
        10'b0100001111: data <= 16'hff87; 
        10'b0100010000: data <= 16'hffcd; 
        10'b0100010001: data <= 16'hff81; 
        10'b0100010010: data <= 16'hff78; 
        10'b0100010011: data <= 16'hff6f; 
        10'b0100010100: data <= 16'hff9d; 
        10'b0100010101: data <= 16'hffd5; 
        10'b0100010110: data <= 16'hffe1; 
        10'b0100010111: data <= 16'h0028; 
        10'b0100011000: data <= 16'h0009; 
        10'b0100011001: data <= 16'hfffe; 
        10'b0100011010: data <= 16'hffed; 
        10'b0100011011: data <= 16'hffe0; 
        10'b0100011100: data <= 16'hff76; 
        10'b0100011101: data <= 16'hffb8; 
        10'b0100011110: data <= 16'h0043; 
        10'b0100011111: data <= 16'h0058; 
        10'b0100100000: data <= 16'h00b3; 
        10'b0100100001: data <= 16'h00b2; 
        10'b0100100010: data <= 16'h0099; 
        10'b0100100011: data <= 16'h00e7; 
        10'b0100100100: data <= 16'h0074; 
        10'b0100100101: data <= 16'h001b; 
        10'b0100100110: data <= 16'h001e; 
        10'b0100100111: data <= 16'hff8b; 
        10'b0100101000: data <= 16'hffba; 
        10'b0100101001: data <= 16'hfff2; 
        10'b0100101010: data <= 16'h0051; 
        10'b0100101011: data <= 16'hfffe; 
        10'b0100101100: data <= 16'h0041; 
        10'b0100101101: data <= 16'hffd9; 
        10'b0100101110: data <= 16'hffb0; 
        10'b0100101111: data <= 16'hffb4; 
        10'b0100110000: data <= 16'hffa0; 
        10'b0100110001: data <= 16'hffe5; 
        10'b0100110010: data <= 16'hffdc; 
        10'b0100110011: data <= 16'h0017; 
        10'b0100110100: data <= 16'hfff8; 
        10'b0100110101: data <= 16'h0009; 
        10'b0100110110: data <= 16'hffeb; 
        10'b0100110111: data <= 16'hfff3; 
        10'b0100111000: data <= 16'hffda; 
        10'b0100111001: data <= 16'h007f; 
        10'b0100111010: data <= 16'h0126; 
        10'b0100111011: data <= 16'h00dc; 
        10'b0100111100: data <= 16'h0159; 
        10'b0100111101: data <= 16'h008a; 
        10'b0100111110: data <= 16'h008f; 
        10'b0100111111: data <= 16'h00f6; 
        10'b0101000000: data <= 16'hffb2; 
        10'b0101000001: data <= 16'hffbd; 
        10'b0101000010: data <= 16'hffdc; 
        10'b0101000011: data <= 16'h0011; 
        10'b0101000100: data <= 16'h005f; 
        10'b0101000101: data <= 16'h014e; 
        10'b0101000110: data <= 16'h009e; 
        10'b0101000111: data <= 16'h00a0; 
        10'b0101001000: data <= 16'h0106; 
        10'b0101001001: data <= 16'h00be; 
        10'b0101001010: data <= 16'h006f; 
        10'b0101001011: data <= 16'h0017; 
        10'b0101001100: data <= 16'hffee; 
        10'b0101001101: data <= 16'hffd3; 
        10'b0101001110: data <= 16'hfffe; 
        10'b0101001111: data <= 16'h0000; 
        10'b0101010000: data <= 16'h0015; 
        10'b0101010001: data <= 16'h002b; 
        10'b0101010010: data <= 16'hffe2; 
        10'b0101010011: data <= 16'hffd1; 
        10'b0101010100: data <= 16'h006b; 
        10'b0101010101: data <= 16'h0117; 
        10'b0101010110: data <= 16'h0143; 
        10'b0101010111: data <= 16'h00c0; 
        10'b0101011000: data <= 16'h00ef; 
        10'b0101011001: data <= 16'h0125; 
        10'b0101011010: data <= 16'h00bb; 
        10'b0101011011: data <= 16'h0002; 
        10'b0101011100: data <= 16'hff44; 
        10'b0101011101: data <= 16'h00a2; 
        10'b0101011110: data <= 16'h015f; 
        10'b0101011111: data <= 16'h0116; 
        10'b0101100000: data <= 16'h00ed; 
        10'b0101100001: data <= 16'h016b; 
        10'b0101100010: data <= 16'h016e; 
        10'b0101100011: data <= 16'h017b; 
        10'b0101100100: data <= 16'h0186; 
        10'b0101100101: data <= 16'h0105; 
        10'b0101100110: data <= 16'h007d; 
        10'b0101100111: data <= 16'h0003; 
        10'b0101101000: data <= 16'hffc6; 
        10'b0101101001: data <= 16'h0009; 
        10'b0101101010: data <= 16'h0015; 
        10'b0101101011: data <= 16'h0017; 
        10'b0101101100: data <= 16'h0030; 
        10'b0101101101: data <= 16'h001e; 
        10'b0101101110: data <= 16'hffd7; 
        10'b0101101111: data <= 16'h000f; 
        10'b0101110000: data <= 16'h00a2; 
        10'b0101110001: data <= 16'h00f4; 
        10'b0101110010: data <= 16'h00e6; 
        10'b0101110011: data <= 16'h0097; 
        10'b0101110100: data <= 16'h00be; 
        10'b0101110101: data <= 16'h007a; 
        10'b0101110110: data <= 16'h006e; 
        10'b0101110111: data <= 16'hffc7; 
        10'b0101111000: data <= 16'hff9e; 
        10'b0101111001: data <= 16'h00ff; 
        10'b0101111010: data <= 16'h015e; 
        10'b0101111011: data <= 16'h00fe; 
        10'b0101111100: data <= 16'h0124; 
        10'b0101111101: data <= 16'h0106; 
        10'b0101111110: data <= 16'h0168; 
        10'b0101111111: data <= 16'h016e; 
        10'b0110000000: data <= 16'h011e; 
        10'b0110000001: data <= 16'h00a7; 
        10'b0110000010: data <= 16'h000a; 
        10'b0110000011: data <= 16'hff8e; 
        10'b0110000100: data <= 16'hffbe; 
        10'b0110000101: data <= 16'hffeb; 
        10'b0110000110: data <= 16'h0016; 
        10'b0110000111: data <= 16'h0016; 
        10'b0110001000: data <= 16'h000a; 
        10'b0110001001: data <= 16'h0005; 
        10'b0110001010: data <= 16'h0021; 
        10'b0110001011: data <= 16'h0015; 
        10'b0110001100: data <= 16'h004a; 
        10'b0110001101: data <= 16'h0046; 
        10'b0110001110: data <= 16'h00bf; 
        10'b0110001111: data <= 16'h0085; 
        10'b0110010000: data <= 16'h0041; 
        10'b0110010001: data <= 16'hffff; 
        10'b0110010010: data <= 16'h0018; 
        10'b0110010011: data <= 16'hfff4; 
        10'b0110010100: data <= 16'hffb8; 
        10'b0110010101: data <= 16'h0053; 
        10'b0110010110: data <= 16'h002f; 
        10'b0110010111: data <= 16'h00e0; 
        10'b0110011000: data <= 16'h00ee; 
        10'b0110011001: data <= 16'h00ee; 
        10'b0110011010: data <= 16'h00a2; 
        10'b0110011011: data <= 16'h0068; 
        10'b0110011100: data <= 16'h0082; 
        10'b0110011101: data <= 16'h0002; 
        10'b0110011110: data <= 16'hff7d; 
        10'b0110011111: data <= 16'hff41; 
        10'b0110100000: data <= 16'hffb1; 
        10'b0110100001: data <= 16'h000d; 
        10'b0110100010: data <= 16'h0007; 
        10'b0110100011: data <= 16'h0009; 
        10'b0110100100: data <= 16'h0025; 
        10'b0110100101: data <= 16'h0021; 
        10'b0110100110: data <= 16'h0016; 
        10'b0110100111: data <= 16'hffe5; 
        10'b0110101000: data <= 16'h0005; 
        10'b0110101001: data <= 16'h0055; 
        10'b0110101010: data <= 16'h0051; 
        10'b0110101011: data <= 16'h0036; 
        10'b0110101100: data <= 16'h0037; 
        10'b0110101101: data <= 16'hff9b; 
        10'b0110101110: data <= 16'hffd1; 
        10'b0110101111: data <= 16'hffd1; 
        10'b0110110000: data <= 16'hffba; 
        10'b0110110001: data <= 16'hffca; 
        10'b0110110010: data <= 16'hffbe; 
        10'b0110110011: data <= 16'h00f5; 
        10'b0110110100: data <= 16'h0166; 
        10'b0110110101: data <= 16'h0157; 
        10'b0110110110: data <= 16'h00ac; 
        10'b0110110111: data <= 16'h0011; 
        10'b0110111000: data <= 16'hffb5; 
        10'b0110111001: data <= 16'hff3b; 
        10'b0110111010: data <= 16'hff0a; 
        10'b0110111011: data <= 16'hff51; 
        10'b0110111100: data <= 16'hffb2; 
        10'b0110111101: data <= 16'h0001; 
        10'b0110111110: data <= 16'h0014; 
        10'b0110111111: data <= 16'hfffd; 
        10'b0111000000: data <= 16'h002a; 
        10'b0111000001: data <= 16'h0004; 
        10'b0111000010: data <= 16'hffe2; 
        10'b0111000011: data <= 16'hfff8; 
        10'b0111000100: data <= 16'h0003; 
        10'b0111000101: data <= 16'h0019; 
        10'b0111000110: data <= 16'hffbe; 
        10'b0111000111: data <= 16'h0034; 
        10'b0111001000: data <= 16'h0093; 
        10'b0111001001: data <= 16'hffde; 
        10'b0111001010: data <= 16'h0054; 
        10'b0111001011: data <= 16'h0076; 
        10'b0111001100: data <= 16'hfff0; 
        10'b0111001101: data <= 16'hff79; 
        10'b0111001110: data <= 16'hffe9; 
        10'b0111001111: data <= 16'h0088; 
        10'b0111010000: data <= 16'h00f4; 
        10'b0111010001: data <= 16'h00f3; 
        10'b0111010010: data <= 16'h003d; 
        10'b0111010011: data <= 16'hff76; 
        10'b0111010100: data <= 16'hff1b; 
        10'b0111010101: data <= 16'hfec3; 
        10'b0111010110: data <= 16'hff22; 
        10'b0111010111: data <= 16'hff4b; 
        10'b0111011000: data <= 16'hff88; 
        10'b0111011001: data <= 16'h0004; 
        10'b0111011010: data <= 16'hffe6; 
        10'b0111011011: data <= 16'h0017; 
        10'b0111011100: data <= 16'h000e; 
        10'b0111011101: data <= 16'hfff7; 
        10'b0111011110: data <= 16'hffdf; 
        10'b0111011111: data <= 16'hffd0; 
        10'b0111100000: data <= 16'hffa6; 
        10'b0111100001: data <= 16'hff92; 
        10'b0111100010: data <= 16'hffa6; 
        10'b0111100011: data <= 16'h0029; 
        10'b0111100100: data <= 16'h004f; 
        10'b0111100101: data <= 16'h005a; 
        10'b0111100110: data <= 16'h008a; 
        10'b0111100111: data <= 16'h00c8; 
        10'b0111101000: data <= 16'h007a; 
        10'b0111101001: data <= 16'h0039; 
        10'b0111101010: data <= 16'h004e; 
        10'b0111101011: data <= 16'h00c7; 
        10'b0111101100: data <= 16'h003b; 
        10'b0111101101: data <= 16'hffd8; 
        10'b0111101110: data <= 16'hffa8; 
        10'b0111101111: data <= 16'hff36; 
        10'b0111110000: data <= 16'hff38; 
        10'b0111110001: data <= 16'hff29; 
        10'b0111110010: data <= 16'hff36; 
        10'b0111110011: data <= 16'hff6b; 
        10'b0111110100: data <= 16'hff94; 
        10'b0111110101: data <= 16'h000b; 
        10'b0111110110: data <= 16'h000b; 
        10'b0111110111: data <= 16'hfff6; 
        10'b0111111000: data <= 16'h0027; 
        10'b0111111001: data <= 16'h0000; 
        10'b0111111010: data <= 16'hffe9; 
        10'b0111111011: data <= 16'hfff7; 
        10'b0111111100: data <= 16'hffb1; 
        10'b0111111101: data <= 16'hff4a; 
        10'b0111111110: data <= 16'hff47; 
        10'b0111111111: data <= 16'hff4a; 
        10'b1000000000: data <= 16'hffb4; 
        10'b1000000001: data <= 16'h001e; 
        10'b1000000010: data <= 16'h00dc; 
        10'b1000000011: data <= 16'h00b1; 
        10'b1000000100: data <= 16'hff94; 
        10'b1000000101: data <= 16'hff92; 
        10'b1000000110: data <= 16'h0007; 
        10'b1000000111: data <= 16'h0084; 
        10'b1000001000: data <= 16'hffaf; 
        10'b1000001001: data <= 16'hffa4; 
        10'b1000001010: data <= 16'hff53; 
        10'b1000001011: data <= 16'hff98; 
        10'b1000001100: data <= 16'hff9f; 
        10'b1000001101: data <= 16'hff68; 
        10'b1000001110: data <= 16'hff60; 
        10'b1000001111: data <= 16'hff58; 
        10'b1000010000: data <= 16'hff89; 
        10'b1000010001: data <= 16'hffed; 
        10'b1000010010: data <= 16'h0002; 
        10'b1000010011: data <= 16'h0023; 
        10'b1000010100: data <= 16'h0019; 
        10'b1000010101: data <= 16'h0032; 
        10'b1000010110: data <= 16'h0009; 
        10'b1000010111: data <= 16'hffd5; 
        10'b1000011000: data <= 16'hffb7; 
        10'b1000011001: data <= 16'hff7f; 
        10'b1000011010: data <= 16'hff35; 
        10'b1000011011: data <= 16'hff2f; 
        10'b1000011100: data <= 16'hff28; 
        10'b1000011101: data <= 16'hff2a; 
        10'b1000011110: data <= 16'hff10; 
        10'b1000011111: data <= 16'hff35; 
        10'b1000100000: data <= 16'hfefa; 
        10'b1000100001: data <= 16'hff49; 
        10'b1000100010: data <= 16'hff65; 
        10'b1000100011: data <= 16'hff50; 
        10'b1000100100: data <= 16'hff68; 
        10'b1000100101: data <= 16'hffce; 
        10'b1000100110: data <= 16'hff8d; 
        10'b1000100111: data <= 16'hffe0; 
        10'b1000101000: data <= 16'hffb3; 
        10'b1000101001: data <= 16'hffa5; 
        10'b1000101010: data <= 16'hffaa; 
        10'b1000101011: data <= 16'hffb3; 
        10'b1000101100: data <= 16'hffd0; 
        10'b1000101101: data <= 16'h000e; 
        10'b1000101110: data <= 16'hfff1; 
        10'b1000101111: data <= 16'h0005; 
        10'b1000110000: data <= 16'hfff7; 
        10'b1000110001: data <= 16'h0007; 
        10'b1000110010: data <= 16'h0015; 
        10'b1000110011: data <= 16'h0002; 
        10'b1000110100: data <= 16'hffb5; 
        10'b1000110101: data <= 16'hff84; 
        10'b1000110110: data <= 16'hff44; 
        10'b1000110111: data <= 16'hfed9; 
        10'b1000111000: data <= 16'hfeae; 
        10'b1000111001: data <= 16'hfe85; 
        10'b1000111010: data <= 16'hfdff; 
        10'b1000111011: data <= 16'hfe77; 
        10'b1000111100: data <= 16'hfe81; 
        10'b1000111101: data <= 16'hff83; 
        10'b1000111110: data <= 16'hff50; 
        10'b1000111111: data <= 16'hffae; 
        10'b1001000000: data <= 16'hff9d; 
        10'b1001000001: data <= 16'hffe5; 
        10'b1001000010: data <= 16'hff58; 
        10'b1001000011: data <= 16'hffc9; 
        10'b1001000100: data <= 16'hffbd; 
        10'b1001000101: data <= 16'hff95; 
        10'b1001000110: data <= 16'hffe2; 
        10'b1001000111: data <= 16'hffcd; 
        10'b1001001000: data <= 16'h0005; 
        10'b1001001001: data <= 16'h002b; 
        10'b1001001010: data <= 16'h001a; 
        10'b1001001011: data <= 16'h0008; 
        10'b1001001100: data <= 16'h0003; 
        10'b1001001101: data <= 16'h0000; 
        10'b1001001110: data <= 16'h002b; 
        10'b1001001111: data <= 16'hffd3; 
        10'b1001010000: data <= 16'hffcd; 
        10'b1001010001: data <= 16'hff86; 
        10'b1001010010: data <= 16'hff53; 
        10'b1001010011: data <= 16'hfef5; 
        10'b1001010100: data <= 16'hfed1; 
        10'b1001010101: data <= 16'hfeb3; 
        10'b1001010110: data <= 16'hfea2; 
        10'b1001010111: data <= 16'hfec6; 
        10'b1001011000: data <= 16'hff38; 
        10'b1001011001: data <= 16'hff3a; 
        10'b1001011010: data <= 16'hff37; 
        10'b1001011011: data <= 16'hff8d; 
        10'b1001011100: data <= 16'hff83; 
        10'b1001011101: data <= 16'hff44; 
        10'b1001011110: data <= 16'hff1d; 
        10'b1001011111: data <= 16'hffa0; 
        10'b1001100000: data <= 16'hffca; 
        10'b1001100001: data <= 16'hffe1; 
        10'b1001100010: data <= 16'h000f; 
        10'b1001100011: data <= 16'hfffc; 
        10'b1001100100: data <= 16'h0013; 
        10'b1001100101: data <= 16'h001a; 
        10'b1001100110: data <= 16'h0001; 
        10'b1001100111: data <= 16'h0003; 
        10'b1001101000: data <= 16'h0021; 
        10'b1001101001: data <= 16'h0008; 
        10'b1001101010: data <= 16'h0009; 
        10'b1001101011: data <= 16'h001f; 
        10'b1001101100: data <= 16'hffec; 
        10'b1001101101: data <= 16'hff9d; 
        10'b1001101110: data <= 16'hff62; 
        10'b1001101111: data <= 16'hff29; 
        10'b1001110000: data <= 16'hff60; 
        10'b1001110001: data <= 16'hff59; 
        10'b1001110010: data <= 16'hff49; 
        10'b1001110011: data <= 16'hff85; 
        10'b1001110100: data <= 16'hff75; 
        10'b1001110101: data <= 16'hff47; 
        10'b1001110110: data <= 16'hff65; 
        10'b1001110111: data <= 16'hff26; 
        10'b1001111000: data <= 16'hff0f; 
        10'b1001111001: data <= 16'hff14; 
        10'b1001111010: data <= 16'hff3c; 
        10'b1001111011: data <= 16'hff52; 
        10'b1001111100: data <= 16'hffd0; 
        10'b1001111101: data <= 16'h003b; 
        10'b1001111110: data <= 16'h0021; 
        10'b1001111111: data <= 16'h0028; 
        10'b1010000000: data <= 16'h0042; 
        10'b1010000001: data <= 16'h000e; 
        10'b1010000010: data <= 16'h000f; 
        10'b1010000011: data <= 16'h0018; 
        10'b1010000100: data <= 16'h0027; 
        10'b1010000101: data <= 16'h001e; 
        10'b1010000110: data <= 16'h000b; 
        10'b1010000111: data <= 16'hfff1; 
        10'b1010001000: data <= 16'hffe4; 
        10'b1010001001: data <= 16'hffab; 
        10'b1010001010: data <= 16'hff9d; 
        10'b1010001011: data <= 16'hff7d; 
        10'b1010001100: data <= 16'hfff6; 
        10'b1010001101: data <= 16'hffcb; 
        10'b1010001110: data <= 16'hffd6; 
        10'b1010001111: data <= 16'hff61; 
        10'b1010010000: data <= 16'hff7f; 
        10'b1010010001: data <= 16'hff5d; 
        10'b1010010010: data <= 16'hff76; 
        10'b1010010011: data <= 16'hff15; 
        10'b1010010100: data <= 16'hff02; 
        10'b1010010101: data <= 16'hff20; 
        10'b1010010110: data <= 16'hff75; 
        10'b1010010111: data <= 16'hfff2; 
        10'b1010011000: data <= 16'h0037; 
        10'b1010011001: data <= 16'h007f; 
        10'b1010011010: data <= 16'h00b6; 
        10'b1010011011: data <= 16'h0099; 
        10'b1010011100: data <= 16'h0047; 
        10'b1010011101: data <= 16'hfffb; 
        10'b1010011110: data <= 16'h0033; 
        10'b1010011111: data <= 16'hfffa; 
        10'b1010100000: data <= 16'h0000; 
        10'b1010100001: data <= 16'hffec; 
        10'b1010100010: data <= 16'hfffb; 
        10'b1010100011: data <= 16'h002b; 
        10'b1010100100: data <= 16'h001f; 
        10'b1010100101: data <= 16'h0031; 
        10'b1010100110: data <= 16'h0023; 
        10'b1010100111: data <= 16'h0033; 
        10'b1010101000: data <= 16'h0049; 
        10'b1010101001: data <= 16'h0027; 
        10'b1010101010: data <= 16'hffe6; 
        10'b1010101011: data <= 16'hffaf; 
        10'b1010101100: data <= 16'hfffa; 
        10'b1010101101: data <= 16'hff83; 
        10'b1010101110: data <= 16'hff62; 
        10'b1010101111: data <= 16'hff59; 
        10'b1010110000: data <= 16'hffb4; 
        10'b1010110001: data <= 16'h0037; 
        10'b1010110010: data <= 16'h005e; 
        10'b1010110011: data <= 16'h0061; 
        10'b1010110100: data <= 16'h00dd; 
        10'b1010110101: data <= 16'h00ed; 
        10'b1010110110: data <= 16'h0089; 
        10'b1010110111: data <= 16'h0054; 
        10'b1010111000: data <= 16'h0042; 
        10'b1010111001: data <= 16'hfff3; 
        10'b1010111010: data <= 16'h001d; 
        10'b1010111011: data <= 16'hfffe; 
        10'b1010111100: data <= 16'h000b; 
        10'b1010111101: data <= 16'h002b; 
        10'b1010111110: data <= 16'h002b; 
        10'b1010111111: data <= 16'hfffb; 
        10'b1011000000: data <= 16'h0004; 
        10'b1011000001: data <= 16'h0049; 
        10'b1011000010: data <= 16'h0038; 
        10'b1011000011: data <= 16'h00a0; 
        10'b1011000100: data <= 16'h00b0; 
        10'b1011000101: data <= 16'h00b3; 
        10'b1011000110: data <= 16'h009b; 
        10'b1011000111: data <= 16'h003d; 
        10'b1011001000: data <= 16'h00a3; 
        10'b1011001001: data <= 16'h0091; 
        10'b1011001010: data <= 16'h008b; 
        10'b1011001011: data <= 16'h0083; 
        10'b1011001100: data <= 16'h00f4; 
        10'b1011001101: data <= 16'h0109; 
        10'b1011001110: data <= 16'h0124; 
        10'b1011001111: data <= 16'h0131; 
        10'b1011010000: data <= 16'h0154; 
        10'b1011010001: data <= 16'h00f1; 
        10'b1011010010: data <= 16'h005e; 
        10'b1011010011: data <= 16'h002d; 
        10'b1011010100: data <= 16'hfffa; 
        10'b1011010101: data <= 16'hfffc; 
        10'b1011010110: data <= 16'h000c; 
        10'b1011010111: data <= 16'h000a; 
        10'b1011011000: data <= 16'h0002; 
        10'b1011011001: data <= 16'h0027; 
        10'b1011011010: data <= 16'h000a; 
        10'b1011011011: data <= 16'hfff2; 
        10'b1011011100: data <= 16'h0027; 
        10'b1011011101: data <= 16'h003d; 
        10'b1011011110: data <= 16'h0055; 
        10'b1011011111: data <= 16'h0076; 
        10'b1011100000: data <= 16'h0087; 
        10'b1011100001: data <= 16'h00cd; 
        10'b1011100010: data <= 16'h00d3; 
        10'b1011100011: data <= 16'h00ed; 
        10'b1011100100: data <= 16'h0119; 
        10'b1011100101: data <= 16'h011b; 
        10'b1011100110: data <= 16'h015b; 
        10'b1011100111: data <= 16'h00c8; 
        10'b1011101000: data <= 16'h0089; 
        10'b1011101001: data <= 16'h0074; 
        10'b1011101010: data <= 16'h00ab; 
        10'b1011101011: data <= 16'h00b8; 
        10'b1011101100: data <= 16'h0086; 
        10'b1011101101: data <= 16'h005d; 
        10'b1011101110: data <= 16'h0027; 
        10'b1011101111: data <= 16'h000e; 
        10'b1011110000: data <= 16'h0009; 
        10'b1011110001: data <= 16'h000f; 
        10'b1011110010: data <= 16'hfff1; 
        10'b1011110011: data <= 16'h0009; 
        10'b1011110100: data <= 16'hfff7; 
        10'b1011110101: data <= 16'h0012; 
        10'b1011110110: data <= 16'hfff0; 
        10'b1011110111: data <= 16'h002f; 
        10'b1011111000: data <= 16'h001b; 
        10'b1011111001: data <= 16'h000f; 
        10'b1011111010: data <= 16'hfff9; 
        10'b1011111011: data <= 16'h002e; 
        10'b1011111100: data <= 16'h0027; 
        10'b1011111101: data <= 16'h001b; 
        10'b1011111110: data <= 16'hfff7; 
        10'b1011111111: data <= 16'hfff6; 
        10'b1100000000: data <= 16'h0009; 
        10'b1100000001: data <= 16'hfff7; 
        10'b1100000010: data <= 16'h000a; 
        10'b1100000011: data <= 16'h001e; 
        10'b1100000100: data <= 16'h0003; 
        10'b1100000101: data <= 16'h0010; 
        10'b1100000110: data <= 16'h0034; 
        10'b1100000111: data <= 16'h002f; 
        10'b1100001000: data <= 16'h001a; 
        10'b1100001001: data <= 16'h0010; 
        10'b1100001010: data <= 16'hfff3; 
        10'b1100001011: data <= 16'h0034; 
        10'b1100001100: data <= 16'h001c; 
        10'b1100001101: data <= 16'hfff6; 
        10'b1100001110: data <= 16'h0004; 
        10'b1100001111: data <= 16'hfffb; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 11) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 17'h00048; 
        10'b0000000001: data <= 17'h0003f; 
        10'b0000000010: data <= 17'h1ffec; 
        10'b0000000011: data <= 17'h0002c; 
        10'b0000000100: data <= 17'h00029; 
        10'b0000000101: data <= 17'h00042; 
        10'b0000000110: data <= 17'h1ffe7; 
        10'b0000000111: data <= 17'h0000c; 
        10'b0000001000: data <= 17'h0004c; 
        10'b0000001001: data <= 17'h1ffe1; 
        10'b0000001010: data <= 17'h1fff7; 
        10'b0000001011: data <= 17'h00021; 
        10'b0000001100: data <= 17'h00060; 
        10'b0000001101: data <= 17'h0003f; 
        10'b0000001110: data <= 17'h1ffd9; 
        10'b0000001111: data <= 17'h1ffee; 
        10'b0000010000: data <= 17'h1ffec; 
        10'b0000010001: data <= 17'h00026; 
        10'b0000010010: data <= 17'h00046; 
        10'b0000010011: data <= 17'h00005; 
        10'b0000010100: data <= 17'h00007; 
        10'b0000010101: data <= 17'h1fffb; 
        10'b0000010110: data <= 17'h1ffe1; 
        10'b0000010111: data <= 17'h0000b; 
        10'b0000011000: data <= 17'h0004e; 
        10'b0000011001: data <= 17'h00018; 
        10'b0000011010: data <= 17'h1ffdc; 
        10'b0000011011: data <= 17'h00027; 
        10'b0000011100: data <= 17'h00041; 
        10'b0000011101: data <= 17'h00036; 
        10'b0000011110: data <= 17'h0001a; 
        10'b0000011111: data <= 17'h1fff1; 
        10'b0000100000: data <= 17'h1ffda; 
        10'b0000100001: data <= 17'h1ffe1; 
        10'b0000100010: data <= 17'h1fffa; 
        10'b0000100011: data <= 17'h00061; 
        10'b0000100100: data <= 17'h1ffdb; 
        10'b0000100101: data <= 17'h0004f; 
        10'b0000100110: data <= 17'h0001e; 
        10'b0000100111: data <= 17'h00031; 
        10'b0000101000: data <= 17'h00026; 
        10'b0000101001: data <= 17'h00037; 
        10'b0000101010: data <= 17'h00001; 
        10'b0000101011: data <= 17'h1ffd5; 
        10'b0000101100: data <= 17'h1ffea; 
        10'b0000101101: data <= 17'h0003c; 
        10'b0000101110: data <= 17'h1fffd; 
        10'b0000101111: data <= 17'h00011; 
        10'b0000110000: data <= 17'h0004c; 
        10'b0000110001: data <= 17'h1fffa; 
        10'b0000110010: data <= 17'h0000d; 
        10'b0000110011: data <= 17'h00007; 
        10'b0000110100: data <= 17'h0002a; 
        10'b0000110101: data <= 17'h00051; 
        10'b0000110110: data <= 17'h1ffff; 
        10'b0000110111: data <= 17'h00011; 
        10'b0000111000: data <= 17'h00056; 
        10'b0000111001: data <= 17'h00058; 
        10'b0000111010: data <= 17'h00007; 
        10'b0000111011: data <= 17'h0003c; 
        10'b0000111100: data <= 17'h00049; 
        10'b0000111101: data <= 17'h1fffd; 
        10'b0000111110: data <= 17'h1fff7; 
        10'b0000111111: data <= 17'h0001a; 
        10'b0001000000: data <= 17'h00049; 
        10'b0001000001: data <= 17'h1fff6; 
        10'b0001000010: data <= 17'h1ffea; 
        10'b0001000011: data <= 17'h00038; 
        10'b0001000100: data <= 17'h00021; 
        10'b0001000101: data <= 17'h00046; 
        10'b0001000110: data <= 17'h1ffd7; 
        10'b0001000111: data <= 17'h0004a; 
        10'b0001001000: data <= 17'h1ffe6; 
        10'b0001001001: data <= 17'h1ffe4; 
        10'b0001001010: data <= 17'h00007; 
        10'b0001001011: data <= 17'h1ffdd; 
        10'b0001001100: data <= 17'h00054; 
        10'b0001001101: data <= 17'h1ffea; 
        10'b0001001110: data <= 17'h1ffe2; 
        10'b0001001111: data <= 17'h00054; 
        10'b0001010000: data <= 17'h0000f; 
        10'b0001010001: data <= 17'h0000f; 
        10'b0001010010: data <= 17'h00013; 
        10'b0001010011: data <= 17'h00025; 
        10'b0001010100: data <= 17'h00069; 
        10'b0001010101: data <= 17'h00004; 
        10'b0001010110: data <= 17'h1fff6; 
        10'b0001010111: data <= 17'h0001f; 
        10'b0001011000: data <= 17'h00021; 
        10'b0001011001: data <= 17'h1ffdd; 
        10'b0001011010: data <= 17'h00056; 
        10'b0001011011: data <= 17'h0002f; 
        10'b0001011100: data <= 17'h1ffef; 
        10'b0001011101: data <= 17'h00056; 
        10'b0001011110: data <= 17'h0001b; 
        10'b0001011111: data <= 17'h00044; 
        10'b0001100000: data <= 17'h1fff9; 
        10'b0001100001: data <= 17'h1ffb2; 
        10'b0001100010: data <= 17'h1fff9; 
        10'b0001100011: data <= 17'h1ff8a; 
        10'b0001100100: data <= 17'h1fff1; 
        10'b0001100101: data <= 17'h1ffc2; 
        10'b0001100110: data <= 17'h00014; 
        10'b0001100111: data <= 17'h0000c; 
        10'b0001101000: data <= 17'h0001a; 
        10'b0001101001: data <= 17'h1fff9; 
        10'b0001101010: data <= 17'h00044; 
        10'b0001101011: data <= 17'h1fff7; 
        10'b0001101100: data <= 17'h1fff6; 
        10'b0001101101: data <= 17'h0005e; 
        10'b0001101110: data <= 17'h00023; 
        10'b0001101111: data <= 17'h0003b; 
        10'b0001110000: data <= 17'h0000b; 
        10'b0001110001: data <= 17'h00013; 
        10'b0001110010: data <= 17'h00005; 
        10'b0001110011: data <= 17'h1ffec; 
        10'b0001110100: data <= 17'h1ffdf; 
        10'b0001110101: data <= 17'h0003c; 
        10'b0001110110: data <= 17'h0002a; 
        10'b0001110111: data <= 17'h1fff8; 
        10'b0001111000: data <= 17'h1ffcb; 
        10'b0001111001: data <= 17'h00014; 
        10'b0001111010: data <= 17'h1ffa8; 
        10'b0001111011: data <= 17'h1ff85; 
        10'b0001111100: data <= 17'h1ff52; 
        10'b0001111101: data <= 17'h1fec5; 
        10'b0001111110: data <= 17'h1fe6f; 
        10'b0001111111: data <= 17'h1fde8; 
        10'b0010000000: data <= 17'h1fe74; 
        10'b0010000001: data <= 17'h1fe73; 
        10'b0010000010: data <= 17'h1fed9; 
        10'b0010000011: data <= 17'h1ff7e; 
        10'b0010000100: data <= 17'h1ffc3; 
        10'b0010000101: data <= 17'h1ffd4; 
        10'b0010000110: data <= 17'h0000f; 
        10'b0010000111: data <= 17'h0004b; 
        10'b0010001000: data <= 17'h0003a; 
        10'b0010001001: data <= 17'h00036; 
        10'b0010001010: data <= 17'h00000; 
        10'b0010001011: data <= 17'h00003; 
        10'b0010001100: data <= 17'h00048; 
        10'b0010001101: data <= 17'h00033; 
        10'b0010001110: data <= 17'h0003c; 
        10'b0010001111: data <= 17'h00026; 
        10'b0010010000: data <= 17'h0002e; 
        10'b0010010001: data <= 17'h1ffc7; 
        10'b0010010010: data <= 17'h1ffcd; 
        10'b0010010011: data <= 17'h1ffc8; 
        10'b0010010100: data <= 17'h1ff4a; 
        10'b0010010101: data <= 17'h1ff4e; 
        10'b0010010110: data <= 17'h1ff3f; 
        10'b0010010111: data <= 17'h1ff03; 
        10'b0010011000: data <= 17'h1fec2; 
        10'b0010011001: data <= 17'h1fe88; 
        10'b0010011010: data <= 17'h1fdc3; 
        10'b0010011011: data <= 17'h1fd95; 
        10'b0010011100: data <= 17'h1fcf1; 
        10'b0010011101: data <= 17'h1fdfc; 
        10'b0010011110: data <= 17'h1febb; 
        10'b0010011111: data <= 17'h1ff62; 
        10'b0010100000: data <= 17'h1ff5a; 
        10'b0010100001: data <= 17'h1ff28; 
        10'b0010100010: data <= 17'h1ff37; 
        10'b0010100011: data <= 17'h1ff70; 
        10'b0010100100: data <= 17'h1ffc7; 
        10'b0010100101: data <= 17'h1ffe5; 
        10'b0010100110: data <= 17'h00009; 
        10'b0010100111: data <= 17'h00033; 
        10'b0010101000: data <= 17'h00041; 
        10'b0010101001: data <= 17'h00043; 
        10'b0010101010: data <= 17'h1ffd6; 
        10'b0010101011: data <= 17'h00043; 
        10'b0010101100: data <= 17'h0002b; 
        10'b0010101101: data <= 17'h1ff3f; 
        10'b0010101110: data <= 17'h1ff15; 
        10'b0010101111: data <= 17'h1feeb; 
        10'b0010110000: data <= 17'h1fec7; 
        10'b0010110001: data <= 17'h1fe80; 
        10'b0010110010: data <= 17'h1fee6; 
        10'b0010110011: data <= 17'h1ffa6; 
        10'b0010110100: data <= 17'h00017; 
        10'b0010110101: data <= 17'h0015a; 
        10'b0010110110: data <= 17'h00205; 
        10'b0010110111: data <= 17'h0019b; 
        10'b0010111000: data <= 17'h00120; 
        10'b0010111001: data <= 17'h000ef; 
        10'b0010111010: data <= 17'h0012f; 
        10'b0010111011: data <= 17'h1ffcd; 
        10'b0010111100: data <= 17'h1ffb7; 
        10'b0010111101: data <= 17'h1ff19; 
        10'b0010111110: data <= 17'h1fe62; 
        10'b0010111111: data <= 17'h1fe7f; 
        10'b0011000000: data <= 17'h1ff23; 
        10'b0011000001: data <= 17'h1ff95; 
        10'b0011000010: data <= 17'h1fff0; 
        10'b0011000011: data <= 17'h00023; 
        10'b0011000100: data <= 17'h00064; 
        10'b0011000101: data <= 17'h1fffc; 
        10'b0011000110: data <= 17'h1ffe0; 
        10'b0011000111: data <= 17'h1ffdc; 
        10'b0011001000: data <= 17'h1ff23; 
        10'b0011001001: data <= 17'h1feb0; 
        10'b0011001010: data <= 17'h1fe74; 
        10'b0011001011: data <= 17'h1fe29; 
        10'b0011001100: data <= 17'h1fe42; 
        10'b0011001101: data <= 17'h1ff63; 
        10'b0011001110: data <= 17'h1fff3; 
        10'b0011001111: data <= 17'h0007a; 
        10'b0011010000: data <= 17'h001d5; 
        10'b0011010001: data <= 17'h00230; 
        10'b0011010010: data <= 17'h00300; 
        10'b0011010011: data <= 17'h00304; 
        10'b0011010100: data <= 17'h00323; 
        10'b0011010101: data <= 17'h0016c; 
        10'b0011010110: data <= 17'h00112; 
        10'b0011010111: data <= 17'h0001e; 
        10'b0011011000: data <= 17'h00047; 
        10'b0011011001: data <= 17'h00051; 
        10'b0011011010: data <= 17'h1feeb; 
        10'b0011011011: data <= 17'h1fe10; 
        10'b0011011100: data <= 17'h1fedc; 
        10'b0011011101: data <= 17'h1ffb7; 
        10'b0011011110: data <= 17'h1ffb5; 
        10'b0011011111: data <= 17'h00042; 
        10'b0011100000: data <= 17'h00061; 
        10'b0011100001: data <= 17'h00061; 
        10'b0011100010: data <= 17'h00031; 
        10'b0011100011: data <= 17'h1ffe2; 
        10'b0011100100: data <= 17'h1ff1a; 
        10'b0011100101: data <= 17'h1fea4; 
        10'b0011100110: data <= 17'h1fe6a; 
        10'b0011100111: data <= 17'h1fdc9; 
        10'b0011101000: data <= 17'h1ff6a; 
        10'b0011101001: data <= 17'h1ffbb; 
        10'b0011101010: data <= 17'h1ffb0; 
        10'b0011101011: data <= 17'h1ff5f; 
        10'b0011101100: data <= 17'h1fff4; 
        10'b0011101101: data <= 17'h000e1; 
        10'b0011101110: data <= 17'h00292; 
        10'b0011101111: data <= 17'h0016b; 
        10'b0011110000: data <= 17'h00172; 
        10'b0011110001: data <= 17'h0004c; 
        10'b0011110010: data <= 17'h0001d; 
        10'b0011110011: data <= 17'h00014; 
        10'b0011110100: data <= 17'h1ff86; 
        10'b0011110101: data <= 17'h0003f; 
        10'b0011110110: data <= 17'h1ff64; 
        10'b0011110111: data <= 17'h1fe75; 
        10'b0011111000: data <= 17'h1feb2; 
        10'b0011111001: data <= 17'h1ff60; 
        10'b0011111010: data <= 17'h1ffba; 
        10'b0011111011: data <= 17'h0005a; 
        10'b0011111100: data <= 17'h0001d; 
        10'b0011111101: data <= 17'h00012; 
        10'b0011111110: data <= 17'h00007; 
        10'b0011111111: data <= 17'h1ff5b; 
        10'b0100000000: data <= 17'h1fe99; 
        10'b0100000001: data <= 17'h1feed; 
        10'b0100000010: data <= 17'h1ffb2; 
        10'b0100000011: data <= 17'h1ff62; 
        10'b0100000100: data <= 17'h1ffa2; 
        10'b0100000101: data <= 17'h1ffd5; 
        10'b0100000110: data <= 17'h000a9; 
        10'b0100000111: data <= 17'h00066; 
        10'b0100001000: data <= 17'h0001e; 
        10'b0100001001: data <= 17'h00110; 
        10'b0100001010: data <= 17'h001c7; 
        10'b0100001011: data <= 17'h00196; 
        10'b0100001100: data <= 17'h1fff0; 
        10'b0100001101: data <= 17'h1ff8c; 
        10'b0100001110: data <= 17'h00004; 
        10'b0100001111: data <= 17'h1ff0e; 
        10'b0100010000: data <= 17'h1ff99; 
        10'b0100010001: data <= 17'h1ff02; 
        10'b0100010010: data <= 17'h1fef0; 
        10'b0100010011: data <= 17'h1fede; 
        10'b0100010100: data <= 17'h1ff3a; 
        10'b0100010101: data <= 17'h1ffaa; 
        10'b0100010110: data <= 17'h1ffc1; 
        10'b0100010111: data <= 17'h00050; 
        10'b0100011000: data <= 17'h00011; 
        10'b0100011001: data <= 17'h1fffd; 
        10'b0100011010: data <= 17'h1ffd9; 
        10'b0100011011: data <= 17'h1ffc1; 
        10'b0100011100: data <= 17'h1feeb; 
        10'b0100011101: data <= 17'h1ff6f; 
        10'b0100011110: data <= 17'h00087; 
        10'b0100011111: data <= 17'h000b1; 
        10'b0100100000: data <= 17'h00166; 
        10'b0100100001: data <= 17'h00164; 
        10'b0100100010: data <= 17'h00132; 
        10'b0100100011: data <= 17'h001cd; 
        10'b0100100100: data <= 17'h000e8; 
        10'b0100100101: data <= 17'h00037; 
        10'b0100100110: data <= 17'h0003b; 
        10'b0100100111: data <= 17'h1ff16; 
        10'b0100101000: data <= 17'h1ff75; 
        10'b0100101001: data <= 17'h1ffe4; 
        10'b0100101010: data <= 17'h000a3; 
        10'b0100101011: data <= 17'h1fffd; 
        10'b0100101100: data <= 17'h00083; 
        10'b0100101101: data <= 17'h1ffb2; 
        10'b0100101110: data <= 17'h1ff5f; 
        10'b0100101111: data <= 17'h1ff68; 
        10'b0100110000: data <= 17'h1ff40; 
        10'b0100110001: data <= 17'h1ffc9; 
        10'b0100110010: data <= 17'h1ffb7; 
        10'b0100110011: data <= 17'h0002e; 
        10'b0100110100: data <= 17'h1fff1; 
        10'b0100110101: data <= 17'h00012; 
        10'b0100110110: data <= 17'h1ffd6; 
        10'b0100110111: data <= 17'h1ffe6; 
        10'b0100111000: data <= 17'h1ffb4; 
        10'b0100111001: data <= 17'h000fe; 
        10'b0100111010: data <= 17'h0024d; 
        10'b0100111011: data <= 17'h001b7; 
        10'b0100111100: data <= 17'h002b2; 
        10'b0100111101: data <= 17'h00115; 
        10'b0100111110: data <= 17'h0011f; 
        10'b0100111111: data <= 17'h001ed; 
        10'b0101000000: data <= 17'h1ff63; 
        10'b0101000001: data <= 17'h1ff7b; 
        10'b0101000010: data <= 17'h1ffb8; 
        10'b0101000011: data <= 17'h00023; 
        10'b0101000100: data <= 17'h000be; 
        10'b0101000101: data <= 17'h0029b; 
        10'b0101000110: data <= 17'h0013b; 
        10'b0101000111: data <= 17'h0013f; 
        10'b0101001000: data <= 17'h0020c; 
        10'b0101001001: data <= 17'h0017b; 
        10'b0101001010: data <= 17'h000dd; 
        10'b0101001011: data <= 17'h0002e; 
        10'b0101001100: data <= 17'h1ffdc; 
        10'b0101001101: data <= 17'h1ffa6; 
        10'b0101001110: data <= 17'h1fffc; 
        10'b0101001111: data <= 17'h00000; 
        10'b0101010000: data <= 17'h0002a; 
        10'b0101010001: data <= 17'h00056; 
        10'b0101010010: data <= 17'h1ffc5; 
        10'b0101010011: data <= 17'h1ffa1; 
        10'b0101010100: data <= 17'h000d7; 
        10'b0101010101: data <= 17'h0022e; 
        10'b0101010110: data <= 17'h00286; 
        10'b0101010111: data <= 17'h0017f; 
        10'b0101011000: data <= 17'h001df; 
        10'b0101011001: data <= 17'h00249; 
        10'b0101011010: data <= 17'h00176; 
        10'b0101011011: data <= 17'h00004; 
        10'b0101011100: data <= 17'h1fe89; 
        10'b0101011101: data <= 17'h00145; 
        10'b0101011110: data <= 17'h002be; 
        10'b0101011111: data <= 17'h0022b; 
        10'b0101100000: data <= 17'h001db; 
        10'b0101100001: data <= 17'h002d6; 
        10'b0101100010: data <= 17'h002db; 
        10'b0101100011: data <= 17'h002f7; 
        10'b0101100100: data <= 17'h0030c; 
        10'b0101100101: data <= 17'h00209; 
        10'b0101100110: data <= 17'h000fb; 
        10'b0101100111: data <= 17'h00007; 
        10'b0101101000: data <= 17'h1ff8c; 
        10'b0101101001: data <= 17'h00013; 
        10'b0101101010: data <= 17'h0002a; 
        10'b0101101011: data <= 17'h0002e; 
        10'b0101101100: data <= 17'h00060; 
        10'b0101101101: data <= 17'h0003b; 
        10'b0101101110: data <= 17'h1ffaf; 
        10'b0101101111: data <= 17'h0001e; 
        10'b0101110000: data <= 17'h00145; 
        10'b0101110001: data <= 17'h001e8; 
        10'b0101110010: data <= 17'h001cc; 
        10'b0101110011: data <= 17'h0012e; 
        10'b0101110100: data <= 17'h0017b; 
        10'b0101110101: data <= 17'h000f3; 
        10'b0101110110: data <= 17'h000dc; 
        10'b0101110111: data <= 17'h1ff8e; 
        10'b0101111000: data <= 17'h1ff3b; 
        10'b0101111001: data <= 17'h001ff; 
        10'b0101111010: data <= 17'h002bc; 
        10'b0101111011: data <= 17'h001fc; 
        10'b0101111100: data <= 17'h00249; 
        10'b0101111101: data <= 17'h0020c; 
        10'b0101111110: data <= 17'h002cf; 
        10'b0101111111: data <= 17'h002dc; 
        10'b0110000000: data <= 17'h0023c; 
        10'b0110000001: data <= 17'h0014e; 
        10'b0110000010: data <= 17'h00013; 
        10'b0110000011: data <= 17'h1ff1c; 
        10'b0110000100: data <= 17'h1ff7b; 
        10'b0110000101: data <= 17'h1ffd7; 
        10'b0110000110: data <= 17'h0002b; 
        10'b0110000111: data <= 17'h0002c; 
        10'b0110001000: data <= 17'h00013; 
        10'b0110001001: data <= 17'h0000a; 
        10'b0110001010: data <= 17'h00042; 
        10'b0110001011: data <= 17'h0002a; 
        10'b0110001100: data <= 17'h00095; 
        10'b0110001101: data <= 17'h0008c; 
        10'b0110001110: data <= 17'h0017d; 
        10'b0110001111: data <= 17'h0010b; 
        10'b0110010000: data <= 17'h00082; 
        10'b0110010001: data <= 17'h1ffff; 
        10'b0110010010: data <= 17'h0002f; 
        10'b0110010011: data <= 17'h1ffe8; 
        10'b0110010100: data <= 17'h1ff70; 
        10'b0110010101: data <= 17'h000a6; 
        10'b0110010110: data <= 17'h0005e; 
        10'b0110010111: data <= 17'h001c0; 
        10'b0110011000: data <= 17'h001db; 
        10'b0110011001: data <= 17'h001dc; 
        10'b0110011010: data <= 17'h00144; 
        10'b0110011011: data <= 17'h000d0; 
        10'b0110011100: data <= 17'h00104; 
        10'b0110011101: data <= 17'h00005; 
        10'b0110011110: data <= 17'h1fefa; 
        10'b0110011111: data <= 17'h1fe83; 
        10'b0110100000: data <= 17'h1ff62; 
        10'b0110100001: data <= 17'h0001a; 
        10'b0110100010: data <= 17'h0000f; 
        10'b0110100011: data <= 17'h00012; 
        10'b0110100100: data <= 17'h00049; 
        10'b0110100101: data <= 17'h00043; 
        10'b0110100110: data <= 17'h0002c; 
        10'b0110100111: data <= 17'h1ffcb; 
        10'b0110101000: data <= 17'h0000b; 
        10'b0110101001: data <= 17'h000aa; 
        10'b0110101010: data <= 17'h000a2; 
        10'b0110101011: data <= 17'h0006b; 
        10'b0110101100: data <= 17'h0006d; 
        10'b0110101101: data <= 17'h1ff37; 
        10'b0110101110: data <= 17'h1ffa3; 
        10'b0110101111: data <= 17'h1ffa2; 
        10'b0110110000: data <= 17'h1ff74; 
        10'b0110110001: data <= 17'h1ff93; 
        10'b0110110010: data <= 17'h1ff7c; 
        10'b0110110011: data <= 17'h001e9; 
        10'b0110110100: data <= 17'h002cc; 
        10'b0110110101: data <= 17'h002af; 
        10'b0110110110: data <= 17'h00158; 
        10'b0110110111: data <= 17'h00021; 
        10'b0110111000: data <= 17'h1ff6b; 
        10'b0110111001: data <= 17'h1fe76; 
        10'b0110111010: data <= 17'h1fe15; 
        10'b0110111011: data <= 17'h1fea1; 
        10'b0110111100: data <= 17'h1ff64; 
        10'b0110111101: data <= 17'h00003; 
        10'b0110111110: data <= 17'h00028; 
        10'b0110111111: data <= 17'h1fffa; 
        10'b0111000000: data <= 17'h00054; 
        10'b0111000001: data <= 17'h00007; 
        10'b0111000010: data <= 17'h1ffc4; 
        10'b0111000011: data <= 17'h1fff1; 
        10'b0111000100: data <= 17'h00005; 
        10'b0111000101: data <= 17'h00033; 
        10'b0111000110: data <= 17'h1ff7d; 
        10'b0111000111: data <= 17'h00068; 
        10'b0111001000: data <= 17'h00126; 
        10'b0111001001: data <= 17'h1ffbb; 
        10'b0111001010: data <= 17'h000a7; 
        10'b0111001011: data <= 17'h000ed; 
        10'b0111001100: data <= 17'h1ffe0; 
        10'b0111001101: data <= 17'h1fef3; 
        10'b0111001110: data <= 17'h1ffd3; 
        10'b0111001111: data <= 17'h00110; 
        10'b0111010000: data <= 17'h001e9; 
        10'b0111010001: data <= 17'h001e6; 
        10'b0111010010: data <= 17'h00079; 
        10'b0111010011: data <= 17'h1feec; 
        10'b0111010100: data <= 17'h1fe36; 
        10'b0111010101: data <= 17'h1fd86; 
        10'b0111010110: data <= 17'h1fe43; 
        10'b0111010111: data <= 17'h1fe97; 
        10'b0111011000: data <= 17'h1ff11; 
        10'b0111011001: data <= 17'h00008; 
        10'b0111011010: data <= 17'h1ffcc; 
        10'b0111011011: data <= 17'h0002d; 
        10'b0111011100: data <= 17'h0001c; 
        10'b0111011101: data <= 17'h1ffed; 
        10'b0111011110: data <= 17'h1ffbe; 
        10'b0111011111: data <= 17'h1ffa0; 
        10'b0111100000: data <= 17'h1ff4c; 
        10'b0111100001: data <= 17'h1ff25; 
        10'b0111100010: data <= 17'h1ff4b; 
        10'b0111100011: data <= 17'h00051; 
        10'b0111100100: data <= 17'h0009f; 
        10'b0111100101: data <= 17'h000b5; 
        10'b0111100110: data <= 17'h00113; 
        10'b0111100111: data <= 17'h00191; 
        10'b0111101000: data <= 17'h000f4; 
        10'b0111101001: data <= 17'h00072; 
        10'b0111101010: data <= 17'h0009b; 
        10'b0111101011: data <= 17'h0018f; 
        10'b0111101100: data <= 17'h00076; 
        10'b0111101101: data <= 17'h1ffaf; 
        10'b0111101110: data <= 17'h1ff50; 
        10'b0111101111: data <= 17'h1fe6b; 
        10'b0111110000: data <= 17'h1fe70; 
        10'b0111110001: data <= 17'h1fe52; 
        10'b0111110010: data <= 17'h1fe6b; 
        10'b0111110011: data <= 17'h1fed6; 
        10'b0111110100: data <= 17'h1ff27; 
        10'b0111110101: data <= 17'h00016; 
        10'b0111110110: data <= 17'h00016; 
        10'b0111110111: data <= 17'h1ffed; 
        10'b0111111000: data <= 17'h0004e; 
        10'b0111111001: data <= 17'h00000; 
        10'b0111111010: data <= 17'h1ffd3; 
        10'b0111111011: data <= 17'h1ffee; 
        10'b0111111100: data <= 17'h1ff62; 
        10'b0111111101: data <= 17'h1fe94; 
        10'b0111111110: data <= 17'h1fe8d; 
        10'b0111111111: data <= 17'h1fe94; 
        10'b1000000000: data <= 17'h1ff67; 
        10'b1000000001: data <= 17'h0003d; 
        10'b1000000010: data <= 17'h001b7; 
        10'b1000000011: data <= 17'h00163; 
        10'b1000000100: data <= 17'h1ff27; 
        10'b1000000101: data <= 17'h1ff24; 
        10'b1000000110: data <= 17'h0000e; 
        10'b1000000111: data <= 17'h00108; 
        10'b1000001000: data <= 17'h1ff5e; 
        10'b1000001001: data <= 17'h1ff47; 
        10'b1000001010: data <= 17'h1fea7; 
        10'b1000001011: data <= 17'h1ff30; 
        10'b1000001100: data <= 17'h1ff3d; 
        10'b1000001101: data <= 17'h1fed0; 
        10'b1000001110: data <= 17'h1fec0; 
        10'b1000001111: data <= 17'h1feb1; 
        10'b1000010000: data <= 17'h1ff13; 
        10'b1000010001: data <= 17'h1ffda; 
        10'b1000010010: data <= 17'h00005; 
        10'b1000010011: data <= 17'h00047; 
        10'b1000010100: data <= 17'h00032; 
        10'b1000010101: data <= 17'h00065; 
        10'b1000010110: data <= 17'h00012; 
        10'b1000010111: data <= 17'h1ffa9; 
        10'b1000011000: data <= 17'h1ff6f; 
        10'b1000011001: data <= 17'h1feff; 
        10'b1000011010: data <= 17'h1fe69; 
        10'b1000011011: data <= 17'h1fe5f; 
        10'b1000011100: data <= 17'h1fe50; 
        10'b1000011101: data <= 17'h1fe53; 
        10'b1000011110: data <= 17'h1fe20; 
        10'b1000011111: data <= 17'h1fe6b; 
        10'b1000100000: data <= 17'h1fdf3; 
        10'b1000100001: data <= 17'h1fe91; 
        10'b1000100010: data <= 17'h1fecb; 
        10'b1000100011: data <= 17'h1fea0; 
        10'b1000100100: data <= 17'h1fed1; 
        10'b1000100101: data <= 17'h1ff9d; 
        10'b1000100110: data <= 17'h1ff19; 
        10'b1000100111: data <= 17'h1ffc0; 
        10'b1000101000: data <= 17'h1ff66; 
        10'b1000101001: data <= 17'h1ff49; 
        10'b1000101010: data <= 17'h1ff53; 
        10'b1000101011: data <= 17'h1ff66; 
        10'b1000101100: data <= 17'h1ff9f; 
        10'b1000101101: data <= 17'h0001c; 
        10'b1000101110: data <= 17'h1ffe2; 
        10'b1000101111: data <= 17'h0000b; 
        10'b1000110000: data <= 17'h1ffed; 
        10'b1000110001: data <= 17'h0000e; 
        10'b1000110010: data <= 17'h0002b; 
        10'b1000110011: data <= 17'h00003; 
        10'b1000110100: data <= 17'h1ff6a; 
        10'b1000110101: data <= 17'h1ff08; 
        10'b1000110110: data <= 17'h1fe87; 
        10'b1000110111: data <= 17'h1fdb2; 
        10'b1000111000: data <= 17'h1fd5c; 
        10'b1000111001: data <= 17'h1fd0a; 
        10'b1000111010: data <= 17'h1fbfe; 
        10'b1000111011: data <= 17'h1fcee; 
        10'b1000111100: data <= 17'h1fd03; 
        10'b1000111101: data <= 17'h1ff06; 
        10'b1000111110: data <= 17'h1fea1; 
        10'b1000111111: data <= 17'h1ff5b; 
        10'b1001000000: data <= 17'h1ff3a; 
        10'b1001000001: data <= 17'h1ffcb; 
        10'b1001000010: data <= 17'h1feb0; 
        10'b1001000011: data <= 17'h1ff91; 
        10'b1001000100: data <= 17'h1ff7a; 
        10'b1001000101: data <= 17'h1ff2a; 
        10'b1001000110: data <= 17'h1ffc4; 
        10'b1001000111: data <= 17'h1ff99; 
        10'b1001001000: data <= 17'h0000a; 
        10'b1001001001: data <= 17'h00056; 
        10'b1001001010: data <= 17'h00034; 
        10'b1001001011: data <= 17'h00010; 
        10'b1001001100: data <= 17'h00007; 
        10'b1001001101: data <= 17'h00000; 
        10'b1001001110: data <= 17'h00056; 
        10'b1001001111: data <= 17'h1ffa5; 
        10'b1001010000: data <= 17'h1ff9b; 
        10'b1001010001: data <= 17'h1ff0b; 
        10'b1001010010: data <= 17'h1fea6; 
        10'b1001010011: data <= 17'h1fdea; 
        10'b1001010100: data <= 17'h1fda2; 
        10'b1001010101: data <= 17'h1fd65; 
        10'b1001010110: data <= 17'h1fd45; 
        10'b1001010111: data <= 17'h1fd8b; 
        10'b1001011000: data <= 17'h1fe6f; 
        10'b1001011001: data <= 17'h1fe75; 
        10'b1001011010: data <= 17'h1fe6e; 
        10'b1001011011: data <= 17'h1ff19; 
        10'b1001011100: data <= 17'h1ff06; 
        10'b1001011101: data <= 17'h1fe88; 
        10'b1001011110: data <= 17'h1fe3a; 
        10'b1001011111: data <= 17'h1ff40; 
        10'b1001100000: data <= 17'h1ff95; 
        10'b1001100001: data <= 17'h1ffc2; 
        10'b1001100010: data <= 17'h0001e; 
        10'b1001100011: data <= 17'h1fff7; 
        10'b1001100100: data <= 17'h00026; 
        10'b1001100101: data <= 17'h00035; 
        10'b1001100110: data <= 17'h00003; 
        10'b1001100111: data <= 17'h00006; 
        10'b1001101000: data <= 17'h00042; 
        10'b1001101001: data <= 17'h00010; 
        10'b1001101010: data <= 17'h00013; 
        10'b1001101011: data <= 17'h0003f; 
        10'b1001101100: data <= 17'h1ffd8; 
        10'b1001101101: data <= 17'h1ff3a; 
        10'b1001101110: data <= 17'h1fec3; 
        10'b1001101111: data <= 17'h1fe51; 
        10'b1001110000: data <= 17'h1febf; 
        10'b1001110001: data <= 17'h1feb1; 
        10'b1001110010: data <= 17'h1fe92; 
        10'b1001110011: data <= 17'h1ff09; 
        10'b1001110100: data <= 17'h1feea; 
        10'b1001110101: data <= 17'h1fe8f; 
        10'b1001110110: data <= 17'h1feca; 
        10'b1001110111: data <= 17'h1fe4d; 
        10'b1001111000: data <= 17'h1fe1f; 
        10'b1001111001: data <= 17'h1fe28; 
        10'b1001111010: data <= 17'h1fe78; 
        10'b1001111011: data <= 17'h1fea3; 
        10'b1001111100: data <= 17'h1ffa0; 
        10'b1001111101: data <= 17'h00075; 
        10'b1001111110: data <= 17'h00041; 
        10'b1001111111: data <= 17'h00051; 
        10'b1010000000: data <= 17'h00084; 
        10'b1010000001: data <= 17'h0001c; 
        10'b1010000010: data <= 17'h0001f; 
        10'b1010000011: data <= 17'h00030; 
        10'b1010000100: data <= 17'h0004d; 
        10'b1010000101: data <= 17'h0003c; 
        10'b1010000110: data <= 17'h00017; 
        10'b1010000111: data <= 17'h1ffe2; 
        10'b1010001000: data <= 17'h1ffc8; 
        10'b1010001001: data <= 17'h1ff56; 
        10'b1010001010: data <= 17'h1ff3a; 
        10'b1010001011: data <= 17'h1fefa; 
        10'b1010001100: data <= 17'h1ffec; 
        10'b1010001101: data <= 17'h1ff96; 
        10'b1010001110: data <= 17'h1ffab; 
        10'b1010001111: data <= 17'h1fec3; 
        10'b1010010000: data <= 17'h1fefe; 
        10'b1010010001: data <= 17'h1feba; 
        10'b1010010010: data <= 17'h1feec; 
        10'b1010010011: data <= 17'h1fe2a; 
        10'b1010010100: data <= 17'h1fe04; 
        10'b1010010101: data <= 17'h1fe41; 
        10'b1010010110: data <= 17'h1fee9; 
        10'b1010010111: data <= 17'h1ffe5; 
        10'b1010011000: data <= 17'h0006d; 
        10'b1010011001: data <= 17'h000fd; 
        10'b1010011010: data <= 17'h0016d; 
        10'b1010011011: data <= 17'h00132; 
        10'b1010011100: data <= 17'h0008f; 
        10'b1010011101: data <= 17'h1fff6; 
        10'b1010011110: data <= 17'h00067; 
        10'b1010011111: data <= 17'h1fff4; 
        10'b1010100000: data <= 17'h00000; 
        10'b1010100001: data <= 17'h1ffd8; 
        10'b1010100010: data <= 17'h1fff5; 
        10'b1010100011: data <= 17'h00056; 
        10'b1010100100: data <= 17'h0003e; 
        10'b1010100101: data <= 17'h00061; 
        10'b1010100110: data <= 17'h00047; 
        10'b1010100111: data <= 17'h00067; 
        10'b1010101000: data <= 17'h00091; 
        10'b1010101001: data <= 17'h0004e; 
        10'b1010101010: data <= 17'h1ffcc; 
        10'b1010101011: data <= 17'h1ff5d; 
        10'b1010101100: data <= 17'h1fff4; 
        10'b1010101101: data <= 17'h1ff06; 
        10'b1010101110: data <= 17'h1fec5; 
        10'b1010101111: data <= 17'h1feb3; 
        10'b1010110000: data <= 17'h1ff69; 
        10'b1010110001: data <= 17'h0006e; 
        10'b1010110010: data <= 17'h000bb; 
        10'b1010110011: data <= 17'h000c1; 
        10'b1010110100: data <= 17'h001b9; 
        10'b1010110101: data <= 17'h001db; 
        10'b1010110110: data <= 17'h00111; 
        10'b1010110111: data <= 17'h000a7; 
        10'b1010111000: data <= 17'h00084; 
        10'b1010111001: data <= 17'h1ffe6; 
        10'b1010111010: data <= 17'h0003b; 
        10'b1010111011: data <= 17'h1fffc; 
        10'b1010111100: data <= 17'h00015; 
        10'b1010111101: data <= 17'h00056; 
        10'b1010111110: data <= 17'h00056; 
        10'b1010111111: data <= 17'h1fff7; 
        10'b1011000000: data <= 17'h00008; 
        10'b1011000001: data <= 17'h00093; 
        10'b1011000010: data <= 17'h0006f; 
        10'b1011000011: data <= 17'h00141; 
        10'b1011000100: data <= 17'h0015f; 
        10'b1011000101: data <= 17'h00166; 
        10'b1011000110: data <= 17'h00136; 
        10'b1011000111: data <= 17'h0007b; 
        10'b1011001000: data <= 17'h00146; 
        10'b1011001001: data <= 17'h00122; 
        10'b1011001010: data <= 17'h00116; 
        10'b1011001011: data <= 17'h00105; 
        10'b1011001100: data <= 17'h001e8; 
        10'b1011001101: data <= 17'h00213; 
        10'b1011001110: data <= 17'h00248; 
        10'b1011001111: data <= 17'h00261; 
        10'b1011010000: data <= 17'h002a8; 
        10'b1011010001: data <= 17'h001e2; 
        10'b1011010010: data <= 17'h000bc; 
        10'b1011010011: data <= 17'h00059; 
        10'b1011010100: data <= 17'h1fff4; 
        10'b1011010101: data <= 17'h1fff9; 
        10'b1011010110: data <= 17'h00019; 
        10'b1011010111: data <= 17'h00015; 
        10'b1011011000: data <= 17'h00004; 
        10'b1011011001: data <= 17'h0004e; 
        10'b1011011010: data <= 17'h00015; 
        10'b1011011011: data <= 17'h1ffe4; 
        10'b1011011100: data <= 17'h0004e; 
        10'b1011011101: data <= 17'h0007a; 
        10'b1011011110: data <= 17'h000ab; 
        10'b1011011111: data <= 17'h000ed; 
        10'b1011100000: data <= 17'h0010e; 
        10'b1011100001: data <= 17'h00199; 
        10'b1011100010: data <= 17'h001a6; 
        10'b1011100011: data <= 17'h001da; 
        10'b1011100100: data <= 17'h00231; 
        10'b1011100101: data <= 17'h00236; 
        10'b1011100110: data <= 17'h002b6; 
        10'b1011100111: data <= 17'h00190; 
        10'b1011101000: data <= 17'h00112; 
        10'b1011101001: data <= 17'h000e7; 
        10'b1011101010: data <= 17'h00155; 
        10'b1011101011: data <= 17'h00170; 
        10'b1011101100: data <= 17'h0010b; 
        10'b1011101101: data <= 17'h000ba; 
        10'b1011101110: data <= 17'h0004d; 
        10'b1011101111: data <= 17'h0001c; 
        10'b1011110000: data <= 17'h00011; 
        10'b1011110001: data <= 17'h0001f; 
        10'b1011110010: data <= 17'h1ffe3; 
        10'b1011110011: data <= 17'h00011; 
        10'b1011110100: data <= 17'h1ffed; 
        10'b1011110101: data <= 17'h00024; 
        10'b1011110110: data <= 17'h1ffe0; 
        10'b1011110111: data <= 17'h0005f; 
        10'b1011111000: data <= 17'h00036; 
        10'b1011111001: data <= 17'h0001e; 
        10'b1011111010: data <= 17'h1fff3; 
        10'b1011111011: data <= 17'h0005c; 
        10'b1011111100: data <= 17'h0004e; 
        10'b1011111101: data <= 17'h00035; 
        10'b1011111110: data <= 17'h1ffef; 
        10'b1011111111: data <= 17'h1ffed; 
        10'b1100000000: data <= 17'h00012; 
        10'b1100000001: data <= 17'h1ffef; 
        10'b1100000010: data <= 17'h00014; 
        10'b1100000011: data <= 17'h0003b; 
        10'b1100000100: data <= 17'h00005; 
        10'b1100000101: data <= 17'h00020; 
        10'b1100000110: data <= 17'h00069; 
        10'b1100000111: data <= 17'h0005d; 
        10'b1100001000: data <= 17'h00035; 
        10'b1100001001: data <= 17'h00020; 
        10'b1100001010: data <= 17'h1ffe6; 
        10'b1100001011: data <= 17'h00068; 
        10'b1100001100: data <= 17'h00038; 
        10'b1100001101: data <= 17'h1ffed; 
        10'b1100001110: data <= 17'h00007; 
        10'b1100001111: data <= 17'h1fff6; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 12) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 18'h00091; 
        10'b0000000001: data <= 18'h0007f; 
        10'b0000000010: data <= 18'h3ffd9; 
        10'b0000000011: data <= 18'h00059; 
        10'b0000000100: data <= 18'h00052; 
        10'b0000000101: data <= 18'h00085; 
        10'b0000000110: data <= 18'h3ffce; 
        10'b0000000111: data <= 18'h00019; 
        10'b0000001000: data <= 18'h00099; 
        10'b0000001001: data <= 18'h3ffc2; 
        10'b0000001010: data <= 18'h3ffee; 
        10'b0000001011: data <= 18'h00043; 
        10'b0000001100: data <= 18'h000c1; 
        10'b0000001101: data <= 18'h0007e; 
        10'b0000001110: data <= 18'h3ffb1; 
        10'b0000001111: data <= 18'h3ffdc; 
        10'b0000010000: data <= 18'h3ffd8; 
        10'b0000010001: data <= 18'h0004c; 
        10'b0000010010: data <= 18'h0008b; 
        10'b0000010011: data <= 18'h0000a; 
        10'b0000010100: data <= 18'h0000e; 
        10'b0000010101: data <= 18'h3fff6; 
        10'b0000010110: data <= 18'h3ffc2; 
        10'b0000010111: data <= 18'h00016; 
        10'b0000011000: data <= 18'h0009c; 
        10'b0000011001: data <= 18'h0002f; 
        10'b0000011010: data <= 18'h3ffb9; 
        10'b0000011011: data <= 18'h0004e; 
        10'b0000011100: data <= 18'h00082; 
        10'b0000011101: data <= 18'h0006c; 
        10'b0000011110: data <= 18'h00034; 
        10'b0000011111: data <= 18'h3ffe2; 
        10'b0000100000: data <= 18'h3ffb5; 
        10'b0000100001: data <= 18'h3ffc3; 
        10'b0000100010: data <= 18'h3fff4; 
        10'b0000100011: data <= 18'h000c2; 
        10'b0000100100: data <= 18'h3ffb7; 
        10'b0000100101: data <= 18'h0009d; 
        10'b0000100110: data <= 18'h0003d; 
        10'b0000100111: data <= 18'h00061; 
        10'b0000101000: data <= 18'h0004c; 
        10'b0000101001: data <= 18'h0006e; 
        10'b0000101010: data <= 18'h00003; 
        10'b0000101011: data <= 18'h3ffab; 
        10'b0000101100: data <= 18'h3ffd4; 
        10'b0000101101: data <= 18'h00078; 
        10'b0000101110: data <= 18'h3fffb; 
        10'b0000101111: data <= 18'h00022; 
        10'b0000110000: data <= 18'h00098; 
        10'b0000110001: data <= 18'h3fff5; 
        10'b0000110010: data <= 18'h0001b; 
        10'b0000110011: data <= 18'h0000e; 
        10'b0000110100: data <= 18'h00054; 
        10'b0000110101: data <= 18'h000a3; 
        10'b0000110110: data <= 18'h3fffe; 
        10'b0000110111: data <= 18'h00023; 
        10'b0000111000: data <= 18'h000ab; 
        10'b0000111001: data <= 18'h000b0; 
        10'b0000111010: data <= 18'h0000d; 
        10'b0000111011: data <= 18'h00078; 
        10'b0000111100: data <= 18'h00091; 
        10'b0000111101: data <= 18'h3fff9; 
        10'b0000111110: data <= 18'h3ffef; 
        10'b0000111111: data <= 18'h00034; 
        10'b0001000000: data <= 18'h00092; 
        10'b0001000001: data <= 18'h3ffeb; 
        10'b0001000010: data <= 18'h3ffd4; 
        10'b0001000011: data <= 18'h0006f; 
        10'b0001000100: data <= 18'h00042; 
        10'b0001000101: data <= 18'h0008b; 
        10'b0001000110: data <= 18'h3ffae; 
        10'b0001000111: data <= 18'h00093; 
        10'b0001001000: data <= 18'h3ffcb; 
        10'b0001001001: data <= 18'h3ffc8; 
        10'b0001001010: data <= 18'h0000d; 
        10'b0001001011: data <= 18'h3ffba; 
        10'b0001001100: data <= 18'h000a9; 
        10'b0001001101: data <= 18'h3ffd4; 
        10'b0001001110: data <= 18'h3ffc3; 
        10'b0001001111: data <= 18'h000a8; 
        10'b0001010000: data <= 18'h0001e; 
        10'b0001010001: data <= 18'h0001d; 
        10'b0001010010: data <= 18'h00025; 
        10'b0001010011: data <= 18'h0004b; 
        10'b0001010100: data <= 18'h000d1; 
        10'b0001010101: data <= 18'h00007; 
        10'b0001010110: data <= 18'h3ffed; 
        10'b0001010111: data <= 18'h0003e; 
        10'b0001011000: data <= 18'h00042; 
        10'b0001011001: data <= 18'h3ffbb; 
        10'b0001011010: data <= 18'h000ab; 
        10'b0001011011: data <= 18'h0005e; 
        10'b0001011100: data <= 18'h3ffde; 
        10'b0001011101: data <= 18'h000ad; 
        10'b0001011110: data <= 18'h00036; 
        10'b0001011111: data <= 18'h00088; 
        10'b0001100000: data <= 18'h3fff2; 
        10'b0001100001: data <= 18'h3ff64; 
        10'b0001100010: data <= 18'h3fff2; 
        10'b0001100011: data <= 18'h3ff13; 
        10'b0001100100: data <= 18'h3ffe3; 
        10'b0001100101: data <= 18'h3ff85; 
        10'b0001100110: data <= 18'h00029; 
        10'b0001100111: data <= 18'h00019; 
        10'b0001101000: data <= 18'h00035; 
        10'b0001101001: data <= 18'h3fff3; 
        10'b0001101010: data <= 18'h00088; 
        10'b0001101011: data <= 18'h3ffef; 
        10'b0001101100: data <= 18'h3ffec; 
        10'b0001101101: data <= 18'h000bb; 
        10'b0001101110: data <= 18'h00046; 
        10'b0001101111: data <= 18'h00077; 
        10'b0001110000: data <= 18'h00017; 
        10'b0001110001: data <= 18'h00027; 
        10'b0001110010: data <= 18'h00009; 
        10'b0001110011: data <= 18'h3ffd8; 
        10'b0001110100: data <= 18'h3ffbd; 
        10'b0001110101: data <= 18'h00079; 
        10'b0001110110: data <= 18'h00053; 
        10'b0001110111: data <= 18'h3fff1; 
        10'b0001111000: data <= 18'h3ff96; 
        10'b0001111001: data <= 18'h00028; 
        10'b0001111010: data <= 18'h3ff51; 
        10'b0001111011: data <= 18'h3ff09; 
        10'b0001111100: data <= 18'h3fea5; 
        10'b0001111101: data <= 18'h3fd8a; 
        10'b0001111110: data <= 18'h3fcdf; 
        10'b0001111111: data <= 18'h3fbd1; 
        10'b0010000000: data <= 18'h3fce8; 
        10'b0010000001: data <= 18'h3fce6; 
        10'b0010000010: data <= 18'h3fdb1; 
        10'b0010000011: data <= 18'h3fefc; 
        10'b0010000100: data <= 18'h3ff86; 
        10'b0010000101: data <= 18'h3ffa8; 
        10'b0010000110: data <= 18'h0001d; 
        10'b0010000111: data <= 18'h00095; 
        10'b0010001000: data <= 18'h00075; 
        10'b0010001001: data <= 18'h0006c; 
        10'b0010001010: data <= 18'h00001; 
        10'b0010001011: data <= 18'h00005; 
        10'b0010001100: data <= 18'h00091; 
        10'b0010001101: data <= 18'h00067; 
        10'b0010001110: data <= 18'h00078; 
        10'b0010001111: data <= 18'h0004c; 
        10'b0010010000: data <= 18'h0005c; 
        10'b0010010001: data <= 18'h3ff8e; 
        10'b0010010010: data <= 18'h3ff9a; 
        10'b0010010011: data <= 18'h3ff8f; 
        10'b0010010100: data <= 18'h3fe94; 
        10'b0010010101: data <= 18'h3fe9c; 
        10'b0010010110: data <= 18'h3fe7f; 
        10'b0010010111: data <= 18'h3fe05; 
        10'b0010011000: data <= 18'h3fd85; 
        10'b0010011001: data <= 18'h3fd11; 
        10'b0010011010: data <= 18'h3fb85; 
        10'b0010011011: data <= 18'h3fb2a; 
        10'b0010011100: data <= 18'h3f9e3; 
        10'b0010011101: data <= 18'h3fbf8; 
        10'b0010011110: data <= 18'h3fd76; 
        10'b0010011111: data <= 18'h3fec5; 
        10'b0010100000: data <= 18'h3feb4; 
        10'b0010100001: data <= 18'h3fe4f; 
        10'b0010100010: data <= 18'h3fe6d; 
        10'b0010100011: data <= 18'h3fee1; 
        10'b0010100100: data <= 18'h3ff8e; 
        10'b0010100101: data <= 18'h3ffcb; 
        10'b0010100110: data <= 18'h00012; 
        10'b0010100111: data <= 18'h00065; 
        10'b0010101000: data <= 18'h00082; 
        10'b0010101001: data <= 18'h00086; 
        10'b0010101010: data <= 18'h3ffac; 
        10'b0010101011: data <= 18'h00087; 
        10'b0010101100: data <= 18'h00056; 
        10'b0010101101: data <= 18'h3fe7d; 
        10'b0010101110: data <= 18'h3fe29; 
        10'b0010101111: data <= 18'h3fdd5; 
        10'b0010110000: data <= 18'h3fd8f; 
        10'b0010110001: data <= 18'h3fd01; 
        10'b0010110010: data <= 18'h3fdcd; 
        10'b0010110011: data <= 18'h3ff4c; 
        10'b0010110100: data <= 18'h0002d; 
        10'b0010110101: data <= 18'h002b5; 
        10'b0010110110: data <= 18'h00409; 
        10'b0010110111: data <= 18'h00336; 
        10'b0010111000: data <= 18'h00240; 
        10'b0010111001: data <= 18'h001de; 
        10'b0010111010: data <= 18'h0025f; 
        10'b0010111011: data <= 18'h3ff9a; 
        10'b0010111100: data <= 18'h3ff6e; 
        10'b0010111101: data <= 18'h3fe32; 
        10'b0010111110: data <= 18'h3fcc5; 
        10'b0010111111: data <= 18'h3fcfe; 
        10'b0011000000: data <= 18'h3fe47; 
        10'b0011000001: data <= 18'h3ff29; 
        10'b0011000010: data <= 18'h3ffdf; 
        10'b0011000011: data <= 18'h00046; 
        10'b0011000100: data <= 18'h000c7; 
        10'b0011000101: data <= 18'h3fff9; 
        10'b0011000110: data <= 18'h3ffbf; 
        10'b0011000111: data <= 18'h3ffb8; 
        10'b0011001000: data <= 18'h3fe46; 
        10'b0011001001: data <= 18'h3fd60; 
        10'b0011001010: data <= 18'h3fce8; 
        10'b0011001011: data <= 18'h3fc52; 
        10'b0011001100: data <= 18'h3fc85; 
        10'b0011001101: data <= 18'h3fec6; 
        10'b0011001110: data <= 18'h3ffe6; 
        10'b0011001111: data <= 18'h000f4; 
        10'b0011010000: data <= 18'h003ab; 
        10'b0011010001: data <= 18'h00460; 
        10'b0011010010: data <= 18'h00600; 
        10'b0011010011: data <= 18'h00608; 
        10'b0011010100: data <= 18'h00646; 
        10'b0011010101: data <= 18'h002d8; 
        10'b0011010110: data <= 18'h00224; 
        10'b0011010111: data <= 18'h0003b; 
        10'b0011011000: data <= 18'h0008e; 
        10'b0011011001: data <= 18'h000a1; 
        10'b0011011010: data <= 18'h3fdd7; 
        10'b0011011011: data <= 18'h3fc21; 
        10'b0011011100: data <= 18'h3fdb8; 
        10'b0011011101: data <= 18'h3ff6e; 
        10'b0011011110: data <= 18'h3ff6a; 
        10'b0011011111: data <= 18'h00083; 
        10'b0011100000: data <= 18'h000c2; 
        10'b0011100001: data <= 18'h000c3; 
        10'b0011100010: data <= 18'h00063; 
        10'b0011100011: data <= 18'h3ffc4; 
        10'b0011100100: data <= 18'h3fe34; 
        10'b0011100101: data <= 18'h3fd47; 
        10'b0011100110: data <= 18'h3fcd5; 
        10'b0011100111: data <= 18'h3fb92; 
        10'b0011101000: data <= 18'h3fed4; 
        10'b0011101001: data <= 18'h3ff75; 
        10'b0011101010: data <= 18'h3ff5f; 
        10'b0011101011: data <= 18'h3febd; 
        10'b0011101100: data <= 18'h3ffe7; 
        10'b0011101101: data <= 18'h001c2; 
        10'b0011101110: data <= 18'h00524; 
        10'b0011101111: data <= 18'h002d7; 
        10'b0011110000: data <= 18'h002e4; 
        10'b0011110001: data <= 18'h00097; 
        10'b0011110010: data <= 18'h0003a; 
        10'b0011110011: data <= 18'h00027; 
        10'b0011110100: data <= 18'h3ff0d; 
        10'b0011110101: data <= 18'h0007e; 
        10'b0011110110: data <= 18'h3fec8; 
        10'b0011110111: data <= 18'h3fce9; 
        10'b0011111000: data <= 18'h3fd64; 
        10'b0011111001: data <= 18'h3fec0; 
        10'b0011111010: data <= 18'h3ff74; 
        10'b0011111011: data <= 18'h000b5; 
        10'b0011111100: data <= 18'h0003b; 
        10'b0011111101: data <= 18'h00023; 
        10'b0011111110: data <= 18'h0000d; 
        10'b0011111111: data <= 18'h3feb7; 
        10'b0100000000: data <= 18'h3fd32; 
        10'b0100000001: data <= 18'h3fdd9; 
        10'b0100000010: data <= 18'h3ff64; 
        10'b0100000011: data <= 18'h3fec4; 
        10'b0100000100: data <= 18'h3ff44; 
        10'b0100000101: data <= 18'h3ffab; 
        10'b0100000110: data <= 18'h00151; 
        10'b0100000111: data <= 18'h000cb; 
        10'b0100001000: data <= 18'h0003c; 
        10'b0100001001: data <= 18'h00220; 
        10'b0100001010: data <= 18'h0038e; 
        10'b0100001011: data <= 18'h0032c; 
        10'b0100001100: data <= 18'h3ffe0; 
        10'b0100001101: data <= 18'h3ff17; 
        10'b0100001110: data <= 18'h00009; 
        10'b0100001111: data <= 18'h3fe1b; 
        10'b0100010000: data <= 18'h3ff32; 
        10'b0100010001: data <= 18'h3fe04; 
        10'b0100010010: data <= 18'h3fde0; 
        10'b0100010011: data <= 18'h3fdbc; 
        10'b0100010100: data <= 18'h3fe74; 
        10'b0100010101: data <= 18'h3ff53; 
        10'b0100010110: data <= 18'h3ff82; 
        10'b0100010111: data <= 18'h000a0; 
        10'b0100011000: data <= 18'h00023; 
        10'b0100011001: data <= 18'h3fff9; 
        10'b0100011010: data <= 18'h3ffb3; 
        10'b0100011011: data <= 18'h3ff82; 
        10'b0100011100: data <= 18'h3fdd7; 
        10'b0100011101: data <= 18'h3fedf; 
        10'b0100011110: data <= 18'h0010e; 
        10'b0100011111: data <= 18'h00161; 
        10'b0100100000: data <= 18'h002cd; 
        10'b0100100001: data <= 18'h002c8; 
        10'b0100100010: data <= 18'h00265; 
        10'b0100100011: data <= 18'h0039b; 
        10'b0100100100: data <= 18'h001d1; 
        10'b0100100101: data <= 18'h0006d; 
        10'b0100100110: data <= 18'h00077; 
        10'b0100100111: data <= 18'h3fe2d; 
        10'b0100101000: data <= 18'h3fee9; 
        10'b0100101001: data <= 18'h3ffc9; 
        10'b0100101010: data <= 18'h00145; 
        10'b0100101011: data <= 18'h3fff9; 
        10'b0100101100: data <= 18'h00106; 
        10'b0100101101: data <= 18'h3ff64; 
        10'b0100101110: data <= 18'h3febf; 
        10'b0100101111: data <= 18'h3fed1; 
        10'b0100110000: data <= 18'h3fe7f; 
        10'b0100110001: data <= 18'h3ff92; 
        10'b0100110010: data <= 18'h3ff6e; 
        10'b0100110011: data <= 18'h0005c; 
        10'b0100110100: data <= 18'h3ffe2; 
        10'b0100110101: data <= 18'h00025; 
        10'b0100110110: data <= 18'h3ffad; 
        10'b0100110111: data <= 18'h3ffcb; 
        10'b0100111000: data <= 18'h3ff68; 
        10'b0100111001: data <= 18'h001fd; 
        10'b0100111010: data <= 18'h00499; 
        10'b0100111011: data <= 18'h0036f; 
        10'b0100111100: data <= 18'h00564; 
        10'b0100111101: data <= 18'h00229; 
        10'b0100111110: data <= 18'h0023e; 
        10'b0100111111: data <= 18'h003da; 
        10'b0101000000: data <= 18'h3fec6; 
        10'b0101000001: data <= 18'h3fef5; 
        10'b0101000010: data <= 18'h3ff70; 
        10'b0101000011: data <= 18'h00046; 
        10'b0101000100: data <= 18'h0017d; 
        10'b0101000101: data <= 18'h00536; 
        10'b0101000110: data <= 18'h00276; 
        10'b0101000111: data <= 18'h0027f; 
        10'b0101001000: data <= 18'h00418; 
        10'b0101001001: data <= 18'h002f6; 
        10'b0101001010: data <= 18'h001bb; 
        10'b0101001011: data <= 18'h0005c; 
        10'b0101001100: data <= 18'h3ffb8; 
        10'b0101001101: data <= 18'h3ff4b; 
        10'b0101001110: data <= 18'h3fff8; 
        10'b0101001111: data <= 18'h00001; 
        10'b0101010000: data <= 18'h00053; 
        10'b0101010001: data <= 18'h000ac; 
        10'b0101010010: data <= 18'h3ff8a; 
        10'b0101010011: data <= 18'h3ff43; 
        10'b0101010100: data <= 18'h001ad; 
        10'b0101010101: data <= 18'h0045c; 
        10'b0101010110: data <= 18'h0050b; 
        10'b0101010111: data <= 18'h002fe; 
        10'b0101011000: data <= 18'h003bd; 
        10'b0101011001: data <= 18'h00493; 
        10'b0101011010: data <= 18'h002ec; 
        10'b0101011011: data <= 18'h00009; 
        10'b0101011100: data <= 18'h3fd12; 
        10'b0101011101: data <= 18'h0028a; 
        10'b0101011110: data <= 18'h0057c; 
        10'b0101011111: data <= 18'h00457; 
        10'b0101100000: data <= 18'h003b6; 
        10'b0101100001: data <= 18'h005ac; 
        10'b0101100010: data <= 18'h005b6; 
        10'b0101100011: data <= 18'h005ed; 
        10'b0101100100: data <= 18'h00618; 
        10'b0101100101: data <= 18'h00412; 
        10'b0101100110: data <= 18'h001f5; 
        10'b0101100111: data <= 18'h0000d; 
        10'b0101101000: data <= 18'h3ff18; 
        10'b0101101001: data <= 18'h00026; 
        10'b0101101010: data <= 18'h00054; 
        10'b0101101011: data <= 18'h0005b; 
        10'b0101101100: data <= 18'h000c1; 
        10'b0101101101: data <= 18'h00077; 
        10'b0101101110: data <= 18'h3ff5e; 
        10'b0101101111: data <= 18'h0003d; 
        10'b0101110000: data <= 18'h00289; 
        10'b0101110001: data <= 18'h003d1; 
        10'b0101110010: data <= 18'h00398; 
        10'b0101110011: data <= 18'h0025c; 
        10'b0101110100: data <= 18'h002f7; 
        10'b0101110101: data <= 18'h001e7; 
        10'b0101110110: data <= 18'h001b8; 
        10'b0101110111: data <= 18'h3ff1c; 
        10'b0101111000: data <= 18'h3fe76; 
        10'b0101111001: data <= 18'h003fd; 
        10'b0101111010: data <= 18'h00579; 
        10'b0101111011: data <= 18'h003f7; 
        10'b0101111100: data <= 18'h00492; 
        10'b0101111101: data <= 18'h00419; 
        10'b0101111110: data <= 18'h0059f; 
        10'b0101111111: data <= 18'h005b8; 
        10'b0110000000: data <= 18'h00478; 
        10'b0110000001: data <= 18'h0029c; 
        10'b0110000010: data <= 18'h00026; 
        10'b0110000011: data <= 18'h3fe39; 
        10'b0110000100: data <= 18'h3fef7; 
        10'b0110000101: data <= 18'h3ffae; 
        10'b0110000110: data <= 18'h00056; 
        10'b0110000111: data <= 18'h00058; 
        10'b0110001000: data <= 18'h00027; 
        10'b0110001001: data <= 18'h00013; 
        10'b0110001010: data <= 18'h00085; 
        10'b0110001011: data <= 18'h00054; 
        10'b0110001100: data <= 18'h00129; 
        10'b0110001101: data <= 18'h00118; 
        10'b0110001110: data <= 18'h002fb; 
        10'b0110001111: data <= 18'h00216; 
        10'b0110010000: data <= 18'h00103; 
        10'b0110010001: data <= 18'h3fffd; 
        10'b0110010010: data <= 18'h0005f; 
        10'b0110010011: data <= 18'h3ffd1; 
        10'b0110010100: data <= 18'h3fee0; 
        10'b0110010101: data <= 18'h0014b; 
        10'b0110010110: data <= 18'h000bc; 
        10'b0110010111: data <= 18'h00380; 
        10'b0110011000: data <= 18'h003b6; 
        10'b0110011001: data <= 18'h003b7; 
        10'b0110011010: data <= 18'h00288; 
        10'b0110011011: data <= 18'h001a0; 
        10'b0110011100: data <= 18'h00208; 
        10'b0110011101: data <= 18'h0000a; 
        10'b0110011110: data <= 18'h3fdf3; 
        10'b0110011111: data <= 18'h3fd06; 
        10'b0110100000: data <= 18'h3fec5; 
        10'b0110100001: data <= 18'h00035; 
        10'b0110100010: data <= 18'h0001e; 
        10'b0110100011: data <= 18'h00024; 
        10'b0110100100: data <= 18'h00092; 
        10'b0110100101: data <= 18'h00085; 
        10'b0110100110: data <= 18'h00058; 
        10'b0110100111: data <= 18'h3ff95; 
        10'b0110101000: data <= 18'h00016; 
        10'b0110101001: data <= 18'h00153; 
        10'b0110101010: data <= 18'h00145; 
        10'b0110101011: data <= 18'h000d7; 
        10'b0110101100: data <= 18'h000db; 
        10'b0110101101: data <= 18'h3fe6e; 
        10'b0110101110: data <= 18'h3ff45; 
        10'b0110101111: data <= 18'h3ff44; 
        10'b0110110000: data <= 18'h3fee7; 
        10'b0110110001: data <= 18'h3ff27; 
        10'b0110110010: data <= 18'h3fef9; 
        10'b0110110011: data <= 18'h003d3; 
        10'b0110110100: data <= 18'h00599; 
        10'b0110110101: data <= 18'h0055d; 
        10'b0110110110: data <= 18'h002af; 
        10'b0110110111: data <= 18'h00042; 
        10'b0110111000: data <= 18'h3fed5; 
        10'b0110111001: data <= 18'h3fced; 
        10'b0110111010: data <= 18'h3fc2a; 
        10'b0110111011: data <= 18'h3fd42; 
        10'b0110111100: data <= 18'h3fec8; 
        10'b0110111101: data <= 18'h00006; 
        10'b0110111110: data <= 18'h00050; 
        10'b0110111111: data <= 18'h3fff5; 
        10'b0111000000: data <= 18'h000a8; 
        10'b0111000001: data <= 18'h0000e; 
        10'b0111000010: data <= 18'h3ff88; 
        10'b0111000011: data <= 18'h3ffe1; 
        10'b0111000100: data <= 18'h0000b; 
        10'b0111000101: data <= 18'h00066; 
        10'b0111000110: data <= 18'h3fefa; 
        10'b0111000111: data <= 18'h000cf; 
        10'b0111001000: data <= 18'h0024d; 
        10'b0111001001: data <= 18'h3ff76; 
        10'b0111001010: data <= 18'h0014e; 
        10'b0111001011: data <= 18'h001da; 
        10'b0111001100: data <= 18'h3ffbf; 
        10'b0111001101: data <= 18'h3fde5; 
        10'b0111001110: data <= 18'h3ffa6; 
        10'b0111001111: data <= 18'h0021f; 
        10'b0111010000: data <= 18'h003d2; 
        10'b0111010001: data <= 18'h003cb; 
        10'b0111010010: data <= 18'h000f3; 
        10'b0111010011: data <= 18'h3fdd8; 
        10'b0111010100: data <= 18'h3fc6b; 
        10'b0111010101: data <= 18'h3fb0d; 
        10'b0111010110: data <= 18'h3fc86; 
        10'b0111010111: data <= 18'h3fd2d; 
        10'b0111011000: data <= 18'h3fe22; 
        10'b0111011001: data <= 18'h00010; 
        10'b0111011010: data <= 18'h3ff98; 
        10'b0111011011: data <= 18'h0005a; 
        10'b0111011100: data <= 18'h00038; 
        10'b0111011101: data <= 18'h3ffdb; 
        10'b0111011110: data <= 18'h3ff7c; 
        10'b0111011111: data <= 18'h3ff40; 
        10'b0111100000: data <= 18'h3fe98; 
        10'b0111100001: data <= 18'h3fe4a; 
        10'b0111100010: data <= 18'h3fe97; 
        10'b0111100011: data <= 18'h000a3; 
        10'b0111100100: data <= 18'h0013d; 
        10'b0111100101: data <= 18'h00169; 
        10'b0111100110: data <= 18'h00227; 
        10'b0111100111: data <= 18'h00322; 
        10'b0111101000: data <= 18'h001e9; 
        10'b0111101001: data <= 18'h000e3; 
        10'b0111101010: data <= 18'h00137; 
        10'b0111101011: data <= 18'h0031d; 
        10'b0111101100: data <= 18'h000ed; 
        10'b0111101101: data <= 18'h3ff5e; 
        10'b0111101110: data <= 18'h3fea0; 
        10'b0111101111: data <= 18'h3fcd7; 
        10'b0111110000: data <= 18'h3fce1; 
        10'b0111110001: data <= 18'h3fca4; 
        10'b0111110010: data <= 18'h3fcd7; 
        10'b0111110011: data <= 18'h3fdac; 
        10'b0111110100: data <= 18'h3fe4e; 
        10'b0111110101: data <= 18'h0002b; 
        10'b0111110110: data <= 18'h0002d; 
        10'b0111110111: data <= 18'h3ffda; 
        10'b0111111000: data <= 18'h0009b; 
        10'b0111111001: data <= 18'h00000; 
        10'b0111111010: data <= 18'h3ffa5; 
        10'b0111111011: data <= 18'h3ffdc; 
        10'b0111111100: data <= 18'h3fec3; 
        10'b0111111101: data <= 18'h3fd29; 
        10'b0111111110: data <= 18'h3fd1b; 
        10'b0111111111: data <= 18'h3fd29; 
        10'b1000000000: data <= 18'h3fecf; 
        10'b1000000001: data <= 18'h00079; 
        10'b1000000010: data <= 18'h0036e; 
        10'b1000000011: data <= 18'h002c6; 
        10'b1000000100: data <= 18'h3fe4f; 
        10'b1000000101: data <= 18'h3fe48; 
        10'b1000000110: data <= 18'h0001b; 
        10'b1000000111: data <= 18'h00210; 
        10'b1000001000: data <= 18'h3febd; 
        10'b1000001001: data <= 18'h3fe8f; 
        10'b1000001010: data <= 18'h3fd4d; 
        10'b1000001011: data <= 18'h3fe60; 
        10'b1000001100: data <= 18'h3fe7a; 
        10'b1000001101: data <= 18'h3fd9f; 
        10'b1000001110: data <= 18'h3fd80; 
        10'b1000001111: data <= 18'h3fd61; 
        10'b1000010000: data <= 18'h3fe26; 
        10'b1000010001: data <= 18'h3ffb5; 
        10'b1000010010: data <= 18'h0000a; 
        10'b1000010011: data <= 18'h0008e; 
        10'b1000010100: data <= 18'h00065; 
        10'b1000010101: data <= 18'h000c9; 
        10'b1000010110: data <= 18'h00024; 
        10'b1000010111: data <= 18'h3ff52; 
        10'b1000011000: data <= 18'h3fedd; 
        10'b1000011001: data <= 18'h3fdfd; 
        10'b1000011010: data <= 18'h3fcd3; 
        10'b1000011011: data <= 18'h3fcbd; 
        10'b1000011100: data <= 18'h3fca0; 
        10'b1000011101: data <= 18'h3fca7; 
        10'b1000011110: data <= 18'h3fc41; 
        10'b1000011111: data <= 18'h3fcd6; 
        10'b1000100000: data <= 18'h3fbe7; 
        10'b1000100001: data <= 18'h3fd23; 
        10'b1000100010: data <= 18'h3fd96; 
        10'b1000100011: data <= 18'h3fd41; 
        10'b1000100100: data <= 18'h3fda1; 
        10'b1000100101: data <= 18'h3ff3a; 
        10'b1000100110: data <= 18'h3fe32; 
        10'b1000100111: data <= 18'h3ff7f; 
        10'b1000101000: data <= 18'h3fecb; 
        10'b1000101001: data <= 18'h3fe92; 
        10'b1000101010: data <= 18'h3fea7; 
        10'b1000101011: data <= 18'h3fecd; 
        10'b1000101100: data <= 18'h3ff3f; 
        10'b1000101101: data <= 18'h00038; 
        10'b1000101110: data <= 18'h3ffc3; 
        10'b1000101111: data <= 18'h00016; 
        10'b1000110000: data <= 18'h3ffda; 
        10'b1000110001: data <= 18'h0001c; 
        10'b1000110010: data <= 18'h00055; 
        10'b1000110011: data <= 18'h00007; 
        10'b1000110100: data <= 18'h3fed3; 
        10'b1000110101: data <= 18'h3fe0f; 
        10'b1000110110: data <= 18'h3fd0f; 
        10'b1000110111: data <= 18'h3fb64; 
        10'b1000111000: data <= 18'h3fab8; 
        10'b1000111001: data <= 18'h3fa14; 
        10'b1000111010: data <= 18'h3f7fb; 
        10'b1000111011: data <= 18'h3f9dd; 
        10'b1000111100: data <= 18'h3fa05; 
        10'b1000111101: data <= 18'h3fe0b; 
        10'b1000111110: data <= 18'h3fd41; 
        10'b1000111111: data <= 18'h3feb6; 
        10'b1001000000: data <= 18'h3fe74; 
        10'b1001000001: data <= 18'h3ff95; 
        10'b1001000010: data <= 18'h3fd5f; 
        10'b1001000011: data <= 18'h3ff22; 
        10'b1001000100: data <= 18'h3fef5; 
        10'b1001000101: data <= 18'h3fe53; 
        10'b1001000110: data <= 18'h3ff87; 
        10'b1001000111: data <= 18'h3ff33; 
        10'b1001001000: data <= 18'h00015; 
        10'b1001001001: data <= 18'h000ab; 
        10'b1001001010: data <= 18'h00067; 
        10'b1001001011: data <= 18'h00020; 
        10'b1001001100: data <= 18'h0000e; 
        10'b1001001101: data <= 18'h00000; 
        10'b1001001110: data <= 18'h000ab; 
        10'b1001001111: data <= 18'h3ff4b; 
        10'b1001010000: data <= 18'h3ff36; 
        10'b1001010001: data <= 18'h3fe16; 
        10'b1001010010: data <= 18'h3fd4c; 
        10'b1001010011: data <= 18'h3fbd4; 
        10'b1001010100: data <= 18'h3fb44; 
        10'b1001010101: data <= 18'h3faca; 
        10'b1001010110: data <= 18'h3fa8a; 
        10'b1001010111: data <= 18'h3fb17; 
        10'b1001011000: data <= 18'h3fcdf; 
        10'b1001011001: data <= 18'h3fce9; 
        10'b1001011010: data <= 18'h3fcdc; 
        10'b1001011011: data <= 18'h3fe33; 
        10'b1001011100: data <= 18'h3fe0c; 
        10'b1001011101: data <= 18'h3fd10; 
        10'b1001011110: data <= 18'h3fc75; 
        10'b1001011111: data <= 18'h3fe80; 
        10'b1001100000: data <= 18'h3ff2a; 
        10'b1001100001: data <= 18'h3ff84; 
        10'b1001100010: data <= 18'h0003d; 
        10'b1001100011: data <= 18'h3ffef; 
        10'b1001100100: data <= 18'h0004d; 
        10'b1001100101: data <= 18'h00069; 
        10'b1001100110: data <= 18'h00006; 
        10'b1001100111: data <= 18'h0000d; 
        10'b1001101000: data <= 18'h00083; 
        10'b1001101001: data <= 18'h00021; 
        10'b1001101010: data <= 18'h00025; 
        10'b1001101011: data <= 18'h0007e; 
        10'b1001101100: data <= 18'h3ffaf; 
        10'b1001101101: data <= 18'h3fe74; 
        10'b1001101110: data <= 18'h3fd87; 
        10'b1001101111: data <= 18'h3fca3; 
        10'b1001110000: data <= 18'h3fd7f; 
        10'b1001110001: data <= 18'h3fd62; 
        10'b1001110010: data <= 18'h3fd25; 
        10'b1001110011: data <= 18'h3fe12; 
        10'b1001110100: data <= 18'h3fdd5; 
        10'b1001110101: data <= 18'h3fd1d; 
        10'b1001110110: data <= 18'h3fd93; 
        10'b1001110111: data <= 18'h3fc9a; 
        10'b1001111000: data <= 18'h3fc3e; 
        10'b1001111001: data <= 18'h3fc51; 
        10'b1001111010: data <= 18'h3fcef; 
        10'b1001111011: data <= 18'h3fd46; 
        10'b1001111100: data <= 18'h3ff41; 
        10'b1001111101: data <= 18'h000eb; 
        10'b1001111110: data <= 18'h00082; 
        10'b1001111111: data <= 18'h000a2; 
        10'b1010000000: data <= 18'h00109; 
        10'b1010000001: data <= 18'h00038; 
        10'b1010000010: data <= 18'h0003e; 
        10'b1010000011: data <= 18'h00061; 
        10'b1010000100: data <= 18'h0009a; 
        10'b1010000101: data <= 18'h00079; 
        10'b1010000110: data <= 18'h0002d; 
        10'b1010000111: data <= 18'h3ffc4; 
        10'b1010001000: data <= 18'h3ff91; 
        10'b1010001001: data <= 18'h3feac; 
        10'b1010001010: data <= 18'h3fe74; 
        10'b1010001011: data <= 18'h3fdf5; 
        10'b1010001100: data <= 18'h3ffd8; 
        10'b1010001101: data <= 18'h3ff2c; 
        10'b1010001110: data <= 18'h3ff57; 
        10'b1010001111: data <= 18'h3fd86; 
        10'b1010010000: data <= 18'h3fdfb; 
        10'b1010010001: data <= 18'h3fd74; 
        10'b1010010010: data <= 18'h3fdd9; 
        10'b1010010011: data <= 18'h3fc53; 
        10'b1010010100: data <= 18'h3fc08; 
        10'b1010010101: data <= 18'h3fc82; 
        10'b1010010110: data <= 18'h3fdd3; 
        10'b1010010111: data <= 18'h3ffca; 
        10'b1010011000: data <= 18'h000da; 
        10'b1010011001: data <= 18'h001fa; 
        10'b1010011010: data <= 18'h002da; 
        10'b1010011011: data <= 18'h00263; 
        10'b1010011100: data <= 18'h0011e; 
        10'b1010011101: data <= 18'h3ffec; 
        10'b1010011110: data <= 18'h000cd; 
        10'b1010011111: data <= 18'h3ffe8; 
        10'b1010100000: data <= 18'h3ffff; 
        10'b1010100001: data <= 18'h3ffaf; 
        10'b1010100010: data <= 18'h3ffea; 
        10'b1010100011: data <= 18'h000ad; 
        10'b1010100100: data <= 18'h0007c; 
        10'b1010100101: data <= 18'h000c3; 
        10'b1010100110: data <= 18'h0008d; 
        10'b1010100111: data <= 18'h000cd; 
        10'b1010101000: data <= 18'h00122; 
        10'b1010101001: data <= 18'h0009d; 
        10'b1010101010: data <= 18'h3ff99; 
        10'b1010101011: data <= 18'h3febb; 
        10'b1010101100: data <= 18'h3ffe9; 
        10'b1010101101: data <= 18'h3fe0d; 
        10'b1010101110: data <= 18'h3fd89; 
        10'b1010101111: data <= 18'h3fd66; 
        10'b1010110000: data <= 18'h3fed2; 
        10'b1010110001: data <= 18'h000db; 
        10'b1010110010: data <= 18'h00176; 
        10'b1010110011: data <= 18'h00183; 
        10'b1010110100: data <= 18'h00373; 
        10'b1010110101: data <= 18'h003b6; 
        10'b1010110110: data <= 18'h00223; 
        10'b1010110111: data <= 18'h0014e; 
        10'b1010111000: data <= 18'h00108; 
        10'b1010111001: data <= 18'h3ffcc; 
        10'b1010111010: data <= 18'h00076; 
        10'b1010111011: data <= 18'h3fff8; 
        10'b1010111100: data <= 18'h0002b; 
        10'b1010111101: data <= 18'h000ab; 
        10'b1010111110: data <= 18'h000ac; 
        10'b1010111111: data <= 18'h3ffee; 
        10'b1011000000: data <= 18'h00010; 
        10'b1011000001: data <= 18'h00125; 
        10'b1011000010: data <= 18'h000de; 
        10'b1011000011: data <= 18'h00281; 
        10'b1011000100: data <= 18'h002bf; 
        10'b1011000101: data <= 18'h002cb; 
        10'b1011000110: data <= 18'h0026b; 
        10'b1011000111: data <= 18'h000f6; 
        10'b1011001000: data <= 18'h0028b; 
        10'b1011001001: data <= 18'h00245; 
        10'b1011001010: data <= 18'h0022c; 
        10'b1011001011: data <= 18'h0020b; 
        10'b1011001100: data <= 18'h003d1; 
        10'b1011001101: data <= 18'h00425; 
        10'b1011001110: data <= 18'h0048f; 
        10'b1011001111: data <= 18'h004c2; 
        10'b1011010000: data <= 18'h00550; 
        10'b1011010001: data <= 18'h003c5; 
        10'b1011010010: data <= 18'h00178; 
        10'b1011010011: data <= 18'h000b3; 
        10'b1011010100: data <= 18'h3ffe8; 
        10'b1011010101: data <= 18'h3fff2; 
        10'b1011010110: data <= 18'h00032; 
        10'b1011010111: data <= 18'h0002a; 
        10'b1011011000: data <= 18'h00007; 
        10'b1011011001: data <= 18'h0009c; 
        10'b1011011010: data <= 18'h0002a; 
        10'b1011011011: data <= 18'h3ffc7; 
        10'b1011011100: data <= 18'h0009d; 
        10'b1011011101: data <= 18'h000f3; 
        10'b1011011110: data <= 18'h00155; 
        10'b1011011111: data <= 18'h001da; 
        10'b1011100000: data <= 18'h0021c; 
        10'b1011100001: data <= 18'h00332; 
        10'b1011100010: data <= 18'h0034c; 
        10'b1011100011: data <= 18'h003b4; 
        10'b1011100100: data <= 18'h00463; 
        10'b1011100101: data <= 18'h0046d; 
        10'b1011100110: data <= 18'h0056b; 
        10'b1011100111: data <= 18'h00320; 
        10'b1011101000: data <= 18'h00224; 
        10'b1011101001: data <= 18'h001cf; 
        10'b1011101010: data <= 18'h002ab; 
        10'b1011101011: data <= 18'h002e1; 
        10'b1011101100: data <= 18'h00217; 
        10'b1011101101: data <= 18'h00175; 
        10'b1011101110: data <= 18'h0009b; 
        10'b1011101111: data <= 18'h00038; 
        10'b1011110000: data <= 18'h00023; 
        10'b1011110001: data <= 18'h0003e; 
        10'b1011110010: data <= 18'h3ffc5; 
        10'b1011110011: data <= 18'h00022; 
        10'b1011110100: data <= 18'h3ffdb; 
        10'b1011110101: data <= 18'h00047; 
        10'b1011110110: data <= 18'h3ffc0; 
        10'b1011110111: data <= 18'h000bd; 
        10'b1011111000: data <= 18'h0006d; 
        10'b1011111001: data <= 18'h0003c; 
        10'b1011111010: data <= 18'h3ffe5; 
        10'b1011111011: data <= 18'h000b8; 
        10'b1011111100: data <= 18'h0009b; 
        10'b1011111101: data <= 18'h0006a; 
        10'b1011111110: data <= 18'h3ffde; 
        10'b1011111111: data <= 18'h3ffda; 
        10'b1100000000: data <= 18'h00025; 
        10'b1100000001: data <= 18'h3ffde; 
        10'b1100000010: data <= 18'h00028; 
        10'b1100000011: data <= 18'h00076; 
        10'b1100000100: data <= 18'h0000b; 
        10'b1100000101: data <= 18'h00040; 
        10'b1100000110: data <= 18'h000d2; 
        10'b1100000111: data <= 18'h000bb; 
        10'b1100001000: data <= 18'h00069; 
        10'b1100001001: data <= 18'h00040; 
        10'b1100001010: data <= 18'h3ffcc; 
        10'b1100001011: data <= 18'h000cf; 
        10'b1100001100: data <= 18'h00071; 
        10'b1100001101: data <= 18'h3ffda; 
        10'b1100001110: data <= 18'h0000e; 
        10'b1100001111: data <= 18'h3ffeb; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 13) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 19'h00121; 
        10'b0000000001: data <= 19'h000fd; 
        10'b0000000010: data <= 19'h7ffb2; 
        10'b0000000011: data <= 19'h000b2; 
        10'b0000000100: data <= 19'h000a4; 
        10'b0000000101: data <= 19'h00109; 
        10'b0000000110: data <= 19'h7ff9d; 
        10'b0000000111: data <= 19'h00031; 
        10'b0000001000: data <= 19'h00132; 
        10'b0000001001: data <= 19'h7ff83; 
        10'b0000001010: data <= 19'h7ffdb; 
        10'b0000001011: data <= 19'h00085; 
        10'b0000001100: data <= 19'h00182; 
        10'b0000001101: data <= 19'h000fb; 
        10'b0000001110: data <= 19'h7ff63; 
        10'b0000001111: data <= 19'h7ffb7; 
        10'b0000010000: data <= 19'h7ffb0; 
        10'b0000010001: data <= 19'h00098; 
        10'b0000010010: data <= 19'h00117; 
        10'b0000010011: data <= 19'h00015; 
        10'b0000010100: data <= 19'h0001c; 
        10'b0000010101: data <= 19'h7ffec; 
        10'b0000010110: data <= 19'h7ff84; 
        10'b0000010111: data <= 19'h0002b; 
        10'b0000011000: data <= 19'h00139; 
        10'b0000011001: data <= 19'h0005f; 
        10'b0000011010: data <= 19'h7ff71; 
        10'b0000011011: data <= 19'h0009b; 
        10'b0000011100: data <= 19'h00103; 
        10'b0000011101: data <= 19'h000d9; 
        10'b0000011110: data <= 19'h00069; 
        10'b0000011111: data <= 19'h7ffc4; 
        10'b0000100000: data <= 19'h7ff6a; 
        10'b0000100001: data <= 19'h7ff85; 
        10'b0000100010: data <= 19'h7ffe7; 
        10'b0000100011: data <= 19'h00184; 
        10'b0000100100: data <= 19'h7ff6e; 
        10'b0000100101: data <= 19'h0013b; 
        10'b0000100110: data <= 19'h00079; 
        10'b0000100111: data <= 19'h000c2; 
        10'b0000101000: data <= 19'h00098; 
        10'b0000101001: data <= 19'h000dc; 
        10'b0000101010: data <= 19'h00006; 
        10'b0000101011: data <= 19'h7ff55; 
        10'b0000101100: data <= 19'h7ffa9; 
        10'b0000101101: data <= 19'h000f0; 
        10'b0000101110: data <= 19'h7fff6; 
        10'b0000101111: data <= 19'h00044; 
        10'b0000110000: data <= 19'h00130; 
        10'b0000110001: data <= 19'h7ffe9; 
        10'b0000110010: data <= 19'h00035; 
        10'b0000110011: data <= 19'h0001c; 
        10'b0000110100: data <= 19'h000a7; 
        10'b0000110101: data <= 19'h00146; 
        10'b0000110110: data <= 19'h7fffc; 
        10'b0000110111: data <= 19'h00045; 
        10'b0000111000: data <= 19'h00157; 
        10'b0000111001: data <= 19'h00160; 
        10'b0000111010: data <= 19'h0001a; 
        10'b0000111011: data <= 19'h000f0; 
        10'b0000111100: data <= 19'h00123; 
        10'b0000111101: data <= 19'h7fff2; 
        10'b0000111110: data <= 19'h7ffde; 
        10'b0000111111: data <= 19'h00068; 
        10'b0001000000: data <= 19'h00124; 
        10'b0001000001: data <= 19'h7ffd6; 
        10'b0001000010: data <= 19'h7ffa7; 
        10'b0001000011: data <= 19'h000df; 
        10'b0001000100: data <= 19'h00084; 
        10'b0001000101: data <= 19'h00117; 
        10'b0001000110: data <= 19'h7ff5c; 
        10'b0001000111: data <= 19'h00126; 
        10'b0001001000: data <= 19'h7ff96; 
        10'b0001001001: data <= 19'h7ff90; 
        10'b0001001010: data <= 19'h0001b; 
        10'b0001001011: data <= 19'h7ff74; 
        10'b0001001100: data <= 19'h00151; 
        10'b0001001101: data <= 19'h7ffa7; 
        10'b0001001110: data <= 19'h7ff87; 
        10'b0001001111: data <= 19'h00150; 
        10'b0001010000: data <= 19'h0003c; 
        10'b0001010001: data <= 19'h0003b; 
        10'b0001010010: data <= 19'h0004b; 
        10'b0001010011: data <= 19'h00096; 
        10'b0001010100: data <= 19'h001a2; 
        10'b0001010101: data <= 19'h0000e; 
        10'b0001010110: data <= 19'h7ffda; 
        10'b0001010111: data <= 19'h0007c; 
        10'b0001011000: data <= 19'h00083; 
        10'b0001011001: data <= 19'h7ff75; 
        10'b0001011010: data <= 19'h00157; 
        10'b0001011011: data <= 19'h000bc; 
        10'b0001011100: data <= 19'h7ffbc; 
        10'b0001011101: data <= 19'h0015a; 
        10'b0001011110: data <= 19'h0006c; 
        10'b0001011111: data <= 19'h00111; 
        10'b0001100000: data <= 19'h7ffe4; 
        10'b0001100001: data <= 19'h7fec8; 
        10'b0001100010: data <= 19'h7ffe4; 
        10'b0001100011: data <= 19'h7fe26; 
        10'b0001100100: data <= 19'h7ffc6; 
        10'b0001100101: data <= 19'h7ff09; 
        10'b0001100110: data <= 19'h00052; 
        10'b0001100111: data <= 19'h00031; 
        10'b0001101000: data <= 19'h0006a; 
        10'b0001101001: data <= 19'h7ffe6; 
        10'b0001101010: data <= 19'h00110; 
        10'b0001101011: data <= 19'h7ffdd; 
        10'b0001101100: data <= 19'h7ffd8; 
        10'b0001101101: data <= 19'h00176; 
        10'b0001101110: data <= 19'h0008b; 
        10'b0001101111: data <= 19'h000ee; 
        10'b0001110000: data <= 19'h0002e; 
        10'b0001110001: data <= 19'h0004d; 
        10'b0001110010: data <= 19'h00013; 
        10'b0001110011: data <= 19'h7ffaf; 
        10'b0001110100: data <= 19'h7ff7b; 
        10'b0001110101: data <= 19'h000f1; 
        10'b0001110110: data <= 19'h000a7; 
        10'b0001110111: data <= 19'h7ffe1; 
        10'b0001111000: data <= 19'h7ff2c; 
        10'b0001111001: data <= 19'h00051; 
        10'b0001111010: data <= 19'h7fea1; 
        10'b0001111011: data <= 19'h7fe12; 
        10'b0001111100: data <= 19'h7fd4a; 
        10'b0001111101: data <= 19'h7fb15; 
        10'b0001111110: data <= 19'h7f9bd; 
        10'b0001111111: data <= 19'h7f7a1; 
        10'b0010000000: data <= 19'h7f9d1; 
        10'b0010000001: data <= 19'h7f9cc; 
        10'b0010000010: data <= 19'h7fb63; 
        10'b0010000011: data <= 19'h7fdf9; 
        10'b0010000100: data <= 19'h7ff0d; 
        10'b0010000101: data <= 19'h7ff51; 
        10'b0010000110: data <= 19'h0003a; 
        10'b0010000111: data <= 19'h0012a; 
        10'b0010001000: data <= 19'h000ea; 
        10'b0010001001: data <= 19'h000d9; 
        10'b0010001010: data <= 19'h00002; 
        10'b0010001011: data <= 19'h0000b; 
        10'b0010001100: data <= 19'h00121; 
        10'b0010001101: data <= 19'h000cd; 
        10'b0010001110: data <= 19'h000f0; 
        10'b0010001111: data <= 19'h00098; 
        10'b0010010000: data <= 19'h000b8; 
        10'b0010010001: data <= 19'h7ff1c; 
        10'b0010010010: data <= 19'h7ff35; 
        10'b0010010011: data <= 19'h7ff1f; 
        10'b0010010100: data <= 19'h7fd29; 
        10'b0010010101: data <= 19'h7fd37; 
        10'b0010010110: data <= 19'h7fcfe; 
        10'b0010010111: data <= 19'h7fc0a; 
        10'b0010011000: data <= 19'h7fb0a; 
        10'b0010011001: data <= 19'h7fa21; 
        10'b0010011010: data <= 19'h7f70a; 
        10'b0010011011: data <= 19'h7f653; 
        10'b0010011100: data <= 19'h7f3c6; 
        10'b0010011101: data <= 19'h7f7f1; 
        10'b0010011110: data <= 19'h7faec; 
        10'b0010011111: data <= 19'h7fd8a; 
        10'b0010100000: data <= 19'h7fd67; 
        10'b0010100001: data <= 19'h7fc9e; 
        10'b0010100010: data <= 19'h7fcda; 
        10'b0010100011: data <= 19'h7fdc1; 
        10'b0010100100: data <= 19'h7ff1b; 
        10'b0010100101: data <= 19'h7ff96; 
        10'b0010100110: data <= 19'h00023; 
        10'b0010100111: data <= 19'h000cb; 
        10'b0010101000: data <= 19'h00104; 
        10'b0010101001: data <= 19'h0010b; 
        10'b0010101010: data <= 19'h7ff58; 
        10'b0010101011: data <= 19'h0010e; 
        10'b0010101100: data <= 19'h000ac; 
        10'b0010101101: data <= 19'h7fcfa; 
        10'b0010101110: data <= 19'h7fc52; 
        10'b0010101111: data <= 19'h7fbab; 
        10'b0010110000: data <= 19'h7fb1d; 
        10'b0010110001: data <= 19'h7fa02; 
        10'b0010110010: data <= 19'h7fb99; 
        10'b0010110011: data <= 19'h7fe98; 
        10'b0010110100: data <= 19'h0005b; 
        10'b0010110101: data <= 19'h00569; 
        10'b0010110110: data <= 19'h00812; 
        10'b0010110111: data <= 19'h0066c; 
        10'b0010111000: data <= 19'h00480; 
        10'b0010111001: data <= 19'h003bd; 
        10'b0010111010: data <= 19'h004be; 
        10'b0010111011: data <= 19'h7ff33; 
        10'b0010111100: data <= 19'h7fedc; 
        10'b0010111101: data <= 19'h7fc65; 
        10'b0010111110: data <= 19'h7f989; 
        10'b0010111111: data <= 19'h7f9fc; 
        10'b0011000000: data <= 19'h7fc8e; 
        10'b0011000001: data <= 19'h7fe53; 
        10'b0011000010: data <= 19'h7ffbf; 
        10'b0011000011: data <= 19'h0008c; 
        10'b0011000100: data <= 19'h0018f; 
        10'b0011000101: data <= 19'h7fff2; 
        10'b0011000110: data <= 19'h7ff7e; 
        10'b0011000111: data <= 19'h7ff70; 
        10'b0011001000: data <= 19'h7fc8b; 
        10'b0011001001: data <= 19'h7fabf; 
        10'b0011001010: data <= 19'h7f9d0; 
        10'b0011001011: data <= 19'h7f8a3; 
        10'b0011001100: data <= 19'h7f909; 
        10'b0011001101: data <= 19'h7fd8b; 
        10'b0011001110: data <= 19'h7ffcd; 
        10'b0011001111: data <= 19'h001e8; 
        10'b0011010000: data <= 19'h00755; 
        10'b0011010001: data <= 19'h008c1; 
        10'b0011010010: data <= 19'h00c00; 
        10'b0011010011: data <= 19'h00c10; 
        10'b0011010100: data <= 19'h00c8d; 
        10'b0011010101: data <= 19'h005b0; 
        10'b0011010110: data <= 19'h00448; 
        10'b0011010111: data <= 19'h00077; 
        10'b0011011000: data <= 19'h0011d; 
        10'b0011011001: data <= 19'h00142; 
        10'b0011011010: data <= 19'h7fbad; 
        10'b0011011011: data <= 19'h7f842; 
        10'b0011011100: data <= 19'h7fb70; 
        10'b0011011101: data <= 19'h7fedc; 
        10'b0011011110: data <= 19'h7fed5; 
        10'b0011011111: data <= 19'h00106; 
        10'b0011100000: data <= 19'h00183; 
        10'b0011100001: data <= 19'h00186; 
        10'b0011100010: data <= 19'h000c6; 
        10'b0011100011: data <= 19'h7ff89; 
        10'b0011100100: data <= 19'h7fc67; 
        10'b0011100101: data <= 19'h7fa8e; 
        10'b0011100110: data <= 19'h7f9a9; 
        10'b0011100111: data <= 19'h7f723; 
        10'b0011101000: data <= 19'h7fda8; 
        10'b0011101001: data <= 19'h7feea; 
        10'b0011101010: data <= 19'h7febf; 
        10'b0011101011: data <= 19'h7fd7a; 
        10'b0011101100: data <= 19'h7ffcf; 
        10'b0011101101: data <= 19'h00383; 
        10'b0011101110: data <= 19'h00a49; 
        10'b0011101111: data <= 19'h005ad; 
        10'b0011110000: data <= 19'h005c8; 
        10'b0011110001: data <= 19'h0012f; 
        10'b0011110010: data <= 19'h00075; 
        10'b0011110011: data <= 19'h0004e; 
        10'b0011110100: data <= 19'h7fe19; 
        10'b0011110101: data <= 19'h000fd; 
        10'b0011110110: data <= 19'h7fd91; 
        10'b0011110111: data <= 19'h7f9d3; 
        10'b0011111000: data <= 19'h7fac8; 
        10'b0011111001: data <= 19'h7fd80; 
        10'b0011111010: data <= 19'h7fee8; 
        10'b0011111011: data <= 19'h00169; 
        10'b0011111100: data <= 19'h00075; 
        10'b0011111101: data <= 19'h00046; 
        10'b0011111110: data <= 19'h0001a; 
        10'b0011111111: data <= 19'h7fd6e; 
        10'b0100000000: data <= 19'h7fa64; 
        10'b0100000001: data <= 19'h7fbb3; 
        10'b0100000010: data <= 19'h7fec8; 
        10'b0100000011: data <= 19'h7fd89; 
        10'b0100000100: data <= 19'h7fe88; 
        10'b0100000101: data <= 19'h7ff56; 
        10'b0100000110: data <= 19'h002a3; 
        10'b0100000111: data <= 19'h00197; 
        10'b0100001000: data <= 19'h00077; 
        10'b0100001001: data <= 19'h0043f; 
        10'b0100001010: data <= 19'h0071d; 
        10'b0100001011: data <= 19'h00657; 
        10'b0100001100: data <= 19'h7ffc1; 
        10'b0100001101: data <= 19'h7fe2f; 
        10'b0100001110: data <= 19'h00012; 
        10'b0100001111: data <= 19'h7fc37; 
        10'b0100010000: data <= 19'h7fe65; 
        10'b0100010001: data <= 19'h7fc08; 
        10'b0100010010: data <= 19'h7fbc0; 
        10'b0100010011: data <= 19'h7fb77; 
        10'b0100010100: data <= 19'h7fce9; 
        10'b0100010101: data <= 19'h7fea6; 
        10'b0100010110: data <= 19'h7ff05; 
        10'b0100010111: data <= 19'h00141; 
        10'b0100011000: data <= 19'h00045; 
        10'b0100011001: data <= 19'h7fff2; 
        10'b0100011010: data <= 19'h7ff65; 
        10'b0100011011: data <= 19'h7ff04; 
        10'b0100011100: data <= 19'h7fbae; 
        10'b0100011101: data <= 19'h7fdbe; 
        10'b0100011110: data <= 19'h0021b; 
        10'b0100011111: data <= 19'h002c3; 
        10'b0100100000: data <= 19'h0059a; 
        10'b0100100001: data <= 19'h00590; 
        10'b0100100010: data <= 19'h004ca; 
        10'b0100100011: data <= 19'h00736; 
        10'b0100100100: data <= 19'h003a1; 
        10'b0100100101: data <= 19'h000db; 
        10'b0100100110: data <= 19'h000ed; 
        10'b0100100111: data <= 19'h7fc5a; 
        10'b0100101000: data <= 19'h7fdd3; 
        10'b0100101001: data <= 19'h7ff92; 
        10'b0100101010: data <= 19'h0028b; 
        10'b0100101011: data <= 19'h7fff2; 
        10'b0100101100: data <= 19'h0020c; 
        10'b0100101101: data <= 19'h7fec7; 
        10'b0100101110: data <= 19'h7fd7e; 
        10'b0100101111: data <= 19'h7fda2; 
        10'b0100110000: data <= 19'h7fcfe; 
        10'b0100110001: data <= 19'h7ff24; 
        10'b0100110010: data <= 19'h7fedd; 
        10'b0100110011: data <= 19'h000b8; 
        10'b0100110100: data <= 19'h7ffc3; 
        10'b0100110101: data <= 19'h0004a; 
        10'b0100110110: data <= 19'h7ff5a; 
        10'b0100110111: data <= 19'h7ff96; 
        10'b0100111000: data <= 19'h7fed1; 
        10'b0100111001: data <= 19'h003fa; 
        10'b0100111010: data <= 19'h00932; 
        10'b0100111011: data <= 19'h006dd; 
        10'b0100111100: data <= 19'h00ac9; 
        10'b0100111101: data <= 19'h00453; 
        10'b0100111110: data <= 19'h0047c; 
        10'b0100111111: data <= 19'h007b3; 
        10'b0101000000: data <= 19'h7fd8d; 
        10'b0101000001: data <= 19'h7fdeb; 
        10'b0101000010: data <= 19'h7fee0; 
        10'b0101000011: data <= 19'h0008b; 
        10'b0101000100: data <= 19'h002fa; 
        10'b0101000101: data <= 19'h00a6c; 
        10'b0101000110: data <= 19'h004ec; 
        10'b0101000111: data <= 19'h004fe; 
        10'b0101001000: data <= 19'h0082f; 
        10'b0101001001: data <= 19'h005ec; 
        10'b0101001010: data <= 19'h00376; 
        10'b0101001011: data <= 19'h000b7; 
        10'b0101001100: data <= 19'h7ff6f; 
        10'b0101001101: data <= 19'h7fe97; 
        10'b0101001110: data <= 19'h7fff0; 
        10'b0101001111: data <= 19'h00002; 
        10'b0101010000: data <= 19'h000a7; 
        10'b0101010001: data <= 19'h00157; 
        10'b0101010010: data <= 19'h7ff13; 
        10'b0101010011: data <= 19'h7fe86; 
        10'b0101010100: data <= 19'h0035b; 
        10'b0101010101: data <= 19'h008b8; 
        10'b0101010110: data <= 19'h00a17; 
        10'b0101010111: data <= 19'h005fc; 
        10'b0101011000: data <= 19'h0077b; 
        10'b0101011001: data <= 19'h00925; 
        10'b0101011010: data <= 19'h005d7; 
        10'b0101011011: data <= 19'h00012; 
        10'b0101011100: data <= 19'h7fa24; 
        10'b0101011101: data <= 19'h00514; 
        10'b0101011110: data <= 19'h00af8; 
        10'b0101011111: data <= 19'h008ad; 
        10'b0101100000: data <= 19'h0076b; 
        10'b0101100001: data <= 19'h00b58; 
        10'b0101100010: data <= 19'h00b6c; 
        10'b0101100011: data <= 19'h00bdb; 
        10'b0101100100: data <= 19'h00c30; 
        10'b0101100101: data <= 19'h00825; 
        10'b0101100110: data <= 19'h003eb; 
        10'b0101100111: data <= 19'h0001a; 
        10'b0101101000: data <= 19'h7fe30; 
        10'b0101101001: data <= 19'h0004c; 
        10'b0101101010: data <= 19'h000a8; 
        10'b0101101011: data <= 19'h000b6; 
        10'b0101101100: data <= 19'h00182; 
        10'b0101101101: data <= 19'h000ed; 
        10'b0101101110: data <= 19'h7febb; 
        10'b0101101111: data <= 19'h0007a; 
        10'b0101110000: data <= 19'h00513; 
        10'b0101110001: data <= 19'h007a1; 
        10'b0101110010: data <= 19'h00731; 
        10'b0101110011: data <= 19'h004b8; 
        10'b0101110100: data <= 19'h005ed; 
        10'b0101110101: data <= 19'h003ce; 
        10'b0101110110: data <= 19'h00370; 
        10'b0101110111: data <= 19'h7fe38; 
        10'b0101111000: data <= 19'h7fcec; 
        10'b0101111001: data <= 19'h007fb; 
        10'b0101111010: data <= 19'h00af2; 
        10'b0101111011: data <= 19'h007ee; 
        10'b0101111100: data <= 19'h00923; 
        10'b0101111101: data <= 19'h00831; 
        10'b0101111110: data <= 19'h00b3d; 
        10'b0101111111: data <= 19'h00b6f; 
        10'b0110000000: data <= 19'h008f0; 
        10'b0110000001: data <= 19'h00538; 
        10'b0110000010: data <= 19'h0004d; 
        10'b0110000011: data <= 19'h7fc72; 
        10'b0110000100: data <= 19'h7fdee; 
        10'b0110000101: data <= 19'h7ff5b; 
        10'b0110000110: data <= 19'h000ad; 
        10'b0110000111: data <= 19'h000af; 
        10'b0110001000: data <= 19'h0004e; 
        10'b0110001001: data <= 19'h00026; 
        10'b0110001010: data <= 19'h0010a; 
        10'b0110001011: data <= 19'h000a9; 
        10'b0110001100: data <= 19'h00252; 
        10'b0110001101: data <= 19'h00230; 
        10'b0110001110: data <= 19'h005f5; 
        10'b0110001111: data <= 19'h0042b; 
        10'b0110010000: data <= 19'h00207; 
        10'b0110010001: data <= 19'h7fffa; 
        10'b0110010010: data <= 19'h000be; 
        10'b0110010011: data <= 19'h7ffa1; 
        10'b0110010100: data <= 19'h7fdc0; 
        10'b0110010101: data <= 19'h00296; 
        10'b0110010110: data <= 19'h00178; 
        10'b0110010111: data <= 19'h00700; 
        10'b0110011000: data <= 19'h0076c; 
        10'b0110011001: data <= 19'h0076f; 
        10'b0110011010: data <= 19'h00510; 
        10'b0110011011: data <= 19'h00341; 
        10'b0110011100: data <= 19'h0040f; 
        10'b0110011101: data <= 19'h00013; 
        10'b0110011110: data <= 19'h7fbe7; 
        10'b0110011111: data <= 19'h7fa0c; 
        10'b0110100000: data <= 19'h7fd89; 
        10'b0110100001: data <= 19'h00069; 
        10'b0110100010: data <= 19'h0003c; 
        10'b0110100011: data <= 19'h00047; 
        10'b0110100100: data <= 19'h00124; 
        10'b0110100101: data <= 19'h0010a; 
        10'b0110100110: data <= 19'h000b0; 
        10'b0110100111: data <= 19'h7ff2b; 
        10'b0110101000: data <= 19'h0002c; 
        10'b0110101001: data <= 19'h002a6; 
        10'b0110101010: data <= 19'h0028a; 
        10'b0110101011: data <= 19'h001ad; 
        10'b0110101100: data <= 19'h001b6; 
        10'b0110101101: data <= 19'h7fcdc; 
        10'b0110101110: data <= 19'h7fe8a; 
        10'b0110101111: data <= 19'h7fe88; 
        10'b0110110000: data <= 19'h7fdcf; 
        10'b0110110001: data <= 19'h7fe4e; 
        10'b0110110010: data <= 19'h7fdf1; 
        10'b0110110011: data <= 19'h007a5; 
        10'b0110110100: data <= 19'h00b31; 
        10'b0110110101: data <= 19'h00aba; 
        10'b0110110110: data <= 19'h0055f; 
        10'b0110110111: data <= 19'h00085; 
        10'b0110111000: data <= 19'h7fdab; 
        10'b0110111001: data <= 19'h7f9d9; 
        10'b0110111010: data <= 19'h7f854; 
        10'b0110111011: data <= 19'h7fa85; 
        10'b0110111100: data <= 19'h7fd90; 
        10'b0110111101: data <= 19'h0000c; 
        10'b0110111110: data <= 19'h000a0; 
        10'b0110111111: data <= 19'h7ffe9; 
        10'b0111000000: data <= 19'h00150; 
        10'b0111000001: data <= 19'h0001c; 
        10'b0111000010: data <= 19'h7ff0f; 
        10'b0111000011: data <= 19'h7ffc2; 
        10'b0111000100: data <= 19'h00015; 
        10'b0111000101: data <= 19'h000cb; 
        10'b0111000110: data <= 19'h7fdf3; 
        10'b0111000111: data <= 19'h0019f; 
        10'b0111001000: data <= 19'h0049a; 
        10'b0111001001: data <= 19'h7feec; 
        10'b0111001010: data <= 19'h0029c; 
        10'b0111001011: data <= 19'h003b3; 
        10'b0111001100: data <= 19'h7ff7f; 
        10'b0111001101: data <= 19'h7fbca; 
        10'b0111001110: data <= 19'h7ff4c; 
        10'b0111001111: data <= 19'h0043f; 
        10'b0111010000: data <= 19'h007a3; 
        10'b0111010001: data <= 19'h00797; 
        10'b0111010010: data <= 19'h001e5; 
        10'b0111010011: data <= 19'h7fbaf; 
        10'b0111010100: data <= 19'h7f8d7; 
        10'b0111010101: data <= 19'h7f619; 
        10'b0111010110: data <= 19'h7f90d; 
        10'b0111010111: data <= 19'h7fa5a; 
        10'b0111011000: data <= 19'h7fc43; 
        10'b0111011001: data <= 19'h00020; 
        10'b0111011010: data <= 19'h7ff2f; 
        10'b0111011011: data <= 19'h000b5; 
        10'b0111011100: data <= 19'h0006f; 
        10'b0111011101: data <= 19'h7ffb6; 
        10'b0111011110: data <= 19'h7fef9; 
        10'b0111011111: data <= 19'h7fe7f; 
        10'b0111100000: data <= 19'h7fd30; 
        10'b0111100001: data <= 19'h7fc94; 
        10'b0111100010: data <= 19'h7fd2e; 
        10'b0111100011: data <= 19'h00146; 
        10'b0111100100: data <= 19'h0027a; 
        10'b0111100101: data <= 19'h002d2; 
        10'b0111100110: data <= 19'h0044e; 
        10'b0111100111: data <= 19'h00643; 
        10'b0111101000: data <= 19'h003d2; 
        10'b0111101001: data <= 19'h001c6; 
        10'b0111101010: data <= 19'h0026d; 
        10'b0111101011: data <= 19'h0063b; 
        10'b0111101100: data <= 19'h001da; 
        10'b0111101101: data <= 19'h7febd; 
        10'b0111101110: data <= 19'h7fd3f; 
        10'b0111101111: data <= 19'h7f9ad; 
        10'b0111110000: data <= 19'h7f9c2; 
        10'b0111110001: data <= 19'h7f948; 
        10'b0111110010: data <= 19'h7f9ae; 
        10'b0111110011: data <= 19'h7fb59; 
        10'b0111110100: data <= 19'h7fc9c; 
        10'b0111110101: data <= 19'h00057; 
        10'b0111110110: data <= 19'h00059; 
        10'b0111110111: data <= 19'h7ffb4; 
        10'b0111111000: data <= 19'h00136; 
        10'b0111111001: data <= 19'h7ffff; 
        10'b0111111010: data <= 19'h7ff4b; 
        10'b0111111011: data <= 19'h7ffb8; 
        10'b0111111100: data <= 19'h7fd87; 
        10'b0111111101: data <= 19'h7fa52; 
        10'b0111111110: data <= 19'h7fa36; 
        10'b0111111111: data <= 19'h7fa52; 
        10'b1000000000: data <= 19'h7fd9d; 
        10'b1000000001: data <= 19'h000f2; 
        10'b1000000010: data <= 19'h006dc; 
        10'b1000000011: data <= 19'h0058c; 
        10'b1000000100: data <= 19'h7fc9d; 
        10'b1000000101: data <= 19'h7fc90; 
        10'b1000000110: data <= 19'h00036; 
        10'b1000000111: data <= 19'h0041f; 
        10'b1000001000: data <= 19'h7fd79; 
        10'b1000001001: data <= 19'h7fd1e; 
        10'b1000001010: data <= 19'h7fa9a; 
        10'b1000001011: data <= 19'h7fcc0; 
        10'b1000001100: data <= 19'h7fcf4; 
        10'b1000001101: data <= 19'h7fb3f; 
        10'b1000001110: data <= 19'h7faff; 
        10'b1000001111: data <= 19'h7fac3; 
        10'b1000010000: data <= 19'h7fc4b; 
        10'b1000010001: data <= 19'h7ff69; 
        10'b1000010010: data <= 19'h00013; 
        10'b1000010011: data <= 19'h0011c; 
        10'b1000010100: data <= 19'h000c9; 
        10'b1000010101: data <= 19'h00192; 
        10'b1000010110: data <= 19'h00047; 
        10'b1000010111: data <= 19'h7fea4; 
        10'b1000011000: data <= 19'h7fdbb; 
        10'b1000011001: data <= 19'h7fbfb; 
        10'b1000011010: data <= 19'h7f9a5; 
        10'b1000011011: data <= 19'h7f97b; 
        10'b1000011100: data <= 19'h7f940; 
        10'b1000011101: data <= 19'h7f94e; 
        10'b1000011110: data <= 19'h7f881; 
        10'b1000011111: data <= 19'h7f9ab; 
        10'b1000100000: data <= 19'h7f7ce; 
        10'b1000100001: data <= 19'h7fa45; 
        10'b1000100010: data <= 19'h7fb2c; 
        10'b1000100011: data <= 19'h7fa82; 
        10'b1000100100: data <= 19'h7fb42; 
        10'b1000100101: data <= 19'h7fe74; 
        10'b1000100110: data <= 19'h7fc65; 
        10'b1000100111: data <= 19'h7fefe; 
        10'b1000101000: data <= 19'h7fd96; 
        10'b1000101001: data <= 19'h7fd24; 
        10'b1000101010: data <= 19'h7fd4d; 
        10'b1000101011: data <= 19'h7fd9a; 
        10'b1000101100: data <= 19'h7fe7e; 
        10'b1000101101: data <= 19'h0006f; 
        10'b1000101110: data <= 19'h7ff86; 
        10'b1000101111: data <= 19'h0002b; 
        10'b1000110000: data <= 19'h7ffb4; 
        10'b1000110001: data <= 19'h00038; 
        10'b1000110010: data <= 19'h000ab; 
        10'b1000110011: data <= 19'h0000d; 
        10'b1000110100: data <= 19'h7fda6; 
        10'b1000110101: data <= 19'h7fc1e; 
        10'b1000110110: data <= 19'h7fa1d; 
        10'b1000110111: data <= 19'h7f6c8; 
        10'b1000111000: data <= 19'h7f571; 
        10'b1000111001: data <= 19'h7f427; 
        10'b1000111010: data <= 19'h7eff7; 
        10'b1000111011: data <= 19'h7f3ba; 
        10'b1000111100: data <= 19'h7f40a; 
        10'b1000111101: data <= 19'h7fc16; 
        10'b1000111110: data <= 19'h7fa83; 
        10'b1000111111: data <= 19'h7fd6c; 
        10'b1001000000: data <= 19'h7fce8; 
        10'b1001000001: data <= 19'h7ff2b; 
        10'b1001000010: data <= 19'h7fabe; 
        10'b1001000011: data <= 19'h7fe45; 
        10'b1001000100: data <= 19'h7fdea; 
        10'b1001000101: data <= 19'h7fca6; 
        10'b1001000110: data <= 19'h7ff0e; 
        10'b1001000111: data <= 19'h7fe65; 
        10'b1001001000: data <= 19'h00029; 
        10'b1001001001: data <= 19'h00157; 
        10'b1001001010: data <= 19'h000ce; 
        10'b1001001011: data <= 19'h00041; 
        10'b1001001100: data <= 19'h0001c; 
        10'b1001001101: data <= 19'h00000; 
        10'b1001001110: data <= 19'h00156; 
        10'b1001001111: data <= 19'h7fe95; 
        10'b1001010000: data <= 19'h7fe6b; 
        10'b1001010001: data <= 19'h7fc2c; 
        10'b1001010010: data <= 19'h7fa98; 
        10'b1001010011: data <= 19'h7f7a8; 
        10'b1001010100: data <= 19'h7f687; 
        10'b1001010101: data <= 19'h7f595; 
        10'b1001010110: data <= 19'h7f514; 
        10'b1001010111: data <= 19'h7f62d; 
        10'b1001011000: data <= 19'h7f9be; 
        10'b1001011001: data <= 19'h7f9d3; 
        10'b1001011010: data <= 19'h7f9b9; 
        10'b1001011011: data <= 19'h7fc66; 
        10'b1001011100: data <= 19'h7fc19; 
        10'b1001011101: data <= 19'h7fa20; 
        10'b1001011110: data <= 19'h7f8ea; 
        10'b1001011111: data <= 19'h7fcff; 
        10'b1001100000: data <= 19'h7fe53; 
        10'b1001100001: data <= 19'h7ff09; 
        10'b1001100010: data <= 19'h00079; 
        10'b1001100011: data <= 19'h7ffde; 
        10'b1001100100: data <= 19'h0009a; 
        10'b1001100101: data <= 19'h000d2; 
        10'b1001100110: data <= 19'h0000c; 
        10'b1001100111: data <= 19'h00019; 
        10'b1001101000: data <= 19'h00107; 
        10'b1001101001: data <= 19'h00042; 
        10'b1001101010: data <= 19'h0004a; 
        10'b1001101011: data <= 19'h000fb; 
        10'b1001101100: data <= 19'h7ff5e; 
        10'b1001101101: data <= 19'h7fce8; 
        10'b1001101110: data <= 19'h7fb0e; 
        10'b1001101111: data <= 19'h7f945; 
        10'b1001110000: data <= 19'h7fafe; 
        10'b1001110001: data <= 19'h7fac5; 
        10'b1001110010: data <= 19'h7fa4a; 
        10'b1001110011: data <= 19'h7fc24; 
        10'b1001110100: data <= 19'h7fbaa; 
        10'b1001110101: data <= 19'h7fa3b; 
        10'b1001110110: data <= 19'h7fb27; 
        10'b1001110111: data <= 19'h7f934; 
        10'b1001111000: data <= 19'h7f87b; 
        10'b1001111001: data <= 19'h7f8a1; 
        10'b1001111010: data <= 19'h7f9df; 
        10'b1001111011: data <= 19'h7fa8d; 
        10'b1001111100: data <= 19'h7fe81; 
        10'b1001111101: data <= 19'h001d5; 
        10'b1001111110: data <= 19'h00105; 
        10'b1001111111: data <= 19'h00144; 
        10'b1010000000: data <= 19'h00211; 
        10'b1010000001: data <= 19'h0006f; 
        10'b1010000010: data <= 19'h0007c; 
        10'b1010000011: data <= 19'h000c1; 
        10'b1010000100: data <= 19'h00134; 
        10'b1010000101: data <= 19'h000f2; 
        10'b1010000110: data <= 19'h0005b; 
        10'b1010000111: data <= 19'h7ff87; 
        10'b1010001000: data <= 19'h7ff22; 
        10'b1010001001: data <= 19'h7fd57; 
        10'b1010001010: data <= 19'h7fce9; 
        10'b1010001011: data <= 19'h7fbea; 
        10'b1010001100: data <= 19'h7ffb1; 
        10'b1010001101: data <= 19'h7fe59; 
        10'b1010001110: data <= 19'h7fead; 
        10'b1010001111: data <= 19'h7fb0c; 
        10'b1010010000: data <= 19'h7fbf7; 
        10'b1010010001: data <= 19'h7fae8; 
        10'b1010010010: data <= 19'h7fbb2; 
        10'b1010010011: data <= 19'h7f8a6; 
        10'b1010010100: data <= 19'h7f811; 
        10'b1010010101: data <= 19'h7f904; 
        10'b1010010110: data <= 19'h7fba6; 
        10'b1010010111: data <= 19'h7ff93; 
        10'b1010011000: data <= 19'h001b4; 
        10'b1010011001: data <= 19'h003f4; 
        10'b1010011010: data <= 19'h005b3; 
        10'b1010011011: data <= 19'h004c6; 
        10'b1010011100: data <= 19'h0023c; 
        10'b1010011101: data <= 19'h7ffd9; 
        10'b1010011110: data <= 19'h0019a; 
        10'b1010011111: data <= 19'h7ffd0; 
        10'b1010100000: data <= 19'h7ffff; 
        10'b1010100001: data <= 19'h7ff5e; 
        10'b1010100010: data <= 19'h7ffd5; 
        10'b1010100011: data <= 19'h0015a; 
        10'b1010100100: data <= 19'h000f8; 
        10'b1010100101: data <= 19'h00185; 
        10'b1010100110: data <= 19'h0011b; 
        10'b1010100111: data <= 19'h0019b; 
        10'b1010101000: data <= 19'h00244; 
        10'b1010101001: data <= 19'h00139; 
        10'b1010101010: data <= 19'h7ff31; 
        10'b1010101011: data <= 19'h7fd76; 
        10'b1010101100: data <= 19'h7ffd2; 
        10'b1010101101: data <= 19'h7fc1a; 
        10'b1010101110: data <= 19'h7fb12; 
        10'b1010101111: data <= 19'h7facc; 
        10'b1010110000: data <= 19'h7fda4; 
        10'b1010110001: data <= 19'h001b6; 
        10'b1010110010: data <= 19'h002ec; 
        10'b1010110011: data <= 19'h00305; 
        10'b1010110100: data <= 19'h006e5; 
        10'b1010110101: data <= 19'h0076c; 
        10'b1010110110: data <= 19'h00446; 
        10'b1010110111: data <= 19'h0029c; 
        10'b1010111000: data <= 19'h00210; 
        10'b1010111001: data <= 19'h7ff98; 
        10'b1010111010: data <= 19'h000ec; 
        10'b1010111011: data <= 19'h7fff0; 
        10'b1010111100: data <= 19'h00056; 
        10'b1010111101: data <= 19'h00157; 
        10'b1010111110: data <= 19'h00158; 
        10'b1010111111: data <= 19'h7ffdc; 
        10'b1011000000: data <= 19'h00020; 
        10'b1011000001: data <= 19'h0024b; 
        10'b1011000010: data <= 19'h001bc; 
        10'b1011000011: data <= 19'h00502; 
        10'b1011000100: data <= 19'h0057e; 
        10'b1011000101: data <= 19'h00597; 
        10'b1011000110: data <= 19'h004d6; 
        10'b1011000111: data <= 19'h001ec; 
        10'b1011001000: data <= 19'h00516; 
        10'b1011001001: data <= 19'h0048a; 
        10'b1011001010: data <= 19'h00458; 
        10'b1011001011: data <= 19'h00415; 
        10'b1011001100: data <= 19'h007a1; 
        10'b1011001101: data <= 19'h0084b; 
        10'b1011001110: data <= 19'h0091e; 
        10'b1011001111: data <= 19'h00984; 
        10'b1011010000: data <= 19'h00aa0; 
        10'b1011010001: data <= 19'h0078a; 
        10'b1011010010: data <= 19'h002f1; 
        10'b1011010011: data <= 19'h00165; 
        10'b1011010100: data <= 19'h7ffd0; 
        10'b1011010101: data <= 19'h7ffe3; 
        10'b1011010110: data <= 19'h00064; 
        10'b1011010111: data <= 19'h00054; 
        10'b1011011000: data <= 19'h0000f; 
        10'b1011011001: data <= 19'h00138; 
        10'b1011011010: data <= 19'h00054; 
        10'b1011011011: data <= 19'h7ff8e; 
        10'b1011011100: data <= 19'h0013a; 
        10'b1011011101: data <= 19'h001e6; 
        10'b1011011110: data <= 19'h002aa; 
        10'b1011011111: data <= 19'h003b4; 
        10'b1011100000: data <= 19'h00437; 
        10'b1011100001: data <= 19'h00664; 
        10'b1011100010: data <= 19'h00699; 
        10'b1011100011: data <= 19'h00769; 
        10'b1011100100: data <= 19'h008c6; 
        10'b1011100101: data <= 19'h008da; 
        10'b1011100110: data <= 19'h00ad6; 
        10'b1011100111: data <= 19'h00640; 
        10'b1011101000: data <= 19'h00448; 
        10'b1011101001: data <= 19'h0039e; 
        10'b1011101010: data <= 19'h00555; 
        10'b1011101011: data <= 19'h005c2; 
        10'b1011101100: data <= 19'h0042e; 
        10'b1011101101: data <= 19'h002e9; 
        10'b1011101110: data <= 19'h00136; 
        10'b1011101111: data <= 19'h00070; 
        10'b1011110000: data <= 19'h00046; 
        10'b1011110001: data <= 19'h0007c; 
        10'b1011110010: data <= 19'h7ff8b; 
        10'b1011110011: data <= 19'h00044; 
        10'b1011110100: data <= 19'h7ffb5; 
        10'b1011110101: data <= 19'h0008f; 
        10'b1011110110: data <= 19'h7ff7f; 
        10'b1011110111: data <= 19'h0017a; 
        10'b1011111000: data <= 19'h000d9; 
        10'b1011111001: data <= 19'h00078; 
        10'b1011111010: data <= 19'h7ffca; 
        10'b1011111011: data <= 19'h00170; 
        10'b1011111100: data <= 19'h00137; 
        10'b1011111101: data <= 19'h000d5; 
        10'b1011111110: data <= 19'h7ffbb; 
        10'b1011111111: data <= 19'h7ffb3; 
        10'b1100000000: data <= 19'h00049; 
        10'b1100000001: data <= 19'h7ffbc; 
        10'b1100000010: data <= 19'h0004f; 
        10'b1100000011: data <= 19'h000ec; 
        10'b1100000100: data <= 19'h00016; 
        10'b1100000101: data <= 19'h00081; 
        10'b1100000110: data <= 19'h001a4; 
        10'b1100000111: data <= 19'h00176; 
        10'b1100001000: data <= 19'h000d3; 
        10'b1100001001: data <= 19'h00081; 
        10'b1100001010: data <= 19'h7ff98; 
        10'b1100001011: data <= 19'h0019f; 
        10'b1100001100: data <= 19'h000e1; 
        10'b1100001101: data <= 19'h7ffb3; 
        10'b1100001110: data <= 19'h0001d; 
        10'b1100001111: data <= 19'h7ffd6; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 14) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 20'h00242; 
        10'b0000000001: data <= 20'h001fb; 
        10'b0000000010: data <= 20'hfff64; 
        10'b0000000011: data <= 20'h00163; 
        10'b0000000100: data <= 20'h00148; 
        10'b0000000101: data <= 20'h00212; 
        10'b0000000110: data <= 20'hfff39; 
        10'b0000000111: data <= 20'h00063; 
        10'b0000001000: data <= 20'h00263; 
        10'b0000001001: data <= 20'hfff06; 
        10'b0000001010: data <= 20'hfffb6; 
        10'b0000001011: data <= 20'h0010b; 
        10'b0000001100: data <= 20'h00303; 
        10'b0000001101: data <= 20'h001f7; 
        10'b0000001110: data <= 20'hffec5; 
        10'b0000001111: data <= 20'hfff6f; 
        10'b0000010000: data <= 20'hfff60; 
        10'b0000010001: data <= 20'h0012f; 
        10'b0000010010: data <= 20'h0022d; 
        10'b0000010011: data <= 20'h00029; 
        10'b0000010100: data <= 20'h00038; 
        10'b0000010101: data <= 20'hfffd8; 
        10'b0000010110: data <= 20'hfff09; 
        10'b0000010111: data <= 20'h00056; 
        10'b0000011000: data <= 20'h00272; 
        10'b0000011001: data <= 20'h000bd; 
        10'b0000011010: data <= 20'hffee2; 
        10'b0000011011: data <= 20'h00136; 
        10'b0000011100: data <= 20'h00206; 
        10'b0000011101: data <= 20'h001b2; 
        10'b0000011110: data <= 20'h000d1; 
        10'b0000011111: data <= 20'hfff87; 
        10'b0000100000: data <= 20'hffed3; 
        10'b0000100001: data <= 20'hfff0a; 
        10'b0000100010: data <= 20'hfffce; 
        10'b0000100011: data <= 20'h00308; 
        10'b0000100100: data <= 20'hffedb; 
        10'b0000100101: data <= 20'h00276; 
        10'b0000100110: data <= 20'h000f3; 
        10'b0000100111: data <= 20'h00184; 
        10'b0000101000: data <= 20'h00130; 
        10'b0000101001: data <= 20'h001b8; 
        10'b0000101010: data <= 20'h0000c; 
        10'b0000101011: data <= 20'hffeab; 
        10'b0000101100: data <= 20'hfff52; 
        10'b0000101101: data <= 20'h001df; 
        10'b0000101110: data <= 20'hfffeb; 
        10'b0000101111: data <= 20'h00088; 
        10'b0000110000: data <= 20'h00260; 
        10'b0000110001: data <= 20'hfffd2; 
        10'b0000110010: data <= 20'h0006a; 
        10'b0000110011: data <= 20'h00037; 
        10'b0000110100: data <= 20'h0014f; 
        10'b0000110101: data <= 20'h0028b; 
        10'b0000110110: data <= 20'hffff8; 
        10'b0000110111: data <= 20'h0008b; 
        10'b0000111000: data <= 20'h002ae; 
        10'b0000111001: data <= 20'h002c0; 
        10'b0000111010: data <= 20'h00035; 
        10'b0000111011: data <= 20'h001df; 
        10'b0000111100: data <= 20'h00245; 
        10'b0000111101: data <= 20'hfffe5; 
        10'b0000111110: data <= 20'hfffbc; 
        10'b0000111111: data <= 20'h000d0; 
        10'b0001000000: data <= 20'h00247; 
        10'b0001000001: data <= 20'hfffac; 
        10'b0001000010: data <= 20'hfff4e; 
        10'b0001000011: data <= 20'h001be; 
        10'b0001000100: data <= 20'h00107; 
        10'b0001000101: data <= 20'h0022d; 
        10'b0001000110: data <= 20'hffeb8; 
        10'b0001000111: data <= 20'h0024c; 
        10'b0001001000: data <= 20'hfff2c; 
        10'b0001001001: data <= 20'hfff1f; 
        10'b0001001010: data <= 20'h00036; 
        10'b0001001011: data <= 20'hffee7; 
        10'b0001001100: data <= 20'h002a3; 
        10'b0001001101: data <= 20'hfff4f; 
        10'b0001001110: data <= 20'hfff0e; 
        10'b0001001111: data <= 20'h002a0; 
        10'b0001010000: data <= 20'h00079; 
        10'b0001010001: data <= 20'h00075; 
        10'b0001010010: data <= 20'h00096; 
        10'b0001010011: data <= 20'h0012b; 
        10'b0001010100: data <= 20'h00345; 
        10'b0001010101: data <= 20'h0001c; 
        10'b0001010110: data <= 20'hfffb3; 
        10'b0001010111: data <= 20'h000f8; 
        10'b0001011000: data <= 20'h00106; 
        10'b0001011001: data <= 20'hffeeb; 
        10'b0001011010: data <= 20'h002ad; 
        10'b0001011011: data <= 20'h00177; 
        10'b0001011100: data <= 20'hfff79; 
        10'b0001011101: data <= 20'h002b4; 
        10'b0001011110: data <= 20'h000d9; 
        10'b0001011111: data <= 20'h00221; 
        10'b0001100000: data <= 20'hfffc8; 
        10'b0001100001: data <= 20'hffd91; 
        10'b0001100010: data <= 20'hfffc8; 
        10'b0001100011: data <= 20'hffc4c; 
        10'b0001100100: data <= 20'hfff8b; 
        10'b0001100101: data <= 20'hffe12; 
        10'b0001100110: data <= 20'h000a4; 
        10'b0001100111: data <= 20'h00063; 
        10'b0001101000: data <= 20'h000d3; 
        10'b0001101001: data <= 20'hfffcb; 
        10'b0001101010: data <= 20'h00220; 
        10'b0001101011: data <= 20'hfffbb; 
        10'b0001101100: data <= 20'hfffb0; 
        10'b0001101101: data <= 20'h002ed; 
        10'b0001101110: data <= 20'h00116; 
        10'b0001101111: data <= 20'h001dc; 
        10'b0001110000: data <= 20'h0005c; 
        10'b0001110001: data <= 20'h0009b; 
        10'b0001110010: data <= 20'h00026; 
        10'b0001110011: data <= 20'hfff5f; 
        10'b0001110100: data <= 20'hffef6; 
        10'b0001110101: data <= 20'h001e2; 
        10'b0001110110: data <= 20'h0014d; 
        10'b0001110111: data <= 20'hfffc3; 
        10'b0001111000: data <= 20'hffe58; 
        10'b0001111001: data <= 20'h000a1; 
        10'b0001111010: data <= 20'hffd43; 
        10'b0001111011: data <= 20'hffc25; 
        10'b0001111100: data <= 20'hffa94; 
        10'b0001111101: data <= 20'hff629; 
        10'b0001111110: data <= 20'hff37a; 
        10'b0001111111: data <= 20'hfef43; 
        10'b0010000000: data <= 20'hff3a1; 
        10'b0010000001: data <= 20'hff398; 
        10'b0010000010: data <= 20'hff6c6; 
        10'b0010000011: data <= 20'hffbf1; 
        10'b0010000100: data <= 20'hffe19; 
        10'b0010000101: data <= 20'hffea2; 
        10'b0010000110: data <= 20'h00075; 
        10'b0010000111: data <= 20'h00255; 
        10'b0010001000: data <= 20'h001d4; 
        10'b0010001001: data <= 20'h001b1; 
        10'b0010001010: data <= 20'h00003; 
        10'b0010001011: data <= 20'h00015; 
        10'b0010001100: data <= 20'h00243; 
        10'b0010001101: data <= 20'h0019b; 
        10'b0010001110: data <= 20'h001e1; 
        10'b0010001111: data <= 20'h00131; 
        10'b0010010000: data <= 20'h00170; 
        10'b0010010001: data <= 20'hffe37; 
        10'b0010010010: data <= 20'hffe6a; 
        10'b0010010011: data <= 20'hffe3d; 
        10'b0010010100: data <= 20'hffa52; 
        10'b0010010101: data <= 20'hffa6f; 
        10'b0010010110: data <= 20'hff9fc; 
        10'b0010010111: data <= 20'hff814; 
        10'b0010011000: data <= 20'hff613; 
        10'b0010011001: data <= 20'hff443; 
        10'b0010011010: data <= 20'hfee15; 
        10'b0010011011: data <= 20'hfeca7; 
        10'b0010011100: data <= 20'hfe78c; 
        10'b0010011101: data <= 20'hfefe1; 
        10'b0010011110: data <= 20'hff5d7; 
        10'b0010011111: data <= 20'hffb14; 
        10'b0010100000: data <= 20'hffacf; 
        10'b0010100001: data <= 20'hff93d; 
        10'b0010100010: data <= 20'hff9b5; 
        10'b0010100011: data <= 20'hffb83; 
        10'b0010100100: data <= 20'hffe36; 
        10'b0010100101: data <= 20'hfff2c; 
        10'b0010100110: data <= 20'h00046; 
        10'b0010100111: data <= 20'h00196; 
        10'b0010101000: data <= 20'h00208; 
        10'b0010101001: data <= 20'h00217; 
        10'b0010101010: data <= 20'hffeb0; 
        10'b0010101011: data <= 20'h0021c; 
        10'b0010101100: data <= 20'h00157; 
        10'b0010101101: data <= 20'hff9f4; 
        10'b0010101110: data <= 20'hff8a4; 
        10'b0010101111: data <= 20'hff755; 
        10'b0010110000: data <= 20'hff63b; 
        10'b0010110001: data <= 20'hff403; 
        10'b0010110010: data <= 20'hff732; 
        10'b0010110011: data <= 20'hffd30; 
        10'b0010110100: data <= 20'h000b5; 
        10'b0010110101: data <= 20'h00ad2; 
        10'b0010110110: data <= 20'h01025; 
        10'b0010110111: data <= 20'h00cd7; 
        10'b0010111000: data <= 20'h008ff; 
        10'b0010111001: data <= 20'h0077a; 
        10'b0010111010: data <= 20'h0097b; 
        10'b0010111011: data <= 20'hffe67; 
        10'b0010111100: data <= 20'hffdb8; 
        10'b0010111101: data <= 20'hff8c9; 
        10'b0010111110: data <= 20'hff312; 
        10'b0010111111: data <= 20'hff3f8; 
        10'b0011000000: data <= 20'hff91c; 
        10'b0011000001: data <= 20'hffca5; 
        10'b0011000010: data <= 20'hfff7e; 
        10'b0011000011: data <= 20'h00118; 
        10'b0011000100: data <= 20'h0031e; 
        10'b0011000101: data <= 20'hfffe3; 
        10'b0011000110: data <= 20'hffefc; 
        10'b0011000111: data <= 20'hffee0; 
        10'b0011001000: data <= 20'hff917; 
        10'b0011001001: data <= 20'hff57e; 
        10'b0011001010: data <= 20'hff3a1; 
        10'b0011001011: data <= 20'hff146; 
        10'b0011001100: data <= 20'hff213; 
        10'b0011001101: data <= 20'hffb17; 
        10'b0011001110: data <= 20'hfff99; 
        10'b0011001111: data <= 20'h003d1; 
        10'b0011010000: data <= 20'h00eaa; 
        10'b0011010001: data <= 20'h01181; 
        10'b0011010010: data <= 20'h01800; 
        10'b0011010011: data <= 20'h01820; 
        10'b0011010100: data <= 20'h01919; 
        10'b0011010101: data <= 20'h00b60; 
        10'b0011010110: data <= 20'h00891; 
        10'b0011010111: data <= 20'h000ed; 
        10'b0011011000: data <= 20'h00239; 
        10'b0011011001: data <= 20'h00285; 
        10'b0011011010: data <= 20'hff75b; 
        10'b0011011011: data <= 20'hff083; 
        10'b0011011100: data <= 20'hff6df; 
        10'b0011011101: data <= 20'hffdb8; 
        10'b0011011110: data <= 20'hffdaa; 
        10'b0011011111: data <= 20'h0020c; 
        10'b0011100000: data <= 20'h00306; 
        10'b0011100001: data <= 20'h0030b; 
        10'b0011100010: data <= 20'h0018c; 
        10'b0011100011: data <= 20'hfff12; 
        10'b0011100100: data <= 20'hff8cf; 
        10'b0011100101: data <= 20'hff51d; 
        10'b0011100110: data <= 20'hff353; 
        10'b0011100111: data <= 20'hfee47; 
        10'b0011101000: data <= 20'hffb51; 
        10'b0011101001: data <= 20'hffdd5; 
        10'b0011101010: data <= 20'hffd7d; 
        10'b0011101011: data <= 20'hffaf5; 
        10'b0011101100: data <= 20'hfff9d; 
        10'b0011101101: data <= 20'h00706; 
        10'b0011101110: data <= 20'h01491; 
        10'b0011101111: data <= 20'h00b5a; 
        10'b0011110000: data <= 20'h00b8f; 
        10'b0011110001: data <= 20'h0025e; 
        10'b0011110010: data <= 20'h000e9; 
        10'b0011110011: data <= 20'h0009d; 
        10'b0011110100: data <= 20'hffc33; 
        10'b0011110101: data <= 20'h001f9; 
        10'b0011110110: data <= 20'hffb21; 
        10'b0011110111: data <= 20'hff3a5; 
        10'b0011111000: data <= 20'hff590; 
        10'b0011111001: data <= 20'hffaff; 
        10'b0011111010: data <= 20'hffdd0; 
        10'b0011111011: data <= 20'h002d2; 
        10'b0011111100: data <= 20'h000eb; 
        10'b0011111101: data <= 20'h0008d; 
        10'b0011111110: data <= 20'h00035; 
        10'b0011111111: data <= 20'hffadb; 
        10'b0100000000: data <= 20'hff4c8; 
        10'b0100000001: data <= 20'hff766; 
        10'b0100000010: data <= 20'hffd90; 
        10'b0100000011: data <= 20'hffb12; 
        10'b0100000100: data <= 20'hffd11; 
        10'b0100000101: data <= 20'hffeab; 
        10'b0100000110: data <= 20'h00546; 
        10'b0100000111: data <= 20'h0032d; 
        10'b0100001000: data <= 20'h000ee; 
        10'b0100001001: data <= 20'h0087f; 
        10'b0100001010: data <= 20'h00e3a; 
        10'b0100001011: data <= 20'h00caf; 
        10'b0100001100: data <= 20'hfff82; 
        10'b0100001101: data <= 20'hffc5d; 
        10'b0100001110: data <= 20'h00024; 
        10'b0100001111: data <= 20'hff86d; 
        10'b0100010000: data <= 20'hffcca; 
        10'b0100010001: data <= 20'hff810; 
        10'b0100010010: data <= 20'hff780; 
        10'b0100010011: data <= 20'hff6ee; 
        10'b0100010100: data <= 20'hff9d1; 
        10'b0100010101: data <= 20'hffd4c; 
        10'b0100010110: data <= 20'hffe0a; 
        10'b0100010111: data <= 20'h00281; 
        10'b0100011000: data <= 20'h0008b; 
        10'b0100011001: data <= 20'hfffe4; 
        10'b0100011010: data <= 20'hffecb; 
        10'b0100011011: data <= 20'hffe08; 
        10'b0100011100: data <= 20'hff75c; 
        10'b0100011101: data <= 20'hffb7b; 
        10'b0100011110: data <= 20'h00437; 
        10'b0100011111: data <= 20'h00585; 
        10'b0100100000: data <= 20'h00b34; 
        10'b0100100001: data <= 20'h00b1f; 
        10'b0100100010: data <= 20'h00994; 
        10'b0100100011: data <= 20'h00e6c; 
        10'b0100100100: data <= 20'h00743; 
        10'b0100100101: data <= 20'h001b6; 
        10'b0100100110: data <= 20'h001db; 
        10'b0100100111: data <= 20'hff8b3; 
        10'b0100101000: data <= 20'hffba6; 
        10'b0100101001: data <= 20'hfff24; 
        10'b0100101010: data <= 20'h00516; 
        10'b0100101011: data <= 20'hfffe4; 
        10'b0100101100: data <= 20'h00417; 
        10'b0100101101: data <= 20'hffd8f; 
        10'b0100101110: data <= 20'hffafb; 
        10'b0100101111: data <= 20'hffb43; 
        10'b0100110000: data <= 20'hff9fc; 
        10'b0100110001: data <= 20'hffe48; 
        10'b0100110010: data <= 20'hffdba; 
        10'b0100110011: data <= 20'h00170; 
        10'b0100110100: data <= 20'hfff87; 
        10'b0100110101: data <= 20'h00093; 
        10'b0100110110: data <= 20'hffeb3; 
        10'b0100110111: data <= 20'hfff2d; 
        10'b0100111000: data <= 20'hffda1; 
        10'b0100111001: data <= 20'h007f3; 
        10'b0100111010: data <= 20'h01265; 
        10'b0100111011: data <= 20'h00dba; 
        10'b0100111100: data <= 20'h01592; 
        10'b0100111101: data <= 20'h008a6; 
        10'b0100111110: data <= 20'h008f7; 
        10'b0100111111: data <= 20'h00f67; 
        10'b0101000000: data <= 20'hffb1a; 
        10'b0101000001: data <= 20'hffbd6; 
        10'b0101000010: data <= 20'hffdc0; 
        10'b0101000011: data <= 20'h00116; 
        10'b0101000100: data <= 20'h005f4; 
        10'b0101000101: data <= 20'h014d8; 
        10'b0101000110: data <= 20'h009d9; 
        10'b0101000111: data <= 20'h009fb; 
        10'b0101001000: data <= 20'h0105e; 
        10'b0101001001: data <= 20'h00bd8; 
        10'b0101001010: data <= 20'h006ec; 
        10'b0101001011: data <= 20'h0016e; 
        10'b0101001100: data <= 20'hffede; 
        10'b0101001101: data <= 20'hffd2e; 
        10'b0101001110: data <= 20'hfffe1; 
        10'b0101001111: data <= 20'h00003; 
        10'b0101010000: data <= 20'h0014d; 
        10'b0101010001: data <= 20'h002af; 
        10'b0101010010: data <= 20'hffe26; 
        10'b0101010011: data <= 20'hffd0c; 
        10'b0101010100: data <= 20'h006b6; 
        10'b0101010101: data <= 20'h01171; 
        10'b0101010110: data <= 20'h0142d; 
        10'b0101010111: data <= 20'h00bf8; 
        10'b0101011000: data <= 20'h00ef6; 
        10'b0101011001: data <= 20'h0124b; 
        10'b0101011010: data <= 20'h00bae; 
        10'b0101011011: data <= 20'h00023; 
        10'b0101011100: data <= 20'hff448; 
        10'b0101011101: data <= 20'h00a27; 
        10'b0101011110: data <= 20'h015ef; 
        10'b0101011111: data <= 20'h0115a; 
        10'b0101100000: data <= 20'h00ed6; 
        10'b0101100001: data <= 20'h016af; 
        10'b0101100010: data <= 20'h016d9; 
        10'b0101100011: data <= 20'h017b6; 
        10'b0101100100: data <= 20'h01860; 
        10'b0101100101: data <= 20'h0104a; 
        10'b0101100110: data <= 20'h007d5; 
        10'b0101100111: data <= 20'h00035; 
        10'b0101101000: data <= 20'hffc5f; 
        10'b0101101001: data <= 20'h00098; 
        10'b0101101010: data <= 20'h00151; 
        10'b0101101011: data <= 20'h0016d; 
        10'b0101101100: data <= 20'h00304; 
        10'b0101101101: data <= 20'h001da; 
        10'b0101101110: data <= 20'hffd76; 
        10'b0101101111: data <= 20'h000f4; 
        10'b0101110000: data <= 20'h00a26; 
        10'b0101110001: data <= 20'h00f43; 
        10'b0101110010: data <= 20'h00e62; 
        10'b0101110011: data <= 20'h00971; 
        10'b0101110100: data <= 20'h00bda; 
        10'b0101110101: data <= 20'h0079c; 
        10'b0101110110: data <= 20'h006e0; 
        10'b0101110111: data <= 20'hffc70; 
        10'b0101111000: data <= 20'hff9d9; 
        10'b0101111001: data <= 20'h00ff5; 
        10'b0101111010: data <= 20'h015e3; 
        10'b0101111011: data <= 20'h00fdc; 
        10'b0101111100: data <= 20'h01247; 
        10'b0101111101: data <= 20'h01063; 
        10'b0101111110: data <= 20'h0167a; 
        10'b0101111111: data <= 20'h016de; 
        10'b0110000000: data <= 20'h011e0; 
        10'b0110000001: data <= 20'h00a71; 
        10'b0110000010: data <= 20'h00099; 
        10'b0110000011: data <= 20'hff8e4; 
        10'b0110000100: data <= 20'hffbdb; 
        10'b0110000101: data <= 20'hffeb7; 
        10'b0110000110: data <= 20'h00159; 
        10'b0110000111: data <= 20'h0015f; 
        10'b0110001000: data <= 20'h0009b; 
        10'b0110001001: data <= 20'h0004d; 
        10'b0110001010: data <= 20'h00213; 
        10'b0110001011: data <= 20'h00151; 
        10'b0110001100: data <= 20'h004a5; 
        10'b0110001101: data <= 20'h00460; 
        10'b0110001110: data <= 20'h00bea; 
        10'b0110001111: data <= 20'h00856; 
        10'b0110010000: data <= 20'h0040d; 
        10'b0110010001: data <= 20'hffff5; 
        10'b0110010010: data <= 20'h0017c; 
        10'b0110010011: data <= 20'hfff43; 
        10'b0110010100: data <= 20'hffb81; 
        10'b0110010101: data <= 20'h0052d; 
        10'b0110010110: data <= 20'h002f0; 
        10'b0110010111: data <= 20'h00dff; 
        10'b0110011000: data <= 20'h00ed8; 
        10'b0110011001: data <= 20'h00edd; 
        10'b0110011010: data <= 20'h00a20; 
        10'b0110011011: data <= 20'h00682; 
        10'b0110011100: data <= 20'h0081e; 
        10'b0110011101: data <= 20'h00026; 
        10'b0110011110: data <= 20'hff7ce; 
        10'b0110011111: data <= 20'hff417; 
        10'b0110100000: data <= 20'hffb13; 
        10'b0110100001: data <= 20'h000d2; 
        10'b0110100010: data <= 20'h00078; 
        10'b0110100011: data <= 20'h0008e; 
        10'b0110100100: data <= 20'h00248; 
        10'b0110100101: data <= 20'h00215; 
        10'b0110100110: data <= 20'h00161; 
        10'b0110100111: data <= 20'hffe56; 
        10'b0110101000: data <= 20'h00057; 
        10'b0110101001: data <= 20'h0054d; 
        10'b0110101010: data <= 20'h00513; 
        10'b0110101011: data <= 20'h0035a; 
        10'b0110101100: data <= 20'h0036b; 
        10'b0110101101: data <= 20'hff9b8; 
        10'b0110101110: data <= 20'hffd15; 
        10'b0110101111: data <= 20'hffd10; 
        10'b0110110000: data <= 20'hffb9d; 
        10'b0110110001: data <= 20'hffc9b; 
        10'b0110110010: data <= 20'hffbe3; 
        10'b0110110011: data <= 20'h00f4a; 
        10'b0110110100: data <= 20'h01662; 
        10'b0110110101: data <= 20'h01575; 
        10'b0110110110: data <= 20'h00abe; 
        10'b0110110111: data <= 20'h00109; 
        10'b0110111000: data <= 20'hffb55; 
        10'b0110111001: data <= 20'hff3b2; 
        10'b0110111010: data <= 20'hff0a7; 
        10'b0110111011: data <= 20'hff50a; 
        10'b0110111100: data <= 20'hffb1f; 
        10'b0110111101: data <= 20'h00017; 
        10'b0110111110: data <= 20'h00141; 
        10'b0110111111: data <= 20'hfffd2; 
        10'b0111000000: data <= 20'h002a1; 
        10'b0111000001: data <= 20'h00038; 
        10'b0111000010: data <= 20'hffe1e; 
        10'b0111000011: data <= 20'hfff84; 
        10'b0111000100: data <= 20'h0002b; 
        10'b0111000101: data <= 20'h00197; 
        10'b0111000110: data <= 20'hffbe6; 
        10'b0111000111: data <= 20'h0033d; 
        10'b0111001000: data <= 20'h00934; 
        10'b0111001001: data <= 20'hffdd8; 
        10'b0111001010: data <= 20'h00538; 
        10'b0111001011: data <= 20'h00767; 
        10'b0111001100: data <= 20'hffefe; 
        10'b0111001101: data <= 20'hff794; 
        10'b0111001110: data <= 20'hffe97; 
        10'b0111001111: data <= 20'h0087d; 
        10'b0111010000: data <= 20'h00f46; 
        10'b0111010001: data <= 20'h00f2d; 
        10'b0111010010: data <= 20'h003ca; 
        10'b0111010011: data <= 20'hff75f; 
        10'b0111010100: data <= 20'hff1ae; 
        10'b0111010101: data <= 20'hfec33; 
        10'b0111010110: data <= 20'hff219; 
        10'b0111010111: data <= 20'hff4b4; 
        10'b0111011000: data <= 20'hff886; 
        10'b0111011001: data <= 20'h0003f; 
        10'b0111011010: data <= 20'hffe5e; 
        10'b0111011011: data <= 20'h0016a; 
        10'b0111011100: data <= 20'h000de; 
        10'b0111011101: data <= 20'hfff6c; 
        10'b0111011110: data <= 20'hffdf2; 
        10'b0111011111: data <= 20'hffcff; 
        10'b0111100000: data <= 20'hffa5f; 
        10'b0111100001: data <= 20'hff927; 
        10'b0111100010: data <= 20'hffa5b; 
        10'b0111100011: data <= 20'h0028b; 
        10'b0111100100: data <= 20'h004f5; 
        10'b0111100101: data <= 20'h005a5; 
        10'b0111100110: data <= 20'h0089b; 
        10'b0111100111: data <= 20'h00c86; 
        10'b0111101000: data <= 20'h007a3; 
        10'b0111101001: data <= 20'h0038d; 
        10'b0111101010: data <= 20'h004da; 
        10'b0111101011: data <= 20'h00c75; 
        10'b0111101100: data <= 20'h003b3; 
        10'b0111101101: data <= 20'hffd7a; 
        10'b0111101110: data <= 20'hffa7f; 
        10'b0111101111: data <= 20'hff35a; 
        10'b0111110000: data <= 20'hff383; 
        10'b0111110001: data <= 20'hff28f; 
        10'b0111110010: data <= 20'hff35c; 
        10'b0111110011: data <= 20'hff6b2; 
        10'b0111110100: data <= 20'hff939; 
        10'b0111110101: data <= 20'h000ad; 
        10'b0111110110: data <= 20'h000b3; 
        10'b0111110111: data <= 20'hfff67; 
        10'b0111111000: data <= 20'h0026d; 
        10'b0111111001: data <= 20'hffffe; 
        10'b0111111010: data <= 20'hffe96; 
        10'b0111111011: data <= 20'hfff70; 
        10'b0111111100: data <= 20'hffb0d; 
        10'b0111111101: data <= 20'hff4a4; 
        10'b0111111110: data <= 20'hff46b; 
        10'b0111111111: data <= 20'hff4a4; 
        10'b1000000000: data <= 20'hffb3a; 
        10'b1000000001: data <= 20'h001e5; 
        10'b1000000010: data <= 20'h00db9; 
        10'b1000000011: data <= 20'h00b17; 
        10'b1000000100: data <= 20'hff93b; 
        10'b1000000101: data <= 20'hff921; 
        10'b1000000110: data <= 20'h0006d; 
        10'b1000000111: data <= 20'h0083f; 
        10'b1000001000: data <= 20'hffaf2; 
        10'b1000001001: data <= 20'hffa3c; 
        10'b1000001010: data <= 20'hff534; 
        10'b1000001011: data <= 20'hff981; 
        10'b1000001100: data <= 20'hff9e8; 
        10'b1000001101: data <= 20'hff67e; 
        10'b1000001110: data <= 20'hff5fe; 
        10'b1000001111: data <= 20'hff586; 
        10'b1000010000: data <= 20'hff897; 
        10'b1000010001: data <= 20'hffed2; 
        10'b1000010010: data <= 20'h00026; 
        10'b1000010011: data <= 20'h00238; 
        10'b1000010100: data <= 20'h00193; 
        10'b1000010101: data <= 20'h00325; 
        10'b1000010110: data <= 20'h0008f; 
        10'b1000010111: data <= 20'hffd48; 
        10'b1000011000: data <= 20'hffb75; 
        10'b1000011001: data <= 20'hff7f6; 
        10'b1000011010: data <= 20'hff34b; 
        10'b1000011011: data <= 20'hff2f5; 
        10'b1000011100: data <= 20'hff27f; 
        10'b1000011101: data <= 20'hff29b; 
        10'b1000011110: data <= 20'hff102; 
        10'b1000011111: data <= 20'hff356; 
        10'b1000100000: data <= 20'hfef9c; 
        10'b1000100001: data <= 20'hff48b; 
        10'b1000100010: data <= 20'hff658; 
        10'b1000100011: data <= 20'hff504; 
        10'b1000100100: data <= 20'hff685; 
        10'b1000100101: data <= 20'hffce7; 
        10'b1000100110: data <= 20'hff8c9; 
        10'b1000100111: data <= 20'hffdfc; 
        10'b1000101000: data <= 20'hffb2d; 
        10'b1000101001: data <= 20'hffa48; 
        10'b1000101010: data <= 20'hffa9a; 
        10'b1000101011: data <= 20'hffb33; 
        10'b1000101100: data <= 20'hffcfb; 
        10'b1000101101: data <= 20'h000de; 
        10'b1000101110: data <= 20'hfff0d; 
        10'b1000101111: data <= 20'h00056; 
        10'b1000110000: data <= 20'hfff69; 
        10'b1000110001: data <= 20'h00070; 
        10'b1000110010: data <= 20'h00156; 
        10'b1000110011: data <= 20'h0001a; 
        10'b1000110100: data <= 20'hffb4c; 
        10'b1000110101: data <= 20'hff83c; 
        10'b1000110110: data <= 20'hff43a; 
        10'b1000110111: data <= 20'hfed8f; 
        10'b1000111000: data <= 20'hfeae1; 
        10'b1000111001: data <= 20'hfe84f; 
        10'b1000111010: data <= 20'hfdfed; 
        10'b1000111011: data <= 20'hfe774; 
        10'b1000111100: data <= 20'hfe815; 
        10'b1000111101: data <= 20'hff82c; 
        10'b1000111110: data <= 20'hff506; 
        10'b1000111111: data <= 20'hffad8; 
        10'b1001000000: data <= 20'hff9d1; 
        10'b1001000001: data <= 20'hffe55; 
        10'b1001000010: data <= 20'hff57d; 
        10'b1001000011: data <= 20'hffc8a; 
        10'b1001000100: data <= 20'hffbd4; 
        10'b1001000101: data <= 20'hff94d; 
        10'b1001000110: data <= 20'hffe1d; 
        10'b1001000111: data <= 20'hffcca; 
        10'b1001001000: data <= 20'h00053; 
        10'b1001001001: data <= 20'h002ad; 
        10'b1001001010: data <= 20'h0019d; 
        10'b1001001011: data <= 20'h00082; 
        10'b1001001100: data <= 20'h00037; 
        10'b1001001101: data <= 20'h00001; 
        10'b1001001110: data <= 20'h002ad; 
        10'b1001001111: data <= 20'hffd2a; 
        10'b1001010000: data <= 20'hffcd6; 
        10'b1001010001: data <= 20'hff858; 
        10'b1001010010: data <= 20'hff530; 
        10'b1001010011: data <= 20'hfef50; 
        10'b1001010100: data <= 20'hfed0f; 
        10'b1001010101: data <= 20'hfeb29; 
        10'b1001010110: data <= 20'hfea28; 
        10'b1001010111: data <= 20'hfec5b; 
        10'b1001011000: data <= 20'hff37c; 
        10'b1001011001: data <= 20'hff3a6; 
        10'b1001011010: data <= 20'hff371; 
        10'b1001011011: data <= 20'hff8cb; 
        10'b1001011100: data <= 20'hff832; 
        10'b1001011101: data <= 20'hff440; 
        10'b1001011110: data <= 20'hff1d3; 
        10'b1001011111: data <= 20'hff9fe; 
        10'b1001100000: data <= 20'hffca6; 
        10'b1001100001: data <= 20'hffe11; 
        10'b1001100010: data <= 20'h000f2; 
        10'b1001100011: data <= 20'hfffbb; 
        10'b1001100100: data <= 20'h00134; 
        10'b1001100101: data <= 20'h001a5; 
        10'b1001100110: data <= 20'h00018; 
        10'b1001100111: data <= 20'h00032; 
        10'b1001101000: data <= 20'h0020e; 
        10'b1001101001: data <= 20'h00083; 
        10'b1001101010: data <= 20'h00094; 
        10'b1001101011: data <= 20'h001f7; 
        10'b1001101100: data <= 20'hffebd; 
        10'b1001101101: data <= 20'hff9d1; 
        10'b1001101110: data <= 20'hff61b; 
        10'b1001101111: data <= 20'hff28b; 
        10'b1001110000: data <= 20'hff5fc; 
        10'b1001110001: data <= 20'hff589; 
        10'b1001110010: data <= 20'hff493; 
        10'b1001110011: data <= 20'hff849; 
        10'b1001110100: data <= 20'hff754; 
        10'b1001110101: data <= 20'hff476; 
        10'b1001110110: data <= 20'hff64d; 
        10'b1001110111: data <= 20'hff268; 
        10'b1001111000: data <= 20'hff0f7; 
        10'b1001111001: data <= 20'hff142; 
        10'b1001111010: data <= 20'hff3be; 
        10'b1001111011: data <= 20'hff51a; 
        10'b1001111100: data <= 20'hffd02; 
        10'b1001111101: data <= 20'h003ab; 
        10'b1001111110: data <= 20'h0020a; 
        10'b1001111111: data <= 20'h00288; 
        10'b1010000000: data <= 20'h00423; 
        10'b1010000001: data <= 20'h000de; 
        10'b1010000010: data <= 20'h000f7; 
        10'b1010000011: data <= 20'h00182; 
        10'b1010000100: data <= 20'h00269; 
        10'b1010000101: data <= 20'h001e4; 
        10'b1010000110: data <= 20'h000b5; 
        10'b1010000111: data <= 20'hfff0e; 
        10'b1010001000: data <= 20'hffe44; 
        10'b1010001001: data <= 20'hffaaf; 
        10'b1010001010: data <= 20'hff9d1; 
        10'b1010001011: data <= 20'hff7d3; 
        10'b1010001100: data <= 20'hfff62; 
        10'b1010001101: data <= 20'hffcb2; 
        10'b1010001110: data <= 20'hffd5a; 
        10'b1010001111: data <= 20'hff618; 
        10'b1010010000: data <= 20'hff7ed; 
        10'b1010010001: data <= 20'hff5d0; 
        10'b1010010010: data <= 20'hff763; 
        10'b1010010011: data <= 20'hff14c; 
        10'b1010010100: data <= 20'hff021; 
        10'b1010010101: data <= 20'hff208; 
        10'b1010010110: data <= 20'hff74c; 
        10'b1010010111: data <= 20'hfff27; 
        10'b1010011000: data <= 20'h00368; 
        10'b1010011001: data <= 20'h007e9; 
        10'b1010011010: data <= 20'h00b67; 
        10'b1010011011: data <= 20'h0098c; 
        10'b1010011100: data <= 20'h00478; 
        10'b1010011101: data <= 20'hfffb2; 
        10'b1010011110: data <= 20'h00334; 
        10'b1010011111: data <= 20'hfffa0; 
        10'b1010100000: data <= 20'hffffd; 
        10'b1010100001: data <= 20'hffebd; 
        10'b1010100010: data <= 20'hfffa9; 
        10'b1010100011: data <= 20'h002b3; 
        10'b1010100100: data <= 20'h001f1; 
        10'b1010100101: data <= 20'h0030a; 
        10'b1010100110: data <= 20'h00236; 
        10'b1010100111: data <= 20'h00335; 
        10'b1010101000: data <= 20'h00489; 
        10'b1010101001: data <= 20'h00272; 
        10'b1010101010: data <= 20'hffe63; 
        10'b1010101011: data <= 20'hffaeb; 
        10'b1010101100: data <= 20'hfffa4; 
        10'b1010101101: data <= 20'hff834; 
        10'b1010101110: data <= 20'hff625; 
        10'b1010101111: data <= 20'hff598; 
        10'b1010110000: data <= 20'hffb48; 
        10'b1010110001: data <= 20'h0036c; 
        10'b1010110010: data <= 20'h005d8; 
        10'b1010110011: data <= 20'h0060a; 
        10'b1010110100: data <= 20'h00dcb; 
        10'b1010110101: data <= 20'h00ed8; 
        10'b1010110110: data <= 20'h0088b; 
        10'b1010110111: data <= 20'h00539; 
        10'b1010111000: data <= 20'h0041f; 
        10'b1010111001: data <= 20'hfff31; 
        10'b1010111010: data <= 20'h001d8; 
        10'b1010111011: data <= 20'hfffe1; 
        10'b1010111100: data <= 20'h000ac; 
        10'b1010111101: data <= 20'h002ad; 
        10'b1010111110: data <= 20'h002af; 
        10'b1010111111: data <= 20'hfffb8; 
        10'b1011000000: data <= 20'h00040; 
        10'b1011000001: data <= 20'h00495; 
        10'b1011000010: data <= 20'h00379; 
        10'b1011000011: data <= 20'h00a05; 
        10'b1011000100: data <= 20'h00afb; 
        10'b1011000101: data <= 20'h00b2e; 
        10'b1011000110: data <= 20'h009ac; 
        10'b1011000111: data <= 20'h003d7; 
        10'b1011001000: data <= 20'h00a2d; 
        10'b1011001001: data <= 20'h00913; 
        10'b1011001010: data <= 20'h008b1; 
        10'b1011001011: data <= 20'h0082b; 
        10'b1011001100: data <= 20'h00f42; 
        10'b1011001101: data <= 20'h01095; 
        10'b1011001110: data <= 20'h0123d; 
        10'b1011001111: data <= 20'h01309; 
        10'b1011010000: data <= 20'h01540; 
        10'b1011010001: data <= 20'h00f14; 
        10'b1011010010: data <= 20'h005e2; 
        10'b1011010011: data <= 20'h002ca; 
        10'b1011010100: data <= 20'hfffa0; 
        10'b1011010101: data <= 20'hfffc7; 
        10'b1011010110: data <= 20'h000c8; 
        10'b1011010111: data <= 20'h000a8; 
        10'b1011011000: data <= 20'h0001d; 
        10'b1011011001: data <= 20'h00270; 
        10'b1011011010: data <= 20'h000a7; 
        10'b1011011011: data <= 20'hfff1d; 
        10'b1011011100: data <= 20'h00274; 
        10'b1011011101: data <= 20'h003cd; 
        10'b1011011110: data <= 20'h00555; 
        10'b1011011111: data <= 20'h00768; 
        10'b1011100000: data <= 20'h0086e; 
        10'b1011100001: data <= 20'h00cc9; 
        10'b1011100010: data <= 20'h00d31; 
        10'b1011100011: data <= 20'h00ed1; 
        10'b1011100100: data <= 20'h0118c; 
        10'b1011100101: data <= 20'h011b4; 
        10'b1011100110: data <= 20'h015ad; 
        10'b1011100111: data <= 20'h00c81; 
        10'b1011101000: data <= 20'h00890; 
        10'b1011101001: data <= 20'h0073b; 
        10'b1011101010: data <= 20'h00aab; 
        10'b1011101011: data <= 20'h00b83; 
        10'b1011101100: data <= 20'h0085c; 
        10'b1011101101: data <= 20'h005d2; 
        10'b1011101110: data <= 20'h0026c; 
        10'b1011101111: data <= 20'h000e0; 
        10'b1011110000: data <= 20'h0008b; 
        10'b1011110001: data <= 20'h000f7; 
        10'b1011110010: data <= 20'hfff16; 
        10'b1011110011: data <= 20'h00089; 
        10'b1011110100: data <= 20'hfff6a; 
        10'b1011110101: data <= 20'h0011d; 
        10'b1011110110: data <= 20'hffeff; 
        10'b1011110111: data <= 20'h002f4; 
        10'b1011111000: data <= 20'h001b2; 
        10'b1011111001: data <= 20'h000f0; 
        10'b1011111010: data <= 20'hfff95; 
        10'b1011111011: data <= 20'h002df; 
        10'b1011111100: data <= 20'h0026e; 
        10'b1011111101: data <= 20'h001a9; 
        10'b1011111110: data <= 20'hfff77; 
        10'b1011111111: data <= 20'hfff67; 
        10'b1100000000: data <= 20'h00092; 
        10'b1100000001: data <= 20'hfff77; 
        10'b1100000010: data <= 20'h0009f; 
        10'b1100000011: data <= 20'h001d8; 
        10'b1100000100: data <= 20'h0002c; 
        10'b1100000101: data <= 20'h00102; 
        10'b1100000110: data <= 20'h00347; 
        10'b1100000111: data <= 20'h002ec; 
        10'b1100001000: data <= 20'h001a5; 
        10'b1100001001: data <= 20'h00101; 
        10'b1100001010: data <= 20'hfff30; 
        10'b1100001011: data <= 20'h0033e; 
        10'b1100001100: data <= 20'h001c3; 
        10'b1100001101: data <= 20'hfff67; 
        10'b1100001110: data <= 20'h00039; 
        10'b1100001111: data <= 20'hfffac; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 15) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 21'h000485; 
        10'b0000000001: data <= 21'h0003f6; 
        10'b0000000010: data <= 21'h1ffec8; 
        10'b0000000011: data <= 21'h0002c6; 
        10'b0000000100: data <= 21'h00028f; 
        10'b0000000101: data <= 21'h000424; 
        10'b0000000110: data <= 21'h1ffe73; 
        10'b0000000111: data <= 21'h0000c5; 
        10'b0000001000: data <= 21'h0004c6; 
        10'b0000001001: data <= 21'h1ffe0d; 
        10'b0000001010: data <= 21'h1fff6c; 
        10'b0000001011: data <= 21'h000216; 
        10'b0000001100: data <= 21'h000607; 
        10'b0000001101: data <= 21'h0003ed; 
        10'b0000001110: data <= 21'h1ffd8a; 
        10'b0000001111: data <= 21'h1ffedd; 
        10'b0000010000: data <= 21'h1ffec0; 
        10'b0000010001: data <= 21'h00025f; 
        10'b0000010010: data <= 21'h00045b; 
        10'b0000010011: data <= 21'h000052; 
        10'b0000010100: data <= 21'h00006f; 
        10'b0000010101: data <= 21'h1fffaf; 
        10'b0000010110: data <= 21'h1ffe12; 
        10'b0000010111: data <= 21'h0000ad; 
        10'b0000011000: data <= 21'h0004e4; 
        10'b0000011001: data <= 21'h00017a; 
        10'b0000011010: data <= 21'h1ffdc5; 
        10'b0000011011: data <= 21'h00026d; 
        10'b0000011100: data <= 21'h00040d; 
        10'b0000011101: data <= 21'h000363; 
        10'b0000011110: data <= 21'h0001a2; 
        10'b0000011111: data <= 21'h1fff0e; 
        10'b0000100000: data <= 21'h1ffda6; 
        10'b0000100001: data <= 21'h1ffe15; 
        10'b0000100010: data <= 21'h1fff9c; 
        10'b0000100011: data <= 21'h000610; 
        10'b0000100100: data <= 21'h1ffdb7; 
        10'b0000100101: data <= 21'h0004eb; 
        10'b0000100110: data <= 21'h0001e5; 
        10'b0000100111: data <= 21'h000309; 
        10'b0000101000: data <= 21'h000260; 
        10'b0000101001: data <= 21'h000371; 
        10'b0000101010: data <= 21'h000018; 
        10'b0000101011: data <= 21'h1ffd55; 
        10'b0000101100: data <= 21'h1ffea3; 
        10'b0000101101: data <= 21'h0003be; 
        10'b0000101110: data <= 21'h1fffd6; 
        10'b0000101111: data <= 21'h000110; 
        10'b0000110000: data <= 21'h0004bf; 
        10'b0000110001: data <= 21'h1fffa4; 
        10'b0000110010: data <= 21'h0000d5; 
        10'b0000110011: data <= 21'h00006e; 
        10'b0000110100: data <= 21'h00029e; 
        10'b0000110101: data <= 21'h000516; 
        10'b0000110110: data <= 21'h1ffff0; 
        10'b0000110111: data <= 21'h000116; 
        10'b0000111000: data <= 21'h00055b; 
        10'b0000111001: data <= 21'h00057f; 
        10'b0000111010: data <= 21'h00006a; 
        10'b0000111011: data <= 21'h0003be; 
        10'b0000111100: data <= 21'h00048a; 
        10'b0000111101: data <= 21'h1fffca; 
        10'b0000111110: data <= 21'h1fff77; 
        10'b0000111111: data <= 21'h0001a1; 
        10'b0001000000: data <= 21'h00048e; 
        10'b0001000001: data <= 21'h1fff58; 
        10'b0001000010: data <= 21'h1ffe9c; 
        10'b0001000011: data <= 21'h00037c; 
        10'b0001000100: data <= 21'h00020e; 
        10'b0001000101: data <= 21'h00045a; 
        10'b0001000110: data <= 21'h1ffd6f; 
        10'b0001000111: data <= 21'h000498; 
        10'b0001001000: data <= 21'h1ffe59; 
        10'b0001001001: data <= 21'h1ffe3e; 
        10'b0001001010: data <= 21'h00006b; 
        10'b0001001011: data <= 21'h1ffdcf; 
        10'b0001001100: data <= 21'h000546; 
        10'b0001001101: data <= 21'h1ffe9e; 
        10'b0001001110: data <= 21'h1ffe1c; 
        10'b0001001111: data <= 21'h00053f; 
        10'b0001010000: data <= 21'h0000f2; 
        10'b0001010001: data <= 21'h0000ea; 
        10'b0001010010: data <= 21'h00012c; 
        10'b0001010011: data <= 21'h000256; 
        10'b0001010100: data <= 21'h00068a; 
        10'b0001010101: data <= 21'h000039; 
        10'b0001010110: data <= 21'h1fff67; 
        10'b0001010111: data <= 21'h0001ef; 
        10'b0001011000: data <= 21'h00020d; 
        10'b0001011001: data <= 21'h1ffdd6; 
        10'b0001011010: data <= 21'h00055b; 
        10'b0001011011: data <= 21'h0002ee; 
        10'b0001011100: data <= 21'h1ffef2; 
        10'b0001011101: data <= 21'h000568; 
        10'b0001011110: data <= 21'h0001b2; 
        10'b0001011111: data <= 21'h000443; 
        10'b0001100000: data <= 21'h1fff90; 
        10'b0001100001: data <= 21'h1ffb21; 
        10'b0001100010: data <= 21'h1fff90; 
        10'b0001100011: data <= 21'h1ff899; 
        10'b0001100100: data <= 21'h1fff17; 
        10'b0001100101: data <= 21'h1ffc24; 
        10'b0001100110: data <= 21'h000148; 
        10'b0001100111: data <= 21'h0000c6; 
        10'b0001101000: data <= 21'h0001a7; 
        10'b0001101001: data <= 21'h1fff96; 
        10'b0001101010: data <= 21'h00043f; 
        10'b0001101011: data <= 21'h1fff75; 
        10'b0001101100: data <= 21'h1fff5f; 
        10'b0001101101: data <= 21'h0005d9; 
        10'b0001101110: data <= 21'h00022d; 
        10'b0001101111: data <= 21'h0003b7; 
        10'b0001110000: data <= 21'h0000b7; 
        10'b0001110001: data <= 21'h000135; 
        10'b0001110010: data <= 21'h00004c; 
        10'b0001110011: data <= 21'h1ffebd; 
        10'b0001110100: data <= 21'h1ffdec; 
        10'b0001110101: data <= 21'h0003c5; 
        10'b0001110110: data <= 21'h00029b; 
        10'b0001110111: data <= 21'h1fff85; 
        10'b0001111000: data <= 21'h1ffcaf; 
        10'b0001111001: data <= 21'h000143; 
        10'b0001111010: data <= 21'h1ffa85; 
        10'b0001111011: data <= 21'h1ff849; 
        10'b0001111100: data <= 21'h1ff528; 
        10'b0001111101: data <= 21'h1fec53; 
        10'b0001111110: data <= 21'h1fe6f4; 
        10'b0001111111: data <= 21'h1fde85; 
        10'b0010000000: data <= 21'h1fe742; 
        10'b0010000001: data <= 21'h1fe72f; 
        10'b0010000010: data <= 21'h1fed8b; 
        10'b0010000011: data <= 21'h1ff7e3; 
        10'b0010000100: data <= 21'h1ffc33; 
        10'b0010000101: data <= 21'h1ffd44; 
        10'b0010000110: data <= 21'h0000e9; 
        10'b0010000111: data <= 21'h0004aa; 
        10'b0010001000: data <= 21'h0003a7; 
        10'b0010001001: data <= 21'h000363; 
        10'b0010001010: data <= 21'h000006; 
        10'b0010001011: data <= 21'h00002a; 
        10'b0010001100: data <= 21'h000486; 
        10'b0010001101: data <= 21'h000336; 
        10'b0010001110: data <= 21'h0003c1; 
        10'b0010001111: data <= 21'h000261; 
        10'b0010010000: data <= 21'h0002df; 
        10'b0010010001: data <= 21'h1ffc6f; 
        10'b0010010010: data <= 21'h1ffcd4; 
        10'b0010010011: data <= 21'h1ffc7b; 
        10'b0010010100: data <= 21'h1ff4a3; 
        10'b0010010101: data <= 21'h1ff4dd; 
        10'b0010010110: data <= 21'h1ff3f8; 
        10'b0010010111: data <= 21'h1ff029; 
        10'b0010011000: data <= 21'h1fec27; 
        10'b0010011001: data <= 21'h1fe885; 
        10'b0010011010: data <= 21'h1fdc29; 
        10'b0010011011: data <= 21'h1fd94d; 
        10'b0010011100: data <= 21'h1fcf18; 
        10'b0010011101: data <= 21'h1fdfc3; 
        10'b0010011110: data <= 21'h1febaf; 
        10'b0010011111: data <= 21'h1ff628; 
        10'b0010100000: data <= 21'h1ff59d; 
        10'b0010100001: data <= 21'h1ff27a; 
        10'b0010100010: data <= 21'h1ff369; 
        10'b0010100011: data <= 21'h1ff706; 
        10'b0010100100: data <= 21'h1ffc6d; 
        10'b0010100101: data <= 21'h1ffe58; 
        10'b0010100110: data <= 21'h00008c; 
        10'b0010100111: data <= 21'h00032b; 
        10'b0010101000: data <= 21'h000410; 
        10'b0010101001: data <= 21'h00042e; 
        10'b0010101010: data <= 21'h1ffd61; 
        10'b0010101011: data <= 21'h000437; 
        10'b0010101100: data <= 21'h0002af; 
        10'b0010101101: data <= 21'h1ff3e9; 
        10'b0010101110: data <= 21'h1ff149; 
        10'b0010101111: data <= 21'h1feeaa; 
        10'b0010110000: data <= 21'h1fec76; 
        10'b0010110001: data <= 21'h1fe807; 
        10'b0010110010: data <= 21'h1fee65; 
        10'b0010110011: data <= 21'h1ffa5f; 
        10'b0010110100: data <= 21'h00016a; 
        10'b0010110101: data <= 21'h0015a4; 
        10'b0010110110: data <= 21'h00204a; 
        10'b0010110111: data <= 21'h0019af; 
        10'b0010111000: data <= 21'h0011ff; 
        10'b0010111001: data <= 21'h000ef4; 
        10'b0010111010: data <= 21'h0012f6; 
        10'b0010111011: data <= 21'h1ffcce; 
        10'b0010111100: data <= 21'h1ffb6f; 
        10'b0010111101: data <= 21'h1ff193; 
        10'b0010111110: data <= 21'h1fe625; 
        10'b0010111111: data <= 21'h1fe7ef; 
        10'b0011000000: data <= 21'h1ff238; 
        10'b0011000001: data <= 21'h1ff94b; 
        10'b0011000010: data <= 21'h1ffefc; 
        10'b0011000011: data <= 21'h000230; 
        10'b0011000100: data <= 21'h00063c; 
        10'b0011000101: data <= 21'h1fffc6; 
        10'b0011000110: data <= 21'h1ffdf9; 
        10'b0011000111: data <= 21'h1ffdc1; 
        10'b0011001000: data <= 21'h1ff22e; 
        10'b0011001001: data <= 21'h1feafc; 
        10'b0011001010: data <= 21'h1fe741; 
        10'b0011001011: data <= 21'h1fe28d; 
        10'b0011001100: data <= 21'h1fe425; 
        10'b0011001101: data <= 21'h1ff62e; 
        10'b0011001110: data <= 21'h1fff33; 
        10'b0011001111: data <= 21'h0007a2; 
        10'b0011010000: data <= 21'h001d54; 
        10'b0011010001: data <= 21'h002303; 
        10'b0011010010: data <= 21'h003000; 
        10'b0011010011: data <= 21'h00303f; 
        10'b0011010100: data <= 21'h003232; 
        10'b0011010101: data <= 21'h0016c0; 
        10'b0011010110: data <= 21'h001121; 
        10'b0011010111: data <= 21'h0001da; 
        10'b0011011000: data <= 21'h000473; 
        10'b0011011001: data <= 21'h00050a; 
        10'b0011011010: data <= 21'h1feeb6; 
        10'b0011011011: data <= 21'h1fe107; 
        10'b0011011100: data <= 21'h1fedbe; 
        10'b0011011101: data <= 21'h1ffb70; 
        10'b0011011110: data <= 21'h1ffb53; 
        10'b0011011111: data <= 21'h000418; 
        10'b0011100000: data <= 21'h00060d; 
        10'b0011100001: data <= 21'h000617; 
        10'b0011100010: data <= 21'h000318; 
        10'b0011100011: data <= 21'h1ffe23; 
        10'b0011100100: data <= 21'h1ff19d; 
        10'b0011100101: data <= 21'h1fea3a; 
        10'b0011100110: data <= 21'h1fe6a6; 
        10'b0011100111: data <= 21'h1fdc8e; 
        10'b0011101000: data <= 21'h1ff6a2; 
        10'b0011101001: data <= 21'h1ffbaa; 
        10'b0011101010: data <= 21'h1ffafa; 
        10'b0011101011: data <= 21'h1ff5ea; 
        10'b0011101100: data <= 21'h1fff3b; 
        10'b0011101101: data <= 21'h000e0d; 
        10'b0011101110: data <= 21'h002922; 
        10'b0011101111: data <= 21'h0016b4; 
        10'b0011110000: data <= 21'h00171e; 
        10'b0011110001: data <= 21'h0004bc; 
        10'b0011110010: data <= 21'h0001d3; 
        10'b0011110011: data <= 21'h00013a; 
        10'b0011110100: data <= 21'h1ff866; 
        10'b0011110101: data <= 21'h0003f2; 
        10'b0011110110: data <= 21'h1ff642; 
        10'b0011110111: data <= 21'h1fe74b; 
        10'b0011111000: data <= 21'h1feb21; 
        10'b0011111001: data <= 21'h1ff5fe; 
        10'b0011111010: data <= 21'h1ffba1; 
        10'b0011111011: data <= 21'h0005a4; 
        10'b0011111100: data <= 21'h0001d6; 
        10'b0011111101: data <= 21'h000119; 
        10'b0011111110: data <= 21'h000069; 
        10'b0011111111: data <= 21'h1ff5b6; 
        10'b0100000000: data <= 21'h1fe991; 
        10'b0100000001: data <= 21'h1feecb; 
        10'b0100000010: data <= 21'h1ffb21; 
        10'b0100000011: data <= 21'h1ff623; 
        10'b0100000100: data <= 21'h1ffa22; 
        10'b0100000101: data <= 21'h1ffd57; 
        10'b0100000110: data <= 21'h000a8c; 
        10'b0100000111: data <= 21'h00065b; 
        10'b0100001000: data <= 21'h0001dd; 
        10'b0100001001: data <= 21'h0010fd; 
        10'b0100001010: data <= 21'h001c73; 
        10'b0100001011: data <= 21'h00195e; 
        10'b0100001100: data <= 21'h1fff03; 
        10'b0100001101: data <= 21'h1ff8ba; 
        10'b0100001110: data <= 21'h000048; 
        10'b0100001111: data <= 21'h1ff0db; 
        10'b0100010000: data <= 21'h1ff993; 
        10'b0100010001: data <= 21'h1ff01f; 
        10'b0100010010: data <= 21'h1fef00; 
        10'b0100010011: data <= 21'h1feddd; 
        10'b0100010100: data <= 21'h1ff3a2; 
        10'b0100010101: data <= 21'h1ffa99; 
        10'b0100010110: data <= 21'h1ffc14; 
        10'b0100010111: data <= 21'h000502; 
        10'b0100011000: data <= 21'h000116; 
        10'b0100011001: data <= 21'h1fffc8; 
        10'b0100011010: data <= 21'h1ffd96; 
        10'b0100011011: data <= 21'h1ffc0f; 
        10'b0100011100: data <= 21'h1feeb8; 
        10'b0100011101: data <= 21'h1ff6f6; 
        10'b0100011110: data <= 21'h00086e; 
        10'b0100011111: data <= 21'h000b0a; 
        10'b0100100000: data <= 21'h001667; 
        10'b0100100001: data <= 21'h00163f; 
        10'b0100100010: data <= 21'h001327; 
        10'b0100100011: data <= 21'h001cd8; 
        10'b0100100100: data <= 21'h000e85; 
        10'b0100100101: data <= 21'h00036b; 
        10'b0100100110: data <= 21'h0003b5; 
        10'b0100100111: data <= 21'h1ff166; 
        10'b0100101000: data <= 21'h1ff74c; 
        10'b0100101001: data <= 21'h1ffe47; 
        10'b0100101010: data <= 21'h000a2c; 
        10'b0100101011: data <= 21'h1fffc8; 
        10'b0100101100: data <= 21'h00082e; 
        10'b0100101101: data <= 21'h1ffb1d; 
        10'b0100101110: data <= 21'h1ff5f6; 
        10'b0100101111: data <= 21'h1ff686; 
        10'b0100110000: data <= 21'h1ff3f8; 
        10'b0100110001: data <= 21'h1ffc91; 
        10'b0100110010: data <= 21'h1ffb74; 
        10'b0100110011: data <= 21'h0002e0; 
        10'b0100110100: data <= 21'h1fff0d; 
        10'b0100110101: data <= 21'h000127; 
        10'b0100110110: data <= 21'h1ffd66; 
        10'b0100110111: data <= 21'h1ffe59; 
        10'b0100111000: data <= 21'h1ffb43; 
        10'b0100111001: data <= 21'h000fe6; 
        10'b0100111010: data <= 21'h0024c9; 
        10'b0100111011: data <= 21'h001b74; 
        10'b0100111100: data <= 21'h002b23; 
        10'b0100111101: data <= 21'h00114b; 
        10'b0100111110: data <= 21'h0011ee; 
        10'b0100111111: data <= 21'h001ecd; 
        10'b0101000000: data <= 21'h1ff634; 
        10'b0101000001: data <= 21'h1ff7ac; 
        10'b0101000010: data <= 21'h1ffb80; 
        10'b0101000011: data <= 21'h00022d; 
        10'b0101000100: data <= 21'h000be8; 
        10'b0101000101: data <= 21'h0029b1; 
        10'b0101000110: data <= 21'h0013b2; 
        10'b0101000111: data <= 21'h0013f7; 
        10'b0101001000: data <= 21'h0020bd; 
        10'b0101001001: data <= 21'h0017b1; 
        10'b0101001010: data <= 21'h000dd7; 
        10'b0101001011: data <= 21'h0002dd; 
        10'b0101001100: data <= 21'h1ffdbc; 
        10'b0101001101: data <= 21'h1ffa5c; 
        10'b0101001110: data <= 21'h1fffc1; 
        10'b0101001111: data <= 21'h000006; 
        10'b0101010000: data <= 21'h00029b; 
        10'b0101010001: data <= 21'h00055e; 
        10'b0101010010: data <= 21'h1ffc4c; 
        10'b0101010011: data <= 21'h1ffa18; 
        10'b0101010100: data <= 21'h000d6c; 
        10'b0101010101: data <= 21'h0022e1; 
        10'b0101010110: data <= 21'h00285b; 
        10'b0101010111: data <= 21'h0017f0; 
        10'b0101011000: data <= 21'h001deb; 
        10'b0101011001: data <= 21'h002496; 
        10'b0101011010: data <= 21'h00175d; 
        10'b0101011011: data <= 21'h000046; 
        10'b0101011100: data <= 21'h1fe890; 
        10'b0101011101: data <= 21'h00144e; 
        10'b0101011110: data <= 21'h002bde; 
        10'b0101011111: data <= 21'h0022b5; 
        10'b0101100000: data <= 21'h001dac; 
        10'b0101100001: data <= 21'h002d5f; 
        10'b0101100010: data <= 21'h002db2; 
        10'b0101100011: data <= 21'h002f6b; 
        10'b0101100100: data <= 21'h0030c0; 
        10'b0101100101: data <= 21'h002094; 
        10'b0101100110: data <= 21'h000fab; 
        10'b0101100111: data <= 21'h00006a; 
        10'b0101101000: data <= 21'h1ff8bf; 
        10'b0101101001: data <= 21'h00012f; 
        10'b0101101010: data <= 21'h0002a2; 
        10'b0101101011: data <= 21'h0002d9; 
        10'b0101101100: data <= 21'h000608; 
        10'b0101101101: data <= 21'h0003b4; 
        10'b0101101110: data <= 21'h1ffaed; 
        10'b0101101111: data <= 21'h0001e8; 
        10'b0101110000: data <= 21'h00144c; 
        10'b0101110001: data <= 21'h001e85; 
        10'b0101110010: data <= 21'h001cc3; 
        10'b0101110011: data <= 21'h0012e1; 
        10'b0101110100: data <= 21'h0017b5; 
        10'b0101110101: data <= 21'h000f38; 
        10'b0101110110: data <= 21'h000dc1; 
        10'b0101110111: data <= 21'h1ff8e1; 
        10'b0101111000: data <= 21'h1ff3b1; 
        10'b0101111001: data <= 21'h001fea; 
        10'b0101111010: data <= 21'h002bc6; 
        10'b0101111011: data <= 21'h001fb8; 
        10'b0101111100: data <= 21'h00248e; 
        10'b0101111101: data <= 21'h0020c5; 
        10'b0101111110: data <= 21'h002cf5; 
        10'b0101111111: data <= 21'h002dbd; 
        10'b0110000000: data <= 21'h0023c0; 
        10'b0110000001: data <= 21'h0014e1; 
        10'b0110000010: data <= 21'h000132; 
        10'b0110000011: data <= 21'h1ff1c7; 
        10'b0110000100: data <= 21'h1ff7b7; 
        10'b0110000101: data <= 21'h1ffd6d; 
        10'b0110000110: data <= 21'h0002b3; 
        10'b0110000111: data <= 21'h0002bd; 
        10'b0110001000: data <= 21'h000137; 
        10'b0110001001: data <= 21'h00009a; 
        10'b0110001010: data <= 21'h000426; 
        10'b0110001011: data <= 21'h0002a3; 
        10'b0110001100: data <= 21'h000949; 
        10'b0110001101: data <= 21'h0008c0; 
        10'b0110001110: data <= 21'h0017d5; 
        10'b0110001111: data <= 21'h0010ac; 
        10'b0110010000: data <= 21'h00081b; 
        10'b0110010001: data <= 21'h1fffea; 
        10'b0110010010: data <= 21'h0002f7; 
        10'b0110010011: data <= 21'h1ffe86; 
        10'b0110010100: data <= 21'h1ff701; 
        10'b0110010101: data <= 21'h000a59; 
        10'b0110010110: data <= 21'h0005e1; 
        10'b0110010111: data <= 21'h001bfe; 
        10'b0110011000: data <= 21'h001db0; 
        10'b0110011001: data <= 21'h001dbb; 
        10'b0110011010: data <= 21'h00143f; 
        10'b0110011011: data <= 21'h000d04; 
        10'b0110011100: data <= 21'h00103d; 
        10'b0110011101: data <= 21'h00004c; 
        10'b0110011110: data <= 21'h1fef9c; 
        10'b0110011111: data <= 21'h1fe82e; 
        10'b0110100000: data <= 21'h1ff626; 
        10'b0110100001: data <= 21'h0001a5; 
        10'b0110100010: data <= 21'h0000f0; 
        10'b0110100011: data <= 21'h00011c; 
        10'b0110100100: data <= 21'h000490; 
        10'b0110100101: data <= 21'h000429; 
        10'b0110100110: data <= 21'h0002c1; 
        10'b0110100111: data <= 21'h1ffcac; 
        10'b0110101000: data <= 21'h0000ae; 
        10'b0110101001: data <= 21'h000a9a; 
        10'b0110101010: data <= 21'h000a27; 
        10'b0110101011: data <= 21'h0006b4; 
        10'b0110101100: data <= 21'h0006d7; 
        10'b0110101101: data <= 21'h1ff36f; 
        10'b0110101110: data <= 21'h1ffa2a; 
        10'b0110101111: data <= 21'h1ffa1f; 
        10'b0110110000: data <= 21'h1ff73a; 
        10'b0110110001: data <= 21'h1ff936; 
        10'b0110110010: data <= 21'h1ff7c6; 
        10'b0110110011: data <= 21'h001e94; 
        10'b0110110100: data <= 21'h002cc5; 
        10'b0110110101: data <= 21'h002ae9; 
        10'b0110110110: data <= 21'h00157c; 
        10'b0110110111: data <= 21'h000213; 
        10'b0110111000: data <= 21'h1ff6ab; 
        10'b0110111001: data <= 21'h1fe765; 
        10'b0110111010: data <= 21'h1fe14e; 
        10'b0110111011: data <= 21'h1fea13; 
        10'b0110111100: data <= 21'h1ff63e; 
        10'b0110111101: data <= 21'h00002e; 
        10'b0110111110: data <= 21'h000282; 
        10'b0110111111: data <= 21'h1fffa5; 
        10'b0111000000: data <= 21'h000541; 
        10'b0111000001: data <= 21'h000070; 
        10'b0111000010: data <= 21'h1ffc3c; 
        10'b0111000011: data <= 21'h1fff09; 
        10'b0111000100: data <= 21'h000055; 
        10'b0111000101: data <= 21'h00032e; 
        10'b0111000110: data <= 21'h1ff7cc; 
        10'b0111000111: data <= 21'h00067b; 
        10'b0111001000: data <= 21'h001267; 
        10'b0111001001: data <= 21'h1ffbb0; 
        10'b0111001010: data <= 21'h000a71; 
        10'b0111001011: data <= 21'h000ece; 
        10'b0111001100: data <= 21'h1ffdfb; 
        10'b0111001101: data <= 21'h1fef29; 
        10'b0111001110: data <= 21'h1ffd2e; 
        10'b0111001111: data <= 21'h0010fa; 
        10'b0111010000: data <= 21'h001e8d; 
        10'b0111010001: data <= 21'h001e5a; 
        10'b0111010010: data <= 21'h000794; 
        10'b0111010011: data <= 21'h1feebd; 
        10'b0111010100: data <= 21'h1fe35b; 
        10'b0111010101: data <= 21'h1fd865; 
        10'b0111010110: data <= 21'h1fe432; 
        10'b0111010111: data <= 21'h1fe969; 
        10'b0111011000: data <= 21'h1ff10d; 
        10'b0111011001: data <= 21'h00007f; 
        10'b0111011010: data <= 21'h1ffcbd; 
        10'b0111011011: data <= 21'h0002d3; 
        10'b0111011100: data <= 21'h0001bc; 
        10'b0111011101: data <= 21'h1ffed7; 
        10'b0111011110: data <= 21'h1ffbe4; 
        10'b0111011111: data <= 21'h1ff9fe; 
        10'b0111100000: data <= 21'h1ff4bf; 
        10'b0111100001: data <= 21'h1ff24f; 
        10'b0111100010: data <= 21'h1ff4b7; 
        10'b0111100011: data <= 21'h000517; 
        10'b0111100100: data <= 21'h0009ea; 
        10'b0111100101: data <= 21'h000b4a; 
        10'b0111100110: data <= 21'h001136; 
        10'b0111100111: data <= 21'h00190c; 
        10'b0111101000: data <= 21'h000f46; 
        10'b0111101001: data <= 21'h000719; 
        10'b0111101010: data <= 21'h0009b4; 
        10'b0111101011: data <= 21'h0018ea; 
        10'b0111101100: data <= 21'h000766; 
        10'b0111101101: data <= 21'h1ffaf3; 
        10'b0111101110: data <= 21'h1ff4fd; 
        10'b0111101111: data <= 21'h1fe6b4; 
        10'b0111110000: data <= 21'h1fe707; 
        10'b0111110001: data <= 21'h1fe51e; 
        10'b0111110010: data <= 21'h1fe6b8; 
        10'b0111110011: data <= 21'h1fed63; 
        10'b0111110100: data <= 21'h1ff272; 
        10'b0111110101: data <= 21'h00015a; 
        10'b0111110110: data <= 21'h000165; 
        10'b0111110111: data <= 21'h1ffece; 
        10'b0111111000: data <= 21'h0004da; 
        10'b0111111001: data <= 21'h1ffffc; 
        10'b0111111010: data <= 21'h1ffd2b; 
        10'b0111111011: data <= 21'h1ffee0; 
        10'b0111111100: data <= 21'h1ff61a; 
        10'b0111111101: data <= 21'h1fe947; 
        10'b0111111110: data <= 21'h1fe8d7; 
        10'b0111111111: data <= 21'h1fe947; 
        10'b1000000000: data <= 21'h1ff674; 
        10'b1000000001: data <= 21'h0003ca; 
        10'b1000000010: data <= 21'h001b72; 
        10'b1000000011: data <= 21'h00162f; 
        10'b1000000100: data <= 21'h1ff276; 
        10'b1000000101: data <= 21'h1ff242; 
        10'b1000000110: data <= 21'h0000da; 
        10'b1000000111: data <= 21'h00107e; 
        10'b1000001000: data <= 21'h1ff5e4; 
        10'b1000001001: data <= 21'h1ff478; 
        10'b1000001010: data <= 21'h1fea68; 
        10'b1000001011: data <= 21'h1ff301; 
        10'b1000001100: data <= 21'h1ff3d1; 
        10'b1000001101: data <= 21'h1fecfb; 
        10'b1000001110: data <= 21'h1febfc; 
        10'b1000001111: data <= 21'h1feb0b; 
        10'b1000010000: data <= 21'h1ff12d; 
        10'b1000010001: data <= 21'h1ffda4; 
        10'b1000010010: data <= 21'h00004c; 
        10'b1000010011: data <= 21'h000470; 
        10'b1000010100: data <= 21'h000326; 
        10'b1000010101: data <= 21'h000649; 
        10'b1000010110: data <= 21'h00011e; 
        10'b1000010111: data <= 21'h1ffa90; 
        10'b1000011000: data <= 21'h1ff6ea; 
        10'b1000011001: data <= 21'h1fefec; 
        10'b1000011010: data <= 21'h1fe696; 
        10'b1000011011: data <= 21'h1fe5eb; 
        10'b1000011100: data <= 21'h1fe4fe; 
        10'b1000011101: data <= 21'h1fe536; 
        10'b1000011110: data <= 21'h1fe205; 
        10'b1000011111: data <= 21'h1fe6ad; 
        10'b1000100000: data <= 21'h1fdf37; 
        10'b1000100001: data <= 21'h1fe915; 
        10'b1000100010: data <= 21'h1fecb0; 
        10'b1000100011: data <= 21'h1fea07; 
        10'b1000100100: data <= 21'h1fed09; 
        10'b1000100101: data <= 21'h1ff9ce; 
        10'b1000100110: data <= 21'h1ff192; 
        10'b1000100111: data <= 21'h1ffbf9; 
        10'b1000101000: data <= 21'h1ff659; 
        10'b1000101001: data <= 21'h1ff491; 
        10'b1000101010: data <= 21'h1ff534; 
        10'b1000101011: data <= 21'h1ff666; 
        10'b1000101100: data <= 21'h1ff9f6; 
        10'b1000101101: data <= 21'h0001bd; 
        10'b1000101110: data <= 21'h1ffe1a; 
        10'b1000101111: data <= 21'h0000ac; 
        10'b1000110000: data <= 21'h1ffed1; 
        10'b1000110001: data <= 21'h0000e1; 
        10'b1000110010: data <= 21'h0002ac; 
        10'b1000110011: data <= 21'h000034; 
        10'b1000110100: data <= 21'h1ff698; 
        10'b1000110101: data <= 21'h1ff079; 
        10'b1000110110: data <= 21'h1fe874; 
        10'b1000110111: data <= 21'h1fdb1e; 
        10'b1000111000: data <= 21'h1fd5c2; 
        10'b1000111001: data <= 21'h1fd09e; 
        10'b1000111010: data <= 21'h1fbfda; 
        10'b1000111011: data <= 21'h1fcee7; 
        10'b1000111100: data <= 21'h1fd029; 
        10'b1000111101: data <= 21'h1ff058; 
        10'b1000111110: data <= 21'h1fea0b; 
        10'b1000111111: data <= 21'h1ff5b0; 
        10'b1001000000: data <= 21'h1ff3a2; 
        10'b1001000001: data <= 21'h1ffcab; 
        10'b1001000010: data <= 21'h1feaf9; 
        10'b1001000011: data <= 21'h1ff913; 
        10'b1001000100: data <= 21'h1ff7a8; 
        10'b1001000101: data <= 21'h1ff299; 
        10'b1001000110: data <= 21'h1ffc39; 
        10'b1001000111: data <= 21'h1ff994; 
        10'b1001001000: data <= 21'h0000a5; 
        10'b1001001001: data <= 21'h00055a; 
        10'b1001001010: data <= 21'h00033a; 
        10'b1001001011: data <= 21'h000103; 
        10'b1001001100: data <= 21'h00006e; 
        10'b1001001101: data <= 21'h000001; 
        10'b1001001110: data <= 21'h00055a; 
        10'b1001001111: data <= 21'h1ffa54; 
        10'b1001010000: data <= 21'h1ff9ac; 
        10'b1001010001: data <= 21'h1ff0b1; 
        10'b1001010010: data <= 21'h1fea60; 
        10'b1001010011: data <= 21'h1fdea0; 
        10'b1001010100: data <= 21'h1fda1d; 
        10'b1001010101: data <= 21'h1fd652; 
        10'b1001010110: data <= 21'h1fd44f; 
        10'b1001010111: data <= 21'h1fd8b5; 
        10'b1001011000: data <= 21'h1fe6f8; 
        10'b1001011001: data <= 21'h1fe74b; 
        10'b1001011010: data <= 21'h1fe6e3; 
        10'b1001011011: data <= 21'h1ff197; 
        10'b1001011100: data <= 21'h1ff064; 
        10'b1001011101: data <= 21'h1fe881; 
        10'b1001011110: data <= 21'h1fe3a6; 
        10'b1001011111: data <= 21'h1ff3fc; 
        10'b1001100000: data <= 21'h1ff94d; 
        10'b1001100001: data <= 21'h1ffc23; 
        10'b1001100010: data <= 21'h0001e4; 
        10'b1001100011: data <= 21'h1fff77; 
        10'b1001100100: data <= 21'h000267; 
        10'b1001100101: data <= 21'h000349; 
        10'b1001100110: data <= 21'h00002f; 
        10'b1001100111: data <= 21'h000065; 
        10'b1001101000: data <= 21'h00041b; 
        10'b1001101001: data <= 21'h000106; 
        10'b1001101010: data <= 21'h000129; 
        10'b1001101011: data <= 21'h0003ee; 
        10'b1001101100: data <= 21'h1ffd79; 
        10'b1001101101: data <= 21'h1ff3a2; 
        10'b1001101110: data <= 21'h1fec36; 
        10'b1001101111: data <= 21'h1fe515; 
        10'b1001110000: data <= 21'h1febf8; 
        10'b1001110001: data <= 21'h1feb13; 
        10'b1001110010: data <= 21'h1fe926; 
        10'b1001110011: data <= 21'h1ff092; 
        10'b1001110100: data <= 21'h1feea8; 
        10'b1001110101: data <= 21'h1fe8ec; 
        10'b1001110110: data <= 21'h1fec9a; 
        10'b1001110111: data <= 21'h1fe4d0; 
        10'b1001111000: data <= 21'h1fe1ed; 
        10'b1001111001: data <= 21'h1fe285; 
        10'b1001111010: data <= 21'h1fe77c; 
        10'b1001111011: data <= 21'h1fea34; 
        10'b1001111100: data <= 21'h1ffa04; 
        10'b1001111101: data <= 21'h000756; 
        10'b1001111110: data <= 21'h000414; 
        10'b1001111111: data <= 21'h00050f; 
        10'b1010000000: data <= 21'h000846; 
        10'b1010000001: data <= 21'h0001bc; 
        10'b1010000010: data <= 21'h0001ee; 
        10'b1010000011: data <= 21'h000304; 
        10'b1010000100: data <= 21'h0004d2; 
        10'b1010000101: data <= 21'h0003c8; 
        10'b1010000110: data <= 21'h00016a; 
        10'b1010000111: data <= 21'h1ffe1c; 
        10'b1010001000: data <= 21'h1ffc87; 
        10'b1010001001: data <= 21'h1ff55d; 
        10'b1010001010: data <= 21'h1ff3a2; 
        10'b1010001011: data <= 21'h1fefa7; 
        10'b1010001100: data <= 21'h1ffec4; 
        10'b1010001101: data <= 21'h1ff964; 
        10'b1010001110: data <= 21'h1ffab4; 
        10'b1010001111: data <= 21'h1fec2f; 
        10'b1010010000: data <= 21'h1fefda; 
        10'b1010010001: data <= 21'h1feba1; 
        10'b1010010010: data <= 21'h1feec7; 
        10'b1010010011: data <= 21'h1fe298; 
        10'b1010010100: data <= 21'h1fe042; 
        10'b1010010101: data <= 21'h1fe40f; 
        10'b1010010110: data <= 21'h1fee98; 
        10'b1010010111: data <= 21'h1ffe4d; 
        10'b1010011000: data <= 21'h0006d1; 
        10'b1010011001: data <= 21'h000fd2; 
        10'b1010011010: data <= 21'h0016cd; 
        10'b1010011011: data <= 21'h001319; 
        10'b1010011100: data <= 21'h0008f0; 
        10'b1010011101: data <= 21'h1fff64; 
        10'b1010011110: data <= 21'h000669; 
        10'b1010011111: data <= 21'h1fff41; 
        10'b1010100000: data <= 21'h1ffffb; 
        10'b1010100001: data <= 21'h1ffd79; 
        10'b1010100010: data <= 21'h1fff52; 
        10'b1010100011: data <= 21'h000566; 
        10'b1010100100: data <= 21'h0003e2; 
        10'b1010100101: data <= 21'h000615; 
        10'b1010100110: data <= 21'h00046b; 
        10'b1010100111: data <= 21'h00066b; 
        10'b1010101000: data <= 21'h000911; 
        10'b1010101001: data <= 21'h0004e5; 
        10'b1010101010: data <= 21'h1ffcc5; 
        10'b1010101011: data <= 21'h1ff5d7; 
        10'b1010101100: data <= 21'h1fff48; 
        10'b1010101101: data <= 21'h1ff068; 
        10'b1010101110: data <= 21'h1fec4a; 
        10'b1010101111: data <= 21'h1feb30; 
        10'b1010110000: data <= 21'h1ff690; 
        10'b1010110001: data <= 21'h0006d9; 
        10'b1010110010: data <= 21'h000bb0; 
        10'b1010110011: data <= 21'h000c15; 
        10'b1010110100: data <= 21'h001b96; 
        10'b1010110101: data <= 21'h001daf; 
        10'b1010110110: data <= 21'h001116; 
        10'b1010110111: data <= 21'h000a72; 
        10'b1010111000: data <= 21'h00083f; 
        10'b1010111001: data <= 21'h1ffe62; 
        10'b1010111010: data <= 21'h0003af; 
        10'b1010111011: data <= 21'h1fffc1; 
        10'b1010111100: data <= 21'h000158; 
        10'b1010111101: data <= 21'h00055b; 
        10'b1010111110: data <= 21'h00055e; 
        10'b1010111111: data <= 21'h1fff6f; 
        10'b1011000000: data <= 21'h000081; 
        10'b1011000001: data <= 21'h00092b; 
        10'b1011000010: data <= 21'h0006f2; 
        10'b1011000011: data <= 21'h00140a; 
        10'b1011000100: data <= 21'h0015f6; 
        10'b1011000101: data <= 21'h00165c; 
        10'b1011000110: data <= 21'h001359; 
        10'b1011000111: data <= 21'h0007ae; 
        10'b1011001000: data <= 21'h00145a; 
        10'b1011001001: data <= 21'h001227; 
        10'b1011001010: data <= 21'h001161; 
        10'b1011001011: data <= 21'h001056; 
        10'b1011001100: data <= 21'h001e85; 
        10'b1011001101: data <= 21'h00212a; 
        10'b1011001110: data <= 21'h00247a; 
        10'b1011001111: data <= 21'h002612; 
        10'b1011010000: data <= 21'h002a7f; 
        10'b1011010001: data <= 21'h001e27; 
        10'b1011010010: data <= 21'h000bc4; 
        10'b1011010011: data <= 21'h000594; 
        10'b1011010100: data <= 21'h1fff41; 
        10'b1011010101: data <= 21'h1fff8d; 
        10'b1011010110: data <= 21'h000190; 
        10'b1011010111: data <= 21'h000150; 
        10'b1011011000: data <= 21'h00003a; 
        10'b1011011001: data <= 21'h0004e1; 
        10'b1011011010: data <= 21'h00014f; 
        10'b1011011011: data <= 21'h1ffe39; 
        10'b1011011100: data <= 21'h0004e8; 
        10'b1011011101: data <= 21'h00079a; 
        10'b1011011110: data <= 21'h000aa9; 
        10'b1011011111: data <= 21'h000ecf; 
        10'b1011100000: data <= 21'h0010dc; 
        10'b1011100001: data <= 21'h001992; 
        10'b1011100010: data <= 21'h001a62; 
        10'b1011100011: data <= 21'h001da2; 
        10'b1011100100: data <= 21'h002318; 
        10'b1011100101: data <= 21'h002367; 
        10'b1011100110: data <= 21'h002b59; 
        10'b1011100111: data <= 21'h001901; 
        10'b1011101000: data <= 21'h001121; 
        10'b1011101001: data <= 21'h000e77; 
        10'b1011101010: data <= 21'h001555; 
        10'b1011101011: data <= 21'h001707; 
        10'b1011101100: data <= 21'h0010b8; 
        10'b1011101101: data <= 21'h000ba5; 
        10'b1011101110: data <= 21'h0004d8; 
        10'b1011101111: data <= 21'h0001bf; 
        10'b1011110000: data <= 21'h000116; 
        10'b1011110001: data <= 21'h0001ee; 
        10'b1011110010: data <= 21'h1ffe2b; 
        10'b1011110011: data <= 21'h000111; 
        10'b1011110100: data <= 21'h1ffed4; 
        10'b1011110101: data <= 21'h00023b; 
        10'b1011110110: data <= 21'h1ffdfd; 
        10'b1011110111: data <= 21'h0005e9; 
        10'b1011111000: data <= 21'h000364; 
        10'b1011111001: data <= 21'h0001e0; 
        10'b1011111010: data <= 21'h1fff29; 
        10'b1011111011: data <= 21'h0005bf; 
        10'b1011111100: data <= 21'h0004db; 
        10'b1011111101: data <= 21'h000352; 
        10'b1011111110: data <= 21'h1ffeee; 
        10'b1011111111: data <= 21'h1ffecd; 
        10'b1100000000: data <= 21'h000124; 
        10'b1100000001: data <= 21'h1ffeef; 
        10'b1100000010: data <= 21'h00013d; 
        10'b1100000011: data <= 21'h0003b0; 
        10'b1100000100: data <= 21'h000057; 
        10'b1100000101: data <= 21'h000203; 
        10'b1100000110: data <= 21'h00068f; 
        10'b1100000111: data <= 21'h0005d7; 
        10'b1100001000: data <= 21'h00034a; 
        10'b1100001001: data <= 21'h000203; 
        10'b1100001010: data <= 21'h1ffe5f; 
        10'b1100001011: data <= 21'h00067b; 
        10'b1100001100: data <= 21'h000386; 
        10'b1100001101: data <= 21'h1ffecd; 
        10'b1100001110: data <= 21'h000073; 
        10'b1100001111: data <= 21'h1fff58; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 16) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 22'h00090a; 
        10'b0000000001: data <= 22'h0007eb; 
        10'b0000000010: data <= 22'h3ffd90; 
        10'b0000000011: data <= 22'h00058d; 
        10'b0000000100: data <= 22'h00051e; 
        10'b0000000101: data <= 22'h000849; 
        10'b0000000110: data <= 22'h3ffce5; 
        10'b0000000111: data <= 22'h00018b; 
        10'b0000001000: data <= 22'h00098d; 
        10'b0000001001: data <= 22'h3ffc19; 
        10'b0000001010: data <= 22'h3ffed9; 
        10'b0000001011: data <= 22'h00042c; 
        10'b0000001100: data <= 22'h000c0e; 
        10'b0000001101: data <= 22'h0007da; 
        10'b0000001110: data <= 22'h3ffb15; 
        10'b0000001111: data <= 22'h3ffdba; 
        10'b0000010000: data <= 22'h3ffd7f; 
        10'b0000010001: data <= 22'h0004be; 
        10'b0000010010: data <= 22'h0008b6; 
        10'b0000010011: data <= 22'h0000a4; 
        10'b0000010100: data <= 22'h0000de; 
        10'b0000010101: data <= 22'h3fff5e; 
        10'b0000010110: data <= 22'h3ffc24; 
        10'b0000010111: data <= 22'h000159; 
        10'b0000011000: data <= 22'h0009c7; 
        10'b0000011001: data <= 22'h0002f4; 
        10'b0000011010: data <= 22'h3ffb8a; 
        10'b0000011011: data <= 22'h0004da; 
        10'b0000011100: data <= 22'h00081a; 
        10'b0000011101: data <= 22'h0006c7; 
        10'b0000011110: data <= 22'h000344; 
        10'b0000011111: data <= 22'h3ffe1c; 
        10'b0000100000: data <= 22'h3ffb4d; 
        10'b0000100001: data <= 22'h3ffc29; 
        10'b0000100010: data <= 22'h3fff39; 
        10'b0000100011: data <= 22'h000c20; 
        10'b0000100100: data <= 22'h3ffb6d; 
        10'b0000100101: data <= 22'h0009d7; 
        10'b0000100110: data <= 22'h0003ca; 
        10'b0000100111: data <= 22'h000612; 
        10'b0000101000: data <= 22'h0004c0; 
        10'b0000101001: data <= 22'h0006e2; 
        10'b0000101010: data <= 22'h000030; 
        10'b0000101011: data <= 22'h3ffaab; 
        10'b0000101100: data <= 22'h3ffd47; 
        10'b0000101101: data <= 22'h00077d; 
        10'b0000101110: data <= 22'h3fffad; 
        10'b0000101111: data <= 22'h000221; 
        10'b0000110000: data <= 22'h00097f; 
        10'b0000110001: data <= 22'h3fff49; 
        10'b0000110010: data <= 22'h0001aa; 
        10'b0000110011: data <= 22'h0000dc; 
        10'b0000110100: data <= 22'h00053c; 
        10'b0000110101: data <= 22'h000a2d; 
        10'b0000110110: data <= 22'h3fffe0; 
        10'b0000110111: data <= 22'h00022b; 
        10'b0000111000: data <= 22'h000ab7; 
        10'b0000111001: data <= 22'h000afe; 
        10'b0000111010: data <= 22'h0000d3; 
        10'b0000111011: data <= 22'h00077d; 
        10'b0000111100: data <= 22'h000915; 
        10'b0000111101: data <= 22'h3fff93; 
        10'b0000111110: data <= 22'h3ffeee; 
        10'b0000111111: data <= 22'h000341; 
        10'b0001000000: data <= 22'h00091d; 
        10'b0001000001: data <= 22'h3ffeb1; 
        10'b0001000010: data <= 22'h3ffd39; 
        10'b0001000011: data <= 22'h0006f8; 
        10'b0001000100: data <= 22'h00041d; 
        10'b0001000101: data <= 22'h0008b4; 
        10'b0001000110: data <= 22'h3ffadf; 
        10'b0001000111: data <= 22'h000930; 
        10'b0001001000: data <= 22'h3ffcb1; 
        10'b0001001001: data <= 22'h3ffc7c; 
        10'b0001001010: data <= 22'h0000d7; 
        10'b0001001011: data <= 22'h3ffb9d; 
        10'b0001001100: data <= 22'h000a8b; 
        10'b0001001101: data <= 22'h3ffd3c; 
        10'b0001001110: data <= 22'h3ffc37; 
        10'b0001001111: data <= 22'h000a7f; 
        10'b0001010000: data <= 22'h0001e3; 
        10'b0001010001: data <= 22'h0001d5; 
        10'b0001010010: data <= 22'h000258; 
        10'b0001010011: data <= 22'h0004ad; 
        10'b0001010100: data <= 22'h000d14; 
        10'b0001010101: data <= 22'h000071; 
        10'b0001010110: data <= 22'h3ffece; 
        10'b0001010111: data <= 22'h0003df; 
        10'b0001011000: data <= 22'h000419; 
        10'b0001011001: data <= 22'h3ffbab; 
        10'b0001011010: data <= 22'h000ab5; 
        10'b0001011011: data <= 22'h0005dc; 
        10'b0001011100: data <= 22'h3ffde4; 
        10'b0001011101: data <= 22'h000ad0; 
        10'b0001011110: data <= 22'h000363; 
        10'b0001011111: data <= 22'h000885; 
        10'b0001100000: data <= 22'h3fff20; 
        10'b0001100001: data <= 22'h3ff642; 
        10'b0001100010: data <= 22'h3fff20; 
        10'b0001100011: data <= 22'h3ff131; 
        10'b0001100100: data <= 22'h3ffe2d; 
        10'b0001100101: data <= 22'h3ff848; 
        10'b0001100110: data <= 22'h000290; 
        10'b0001100111: data <= 22'h00018b; 
        10'b0001101000: data <= 22'h00034e; 
        10'b0001101001: data <= 22'h3fff2d; 
        10'b0001101010: data <= 22'h00087f; 
        10'b0001101011: data <= 22'h3ffeeb; 
        10'b0001101100: data <= 22'h3ffebe; 
        10'b0001101101: data <= 22'h000bb2; 
        10'b0001101110: data <= 22'h000459; 
        10'b0001101111: data <= 22'h00076e; 
        10'b0001110000: data <= 22'h00016f; 
        10'b0001110001: data <= 22'h00026a; 
        10'b0001110010: data <= 22'h000098; 
        10'b0001110011: data <= 22'h3ffd7a; 
        10'b0001110100: data <= 22'h3ffbd8; 
        10'b0001110101: data <= 22'h00078a; 
        10'b0001110110: data <= 22'h000536; 
        10'b0001110111: data <= 22'h3fff0a; 
        10'b0001111000: data <= 22'h3ff95f; 
        10'b0001111001: data <= 22'h000285; 
        10'b0001111010: data <= 22'h3ff50b; 
        10'b0001111011: data <= 22'h3ff093; 
        10'b0001111100: data <= 22'h3fea50; 
        10'b0001111101: data <= 22'h3fd8a6; 
        10'b0001111110: data <= 22'h3fcde9; 
        10'b0001111111: data <= 22'h3fbd0b; 
        10'b0010000000: data <= 22'h3fce84; 
        10'b0010000001: data <= 22'h3fce5f; 
        10'b0010000010: data <= 22'h3fdb17; 
        10'b0010000011: data <= 22'h3fefc6; 
        10'b0010000100: data <= 22'h3ff866; 
        10'b0010000101: data <= 22'h3ffa88; 
        10'b0010000110: data <= 22'h0001d3; 
        10'b0010000111: data <= 22'h000954; 
        10'b0010001000: data <= 22'h00074e; 
        10'b0010001001: data <= 22'h0006c5; 
        10'b0010001010: data <= 22'h00000c; 
        10'b0010001011: data <= 22'h000055; 
        10'b0010001100: data <= 22'h00090b; 
        10'b0010001101: data <= 22'h00066b; 
        10'b0010001110: data <= 22'h000783; 
        10'b0010001111: data <= 22'h0004c2; 
        10'b0010010000: data <= 22'h0005be; 
        10'b0010010001: data <= 22'h3ff8dd; 
        10'b0010010010: data <= 22'h3ff9a8; 
        10'b0010010011: data <= 22'h3ff8f6; 
        10'b0010010100: data <= 22'h3fe947; 
        10'b0010010101: data <= 22'h3fe9bb; 
        10'b0010010110: data <= 22'h3fe7ef; 
        10'b0010010111: data <= 22'h3fe052; 
        10'b0010011000: data <= 22'h3fd84d; 
        10'b0010011001: data <= 22'h3fd10b; 
        10'b0010011010: data <= 22'h3fb852; 
        10'b0010011011: data <= 22'h3fb29a; 
        10'b0010011100: data <= 22'h3f9e2f; 
        10'b0010011101: data <= 22'h3fbf85; 
        10'b0010011110: data <= 22'h3fd75e; 
        10'b0010011111: data <= 22'h3fec4f; 
        10'b0010100000: data <= 22'h3feb3a; 
        10'b0010100001: data <= 22'h3fe4f4; 
        10'b0010100010: data <= 22'h3fe6d3; 
        10'b0010100011: data <= 22'h3fee0c; 
        10'b0010100100: data <= 22'h3ff8d9; 
        10'b0010100101: data <= 22'h3ffcb0; 
        10'b0010100110: data <= 22'h000118; 
        10'b0010100111: data <= 22'h000656; 
        10'b0010101000: data <= 22'h000820; 
        10'b0010101001: data <= 22'h00085c; 
        10'b0010101010: data <= 22'h3ffac2; 
        10'b0010101011: data <= 22'h00086f; 
        10'b0010101100: data <= 22'h00055e; 
        10'b0010101101: data <= 22'h3fe7d1; 
        10'b0010101110: data <= 22'h3fe291; 
        10'b0010101111: data <= 22'h3fdd55; 
        10'b0010110000: data <= 22'h3fd8eb; 
        10'b0010110001: data <= 22'h3fd00e; 
        10'b0010110010: data <= 22'h3fdcc9; 
        10'b0010110011: data <= 22'h3ff4be; 
        10'b0010110100: data <= 22'h0002d4; 
        10'b0010110101: data <= 22'h002b49; 
        10'b0010110110: data <= 22'h004093; 
        10'b0010110111: data <= 22'h00335e; 
        10'b0010111000: data <= 22'h0023fe; 
        10'b0010111001: data <= 22'h001de8; 
        10'b0010111010: data <= 22'h0025ed; 
        10'b0010111011: data <= 22'h3ff99b; 
        10'b0010111100: data <= 22'h3ff6df; 
        10'b0010111101: data <= 22'h3fe326; 
        10'b0010111110: data <= 22'h3fcc4a; 
        10'b0010111111: data <= 22'h3fcfdf; 
        10'b0011000000: data <= 22'h3fe470; 
        10'b0011000001: data <= 22'h3ff296; 
        10'b0011000010: data <= 22'h3ffdf7; 
        10'b0011000011: data <= 22'h000460; 
        10'b0011000100: data <= 22'h000c78; 
        10'b0011000101: data <= 22'h3fff8c; 
        10'b0011000110: data <= 22'h3ffbf2; 
        10'b0011000111: data <= 22'h3ffb82; 
        10'b0011001000: data <= 22'h3fe45c; 
        10'b0011001001: data <= 22'h3fd5f8; 
        10'b0011001010: data <= 22'h3fce83; 
        10'b0011001011: data <= 22'h3fc519; 
        10'b0011001100: data <= 22'h3fc84b; 
        10'b0011001101: data <= 22'h3fec5b; 
        10'b0011001110: data <= 22'h3ffe65; 
        10'b0011001111: data <= 22'h000f44; 
        10'b0011010000: data <= 22'h003aa9; 
        10'b0011010001: data <= 22'h004605; 
        10'b0011010010: data <= 22'h006000; 
        10'b0011010011: data <= 22'h00607e; 
        10'b0011010100: data <= 22'h006464; 
        10'b0011010101: data <= 22'h002d80; 
        10'b0011010110: data <= 22'h002242; 
        10'b0011010111: data <= 22'h0003b4; 
        10'b0011011000: data <= 22'h0008e6; 
        10'b0011011001: data <= 22'h000a13; 
        10'b0011011010: data <= 22'h3fdd6c; 
        10'b0011011011: data <= 22'h3fc20e; 
        10'b0011011100: data <= 22'h3fdb7d; 
        10'b0011011101: data <= 22'h3ff6e0; 
        10'b0011011110: data <= 22'h3ff6a7; 
        10'b0011011111: data <= 22'h000831; 
        10'b0011100000: data <= 22'h000c19; 
        10'b0011100001: data <= 22'h000c2e; 
        10'b0011100010: data <= 22'h00062f; 
        10'b0011100011: data <= 22'h3ffc47; 
        10'b0011100100: data <= 22'h3fe33b; 
        10'b0011100101: data <= 22'h3fd473; 
        10'b0011100110: data <= 22'h3fcd4b; 
        10'b0011100111: data <= 22'h3fb91b; 
        10'b0011101000: data <= 22'h3fed44; 
        10'b0011101001: data <= 22'h3ff753; 
        10'b0011101010: data <= 22'h3ff5f5; 
        10'b0011101011: data <= 22'h3febd3; 
        10'b0011101100: data <= 22'h3ffe75; 
        10'b0011101101: data <= 22'h001c19; 
        10'b0011101110: data <= 22'h005245; 
        10'b0011101111: data <= 22'h002d69; 
        10'b0011110000: data <= 22'h002e3c; 
        10'b0011110001: data <= 22'h000977; 
        10'b0011110010: data <= 22'h0003a6; 
        10'b0011110011: data <= 22'h000273; 
        10'b0011110100: data <= 22'h3ff0cb; 
        10'b0011110101: data <= 22'h0007e5; 
        10'b0011110110: data <= 22'h3fec85; 
        10'b0011110111: data <= 22'h3fce96; 
        10'b0011111000: data <= 22'h3fd641; 
        10'b0011111001: data <= 22'h3febfd; 
        10'b0011111010: data <= 22'h3ff741; 
        10'b0011111011: data <= 22'h000b48; 
        10'b0011111100: data <= 22'h0003ac; 
        10'b0011111101: data <= 22'h000233; 
        10'b0011111110: data <= 22'h0000d2; 
        10'b0011111111: data <= 22'h3feb6c; 
        10'b0100000000: data <= 22'h3fd322; 
        10'b0100000001: data <= 22'h3fdd97; 
        10'b0100000010: data <= 22'h3ff641; 
        10'b0100000011: data <= 22'h3fec47; 
        10'b0100000100: data <= 22'h3ff443; 
        10'b0100000101: data <= 22'h3ffaad; 
        10'b0100000110: data <= 22'h001517; 
        10'b0100000111: data <= 22'h000cb5; 
        10'b0100001000: data <= 22'h0003ba; 
        10'b0100001001: data <= 22'h0021fb; 
        10'b0100001010: data <= 22'h0038e6; 
        10'b0100001011: data <= 22'h0032bb; 
        10'b0100001100: data <= 22'h3ffe07; 
        10'b0100001101: data <= 22'h3ff175; 
        10'b0100001110: data <= 22'h000090; 
        10'b0100001111: data <= 22'h3fe1b5; 
        10'b0100010000: data <= 22'h3ff326; 
        10'b0100010001: data <= 22'h3fe03e; 
        10'b0100010010: data <= 22'h3fddff; 
        10'b0100010011: data <= 22'h3fdbb9; 
        10'b0100010100: data <= 22'h3fe744; 
        10'b0100010101: data <= 22'h3ff531; 
        10'b0100010110: data <= 22'h3ff827; 
        10'b0100010111: data <= 22'h000a05; 
        10'b0100011000: data <= 22'h00022c; 
        10'b0100011001: data <= 22'h3fff90; 
        10'b0100011010: data <= 22'h3ffb2b; 
        10'b0100011011: data <= 22'h3ff81e; 
        10'b0100011100: data <= 22'h3fdd6f; 
        10'b0100011101: data <= 22'h3fedec; 
        10'b0100011110: data <= 22'h0010db; 
        10'b0100011111: data <= 22'h001614; 
        10'b0100100000: data <= 22'h002cce; 
        10'b0100100001: data <= 22'h002c7e; 
        10'b0100100010: data <= 22'h00264f; 
        10'b0100100011: data <= 22'h0039b0; 
        10'b0100100100: data <= 22'h001d0a; 
        10'b0100100101: data <= 22'h0006d7; 
        10'b0100100110: data <= 22'h00076a; 
        10'b0100100111: data <= 22'h3fe2cd; 
        10'b0100101000: data <= 22'h3fee97; 
        10'b0100101001: data <= 22'h3ffc8e; 
        10'b0100101010: data <= 22'h001457; 
        10'b0100101011: data <= 22'h3fff91; 
        10'b0100101100: data <= 22'h00105d; 
        10'b0100101101: data <= 22'h3ff63a; 
        10'b0100101110: data <= 22'h3febec; 
        10'b0100101111: data <= 22'h3fed0d; 
        10'b0100110000: data <= 22'h3fe7f1; 
        10'b0100110001: data <= 22'h3ff921; 
        10'b0100110010: data <= 22'h3ff6e8; 
        10'b0100110011: data <= 22'h0005c0; 
        10'b0100110100: data <= 22'h3ffe1a; 
        10'b0100110101: data <= 22'h00024e; 
        10'b0100110110: data <= 22'h3ffacd; 
        10'b0100110111: data <= 22'h3ffcb2; 
        10'b0100111000: data <= 22'h3ff685; 
        10'b0100111001: data <= 22'h001fcd; 
        10'b0100111010: data <= 22'h004992; 
        10'b0100111011: data <= 22'h0036e9; 
        10'b0100111100: data <= 22'h005646; 
        10'b0100111101: data <= 22'h002296; 
        10'b0100111110: data <= 22'h0023dc; 
        10'b0100111111: data <= 22'h003d9b; 
        10'b0101000000: data <= 22'h3fec67; 
        10'b0101000001: data <= 22'h3fef58; 
        10'b0101000010: data <= 22'h3ff700; 
        10'b0101000011: data <= 22'h00045a; 
        10'b0101000100: data <= 22'h0017cf; 
        10'b0101000101: data <= 22'h005362; 
        10'b0101000110: data <= 22'h002763; 
        10'b0101000111: data <= 22'h0027ed; 
        10'b0101001000: data <= 22'h004179; 
        10'b0101001001: data <= 22'h002f61; 
        10'b0101001010: data <= 22'h001bae; 
        10'b0101001011: data <= 22'h0005b9; 
        10'b0101001100: data <= 22'h3ffb78; 
        10'b0101001101: data <= 22'h3ff4b8; 
        10'b0101001110: data <= 22'h3fff82; 
        10'b0101001111: data <= 22'h00000d; 
        10'b0101010000: data <= 22'h000536; 
        10'b0101010001: data <= 22'h000abb; 
        10'b0101010010: data <= 22'h3ff899; 
        10'b0101010011: data <= 22'h3ff42f; 
        10'b0101010100: data <= 22'h001ad8; 
        10'b0101010101: data <= 22'h0045c2; 
        10'b0101010110: data <= 22'h0050b6; 
        10'b0101010111: data <= 22'h002fe0; 
        10'b0101011000: data <= 22'h003bd6; 
        10'b0101011001: data <= 22'h00492b; 
        10'b0101011010: data <= 22'h002eba; 
        10'b0101011011: data <= 22'h00008c; 
        10'b0101011100: data <= 22'h3fd11f; 
        10'b0101011101: data <= 22'h00289c; 
        10'b0101011110: data <= 22'h0057bd; 
        10'b0101011111: data <= 22'h004569; 
        10'b0101100000: data <= 22'h003b59; 
        10'b0101100001: data <= 22'h005abd; 
        10'b0101100010: data <= 22'h005b64; 
        10'b0101100011: data <= 22'h005ed7; 
        10'b0101100100: data <= 22'h006180; 
        10'b0101100101: data <= 22'h004127; 
        10'b0101100110: data <= 22'h001f56; 
        10'b0101100111: data <= 22'h0000d4; 
        10'b0101101000: data <= 22'h3ff17e; 
        10'b0101101001: data <= 22'h00025e; 
        10'b0101101010: data <= 22'h000543; 
        10'b0101101011: data <= 22'h0005b2; 
        10'b0101101100: data <= 22'h000c10; 
        10'b0101101101: data <= 22'h000768; 
        10'b0101101110: data <= 22'h3ff5da; 
        10'b0101101111: data <= 22'h0003cf; 
        10'b0101110000: data <= 22'h002897; 
        10'b0101110001: data <= 22'h003d0b; 
        10'b0101110010: data <= 22'h003986; 
        10'b0101110011: data <= 22'h0025c3; 
        10'b0101110100: data <= 22'h002f6a; 
        10'b0101110101: data <= 22'h001e70; 
        10'b0101110110: data <= 22'h001b81; 
        10'b0101110111: data <= 22'h3ff1c1; 
        10'b0101111000: data <= 22'h3fe762; 
        10'b0101111001: data <= 22'h003fd4; 
        10'b0101111010: data <= 22'h00578d; 
        10'b0101111011: data <= 22'h003f70; 
        10'b0101111100: data <= 22'h00491c; 
        10'b0101111101: data <= 22'h00418b; 
        10'b0101111110: data <= 22'h0059ea; 
        10'b0101111111: data <= 22'h005b7a; 
        10'b0110000000: data <= 22'h004780; 
        10'b0110000001: data <= 22'h0029c3; 
        10'b0110000010: data <= 22'h000264; 
        10'b0110000011: data <= 22'h3fe38f; 
        10'b0110000100: data <= 22'h3fef6e; 
        10'b0110000101: data <= 22'h3ffada; 
        10'b0110000110: data <= 22'h000565; 
        10'b0110000111: data <= 22'h00057b; 
        10'b0110001000: data <= 22'h00026d; 
        10'b0110001001: data <= 22'h000133; 
        10'b0110001010: data <= 22'h00084c; 
        10'b0110001011: data <= 22'h000546; 
        10'b0110001100: data <= 22'h001292; 
        10'b0110001101: data <= 22'h001181; 
        10'b0110001110: data <= 22'h002faa; 
        10'b0110001111: data <= 22'h002159; 
        10'b0110010000: data <= 22'h001036; 
        10'b0110010001: data <= 22'h3fffd3; 
        10'b0110010010: data <= 22'h0005ef; 
        10'b0110010011: data <= 22'h3ffd0b; 
        10'b0110010100: data <= 22'h3fee02; 
        10'b0110010101: data <= 22'h0014b2; 
        10'b0110010110: data <= 22'h000bc1; 
        10'b0110010111: data <= 22'h0037fc; 
        10'b0110011000: data <= 22'h003b61; 
        10'b0110011001: data <= 22'h003b76; 
        10'b0110011010: data <= 22'h00287f; 
        10'b0110011011: data <= 22'h001a07; 
        10'b0110011100: data <= 22'h00207a; 
        10'b0110011101: data <= 22'h000098; 
        10'b0110011110: data <= 22'h3fdf37; 
        10'b0110011111: data <= 22'h3fd05d; 
        10'b0110100000: data <= 22'h3fec4b; 
        10'b0110100001: data <= 22'h00034a; 
        10'b0110100010: data <= 22'h0001e0; 
        10'b0110100011: data <= 22'h000238; 
        10'b0110100100: data <= 22'h000921; 
        10'b0110100101: data <= 22'h000853; 
        10'b0110100110: data <= 22'h000583; 
        10'b0110100111: data <= 22'h3ff958; 
        10'b0110101000: data <= 22'h00015c; 
        10'b0110101001: data <= 22'h001533; 
        10'b0110101010: data <= 22'h00144e; 
        10'b0110101011: data <= 22'h000d69; 
        10'b0110101100: data <= 22'h000dad; 
        10'b0110101101: data <= 22'h3fe6df; 
        10'b0110101110: data <= 22'h3ff454; 
        10'b0110101111: data <= 22'h3ff43f; 
        10'b0110110000: data <= 22'h3fee75; 
        10'b0110110001: data <= 22'h3ff26d; 
        10'b0110110010: data <= 22'h3fef8c; 
        10'b0110110011: data <= 22'h003d29; 
        10'b0110110100: data <= 22'h00598a; 
        10'b0110110101: data <= 22'h0055d2; 
        10'b0110110110: data <= 22'h002af8; 
        10'b0110110111: data <= 22'h000426; 
        10'b0110111000: data <= 22'h3fed56; 
        10'b0110111001: data <= 22'h3fcec9; 
        10'b0110111010: data <= 22'h3fc29c; 
        10'b0110111011: data <= 22'h3fd426; 
        10'b0110111100: data <= 22'h3fec7c; 
        10'b0110111101: data <= 22'h00005c; 
        10'b0110111110: data <= 22'h000504; 
        10'b0110111111: data <= 22'h3fff4a; 
        10'b0111000000: data <= 22'h000a82; 
        10'b0111000001: data <= 22'h0000e1; 
        10'b0111000010: data <= 22'h3ff879; 
        10'b0111000011: data <= 22'h3ffe11; 
        10'b0111000100: data <= 22'h0000ab; 
        10'b0111000101: data <= 22'h00065b; 
        10'b0111000110: data <= 22'h3fef98; 
        10'b0111000111: data <= 22'h000cf5; 
        10'b0111001000: data <= 22'h0024cf; 
        10'b0111001001: data <= 22'h3ff760; 
        10'b0111001010: data <= 22'h0014e2; 
        10'b0111001011: data <= 22'h001d9b; 
        10'b0111001100: data <= 22'h3ffbf7; 
        10'b0111001101: data <= 22'h3fde51; 
        10'b0111001110: data <= 22'h3ffa5d; 
        10'b0111001111: data <= 22'h0021f4; 
        10'b0111010000: data <= 22'h003d19; 
        10'b0111010001: data <= 22'h003cb4; 
        10'b0111010010: data <= 22'h000f29; 
        10'b0111010011: data <= 22'h3fdd7b; 
        10'b0111010100: data <= 22'h3fc6b6; 
        10'b0111010101: data <= 22'h3fb0cb; 
        10'b0111010110: data <= 22'h3fc864; 
        10'b0111010111: data <= 22'h3fd2d1; 
        10'b0111011000: data <= 22'h3fe21a; 
        10'b0111011001: data <= 22'h0000fd; 
        10'b0111011010: data <= 22'h3ff979; 
        10'b0111011011: data <= 22'h0005a6; 
        10'b0111011100: data <= 22'h000378; 
        10'b0111011101: data <= 22'h3ffdaf; 
        10'b0111011110: data <= 22'h3ff7c7; 
        10'b0111011111: data <= 22'h3ff3fb; 
        10'b0111100000: data <= 22'h3fe97e; 
        10'b0111100001: data <= 22'h3fe49d; 
        10'b0111100010: data <= 22'h3fe96d; 
        10'b0111100011: data <= 22'h000a2e; 
        10'b0111100100: data <= 22'h0013d3; 
        10'b0111100101: data <= 22'h001694; 
        10'b0111100110: data <= 22'h00226d; 
        10'b0111100111: data <= 22'h003218; 
        10'b0111101000: data <= 22'h001e8d; 
        10'b0111101001: data <= 22'h000e33; 
        10'b0111101010: data <= 22'h001368; 
        10'b0111101011: data <= 22'h0031d4; 
        10'b0111101100: data <= 22'h000ecc; 
        10'b0111101101: data <= 22'h3ff5e7; 
        10'b0111101110: data <= 22'h3fe9fb; 
        10'b0111101111: data <= 22'h3fcd68; 
        10'b0111110000: data <= 22'h3fce0e; 
        10'b0111110001: data <= 22'h3fca3c; 
        10'b0111110010: data <= 22'h3fcd6f; 
        10'b0111110011: data <= 22'h3fdac6; 
        10'b0111110100: data <= 22'h3fe4e4; 
        10'b0111110101: data <= 22'h0002b5; 
        10'b0111110110: data <= 22'h0002cb; 
        10'b0111110111: data <= 22'h3ffd9d; 
        10'b0111111000: data <= 22'h0009b4; 
        10'b0111111001: data <= 22'h3ffff8; 
        10'b0111111010: data <= 22'h3ffa56; 
        10'b0111111011: data <= 22'h3ffdbf; 
        10'b0111111100: data <= 22'h3fec35; 
        10'b0111111101: data <= 22'h3fd28f; 
        10'b0111111110: data <= 22'h3fd1ad; 
        10'b0111111111: data <= 22'h3fd28e; 
        10'b1000000000: data <= 22'h3fece9; 
        10'b1000000001: data <= 22'h000793; 
        10'b1000000010: data <= 22'h0036e4; 
        10'b1000000011: data <= 22'h002c5e; 
        10'b1000000100: data <= 22'h3fe4eb; 
        10'b1000000101: data <= 22'h3fe483; 
        10'b1000000110: data <= 22'h0001b3; 
        10'b1000000111: data <= 22'h0020fc; 
        10'b1000001000: data <= 22'h3febc8; 
        10'b1000001001: data <= 22'h3fe8f0; 
        10'b1000001010: data <= 22'h3fd4d1; 
        10'b1000001011: data <= 22'h3fe603; 
        10'b1000001100: data <= 22'h3fe7a2; 
        10'b1000001101: data <= 22'h3fd9f7; 
        10'b1000001110: data <= 22'h3fd7f9; 
        10'b1000001111: data <= 22'h3fd617; 
        10'b1000010000: data <= 22'h3fe25a; 
        10'b1000010001: data <= 22'h3ffb49; 
        10'b1000010010: data <= 22'h000099; 
        10'b1000010011: data <= 22'h0008df; 
        10'b1000010100: data <= 22'h00064b; 
        10'b1000010101: data <= 22'h000c93; 
        10'b1000010110: data <= 22'h00023b; 
        10'b1000010111: data <= 22'h3ff521; 
        10'b1000011000: data <= 22'h3fedd5; 
        10'b1000011001: data <= 22'h3fdfd7; 
        10'b1000011010: data <= 22'h3fcd2c; 
        10'b1000011011: data <= 22'h3fcbd6; 
        10'b1000011100: data <= 22'h3fc9fd; 
        10'b1000011101: data <= 22'h3fca6c; 
        10'b1000011110: data <= 22'h3fc409; 
        10'b1000011111: data <= 22'h3fcd59; 
        10'b1000100000: data <= 22'h3fbe6e; 
        10'b1000100001: data <= 22'h3fd22b; 
        10'b1000100010: data <= 22'h3fd95f; 
        10'b1000100011: data <= 22'h3fd40e; 
        10'b1000100100: data <= 22'h3fda13; 
        10'b1000100101: data <= 22'h3ff39c; 
        10'b1000100110: data <= 22'h3fe324; 
        10'b1000100111: data <= 22'h3ff7f1; 
        10'b1000101000: data <= 22'h3fecb3; 
        10'b1000101001: data <= 22'h3fe921; 
        10'b1000101010: data <= 22'h3fea69; 
        10'b1000101011: data <= 22'h3feccc; 
        10'b1000101100: data <= 22'h3ff3ec; 
        10'b1000101101: data <= 22'h000379; 
        10'b1000101110: data <= 22'h3ffc33; 
        10'b1000101111: data <= 22'h000159; 
        10'b1000110000: data <= 22'h3ffda2; 
        10'b1000110001: data <= 22'h0001c1; 
        10'b1000110010: data <= 22'h000557; 
        10'b1000110011: data <= 22'h000068; 
        10'b1000110100: data <= 22'h3fed31; 
        10'b1000110101: data <= 22'h3fe0f2; 
        10'b1000110110: data <= 22'h3fd0e9; 
        10'b1000110111: data <= 22'h3fb63d; 
        10'b1000111000: data <= 22'h3fab85; 
        10'b1000111001: data <= 22'h3fa13b; 
        10'b1000111010: data <= 22'h3f7fb4; 
        10'b1000111011: data <= 22'h3f9dcf; 
        10'b1000111100: data <= 22'h3fa052; 
        10'b1000111101: data <= 22'h3fe0b1; 
        10'b1000111110: data <= 22'h3fd417; 
        10'b1000111111: data <= 22'h3feb60; 
        10'b1001000000: data <= 22'h3fe744; 
        10'b1001000001: data <= 22'h3ff956; 
        10'b1001000010: data <= 22'h3fd5f3; 
        10'b1001000011: data <= 22'h3ff227; 
        10'b1001000100: data <= 22'h3fef4f; 
        10'b1001000101: data <= 22'h3fe533; 
        10'b1001000110: data <= 22'h3ff872; 
        10'b1001000111: data <= 22'h3ff329; 
        10'b1001001000: data <= 22'h00014b; 
        10'b1001001001: data <= 22'h000ab4; 
        10'b1001001010: data <= 22'h000674; 
        10'b1001001011: data <= 22'h000206; 
        10'b1001001100: data <= 22'h0000dc; 
        10'b1001001101: data <= 22'h000002; 
        10'b1001001110: data <= 22'h000ab4; 
        10'b1001001111: data <= 22'h3ff4a8; 
        10'b1001010000: data <= 22'h3ff358; 
        10'b1001010001: data <= 22'h3fe161; 
        10'b1001010010: data <= 22'h3fd4c1; 
        10'b1001010011: data <= 22'h3fbd41; 
        10'b1001010100: data <= 22'h3fb43a; 
        10'b1001010101: data <= 22'h3faca4; 
        10'b1001010110: data <= 22'h3fa89e; 
        10'b1001010111: data <= 22'h3fb16a; 
        10'b1001011000: data <= 22'h3fcdef; 
        10'b1001011001: data <= 22'h3fce96; 
        10'b1001011010: data <= 22'h3fcdc5; 
        10'b1001011011: data <= 22'h3fe32e; 
        10'b1001011100: data <= 22'h3fe0c8; 
        10'b1001011101: data <= 22'h3fd102; 
        10'b1001011110: data <= 22'h3fc74c; 
        10'b1001011111: data <= 22'h3fe7f9; 
        10'b1001100000: data <= 22'h3ff299; 
        10'b1001100001: data <= 22'h3ff846; 
        10'b1001100010: data <= 22'h0003c9; 
        10'b1001100011: data <= 22'h3ffeee; 
        10'b1001100100: data <= 22'h0004cf; 
        10'b1001100101: data <= 22'h000693; 
        10'b1001100110: data <= 22'h00005f; 
        10'b1001100111: data <= 22'h0000c9; 
        10'b1001101000: data <= 22'h000836; 
        10'b1001101001: data <= 22'h00020d; 
        10'b1001101010: data <= 22'h000251; 
        10'b1001101011: data <= 22'h0007dc; 
        10'b1001101100: data <= 22'h3ffaf3; 
        10'b1001101101: data <= 22'h3fe744; 
        10'b1001101110: data <= 22'h3fd86d; 
        10'b1001101111: data <= 22'h3fca2b; 
        10'b1001110000: data <= 22'h3fd7f0; 
        10'b1001110001: data <= 22'h3fd625; 
        10'b1001110010: data <= 22'h3fd24c; 
        10'b1001110011: data <= 22'h3fe124; 
        10'b1001110100: data <= 22'h3fdd4f; 
        10'b1001110101: data <= 22'h3fd1d7; 
        10'b1001110110: data <= 22'h3fd935; 
        10'b1001110111: data <= 22'h3fc9a0; 
        10'b1001111000: data <= 22'h3fc3db; 
        10'b1001111001: data <= 22'h3fc50a; 
        10'b1001111010: data <= 22'h3fcef7; 
        10'b1001111011: data <= 22'h3fd467; 
        10'b1001111100: data <= 22'h3ff408; 
        10'b1001111101: data <= 22'h000eac; 
        10'b1001111110: data <= 22'h000828; 
        10'b1001111111: data <= 22'h000a1f; 
        10'b1010000000: data <= 22'h00108b; 
        10'b1010000001: data <= 22'h000378; 
        10'b1010000010: data <= 22'h0003dc; 
        10'b1010000011: data <= 22'h000609; 
        10'b1010000100: data <= 22'h0009a3; 
        10'b1010000101: data <= 22'h000790; 
        10'b1010000110: data <= 22'h0002d5; 
        10'b1010000111: data <= 22'h3ffc39; 
        10'b1010001000: data <= 22'h3ff90f; 
        10'b1010001001: data <= 22'h3feabb; 
        10'b1010001010: data <= 22'h3fe745; 
        10'b1010001011: data <= 22'h3fdf4d; 
        10'b1010001100: data <= 22'h3ffd88; 
        10'b1010001101: data <= 22'h3ff2c7; 
        10'b1010001110: data <= 22'h3ff568; 
        10'b1010001111: data <= 22'h3fd85f; 
        10'b1010010000: data <= 22'h3fdfb5; 
        10'b1010010001: data <= 22'h3fd742; 
        10'b1010010010: data <= 22'h3fdd8e; 
        10'b1010010011: data <= 22'h3fc530; 
        10'b1010010100: data <= 22'h3fc084; 
        10'b1010010101: data <= 22'h3fc81f; 
        10'b1010010110: data <= 22'h3fdd2f; 
        10'b1010010111: data <= 22'h3ffc9b; 
        10'b1010011000: data <= 22'h000da2; 
        10'b1010011001: data <= 22'h001fa3; 
        10'b1010011010: data <= 22'h002d9a; 
        10'b1010011011: data <= 22'h002632; 
        10'b1010011100: data <= 22'h0011e0; 
        10'b1010011101: data <= 22'h3ffec7; 
        10'b1010011110: data <= 22'h000cd1; 
        10'b1010011111: data <= 22'h3ffe82; 
        10'b1010100000: data <= 22'h3ffff5; 
        10'b1010100001: data <= 22'h3ffaf2; 
        10'b1010100010: data <= 22'h3ffea5; 
        10'b1010100011: data <= 22'h000acc; 
        10'b1010100100: data <= 22'h0007c3; 
        10'b1010100101: data <= 22'h000c29; 
        10'b1010100110: data <= 22'h0008d6; 
        10'b1010100111: data <= 22'h000cd5; 
        10'b1010101000: data <= 22'h001222; 
        10'b1010101001: data <= 22'h0009ca; 
        10'b1010101010: data <= 22'h3ff98b; 
        10'b1010101011: data <= 22'h3febad; 
        10'b1010101100: data <= 22'h3ffe90; 
        10'b1010101101: data <= 22'h3fe0cf; 
        10'b1010101110: data <= 22'h3fd893; 
        10'b1010101111: data <= 22'h3fd660; 
        10'b1010110000: data <= 22'h3fed20; 
        10'b1010110001: data <= 22'h000db2; 
        10'b1010110010: data <= 22'h001760; 
        10'b1010110011: data <= 22'h001829; 
        10'b1010110100: data <= 22'h00372b; 
        10'b1010110101: data <= 22'h003b5f; 
        10'b1010110110: data <= 22'h00222d; 
        10'b1010110111: data <= 22'h0014e3; 
        10'b1010111000: data <= 22'h00107e; 
        10'b1010111001: data <= 22'h3ffcc4; 
        10'b1010111010: data <= 22'h00075f; 
        10'b1010111011: data <= 22'h3fff83; 
        10'b1010111100: data <= 22'h0002b0; 
        10'b1010111101: data <= 22'h000ab5; 
        10'b1010111110: data <= 22'h000abd; 
        10'b1010111111: data <= 22'h3ffede; 
        10'b1011000000: data <= 22'h000102; 
        10'b1011000001: data <= 22'h001255; 
        10'b1011000010: data <= 22'h000de3; 
        10'b1011000011: data <= 22'h002814; 
        10'b1011000100: data <= 22'h002bed; 
        10'b1011000101: data <= 22'h002cb8; 
        10'b1011000110: data <= 22'h0026b1; 
        10'b1011000111: data <= 22'h000f5d; 
        10'b1011001000: data <= 22'h0028b3; 
        10'b1011001001: data <= 22'h00244e; 
        10'b1011001010: data <= 22'h0022c2; 
        10'b1011001011: data <= 22'h0020ac; 
        10'b1011001100: data <= 22'h003d09; 
        10'b1011001101: data <= 22'h004254; 
        10'b1011001110: data <= 22'h0048f3; 
        10'b1011001111: data <= 22'h004c24; 
        10'b1011010000: data <= 22'h0054fe; 
        10'b1011010001: data <= 22'h003c4f; 
        10'b1011010010: data <= 22'h001788; 
        10'b1011010011: data <= 22'h000b28; 
        10'b1011010100: data <= 22'h3ffe81; 
        10'b1011010101: data <= 22'h3fff1a; 
        10'b1011010110: data <= 22'h000320; 
        10'b1011010111: data <= 22'h0002a0; 
        10'b1011011000: data <= 22'h000074; 
        10'b1011011001: data <= 22'h0009c1; 
        10'b1011011010: data <= 22'h00029e; 
        10'b1011011011: data <= 22'h3ffc72; 
        10'b1011011100: data <= 22'h0009d0; 
        10'b1011011101: data <= 22'h000f33; 
        10'b1011011110: data <= 22'h001553; 
        10'b1011011111: data <= 22'h001d9e; 
        10'b1011100000: data <= 22'h0021b8; 
        10'b1011100001: data <= 22'h003323; 
        10'b1011100010: data <= 22'h0034c4; 
        10'b1011100011: data <= 22'h003b45; 
        10'b1011100100: data <= 22'h00462f; 
        10'b1011100101: data <= 22'h0046ce; 
        10'b1011100110: data <= 22'h0056b2; 
        10'b1011100111: data <= 22'h003203; 
        10'b1011101000: data <= 22'h002241; 
        10'b1011101001: data <= 22'h001cee; 
        10'b1011101010: data <= 22'h002aaa; 
        10'b1011101011: data <= 22'h002e0e; 
        10'b1011101100: data <= 22'h00216f; 
        10'b1011101101: data <= 22'h00174a; 
        10'b1011101110: data <= 22'h0009b0; 
        10'b1011101111: data <= 22'h00037e; 
        10'b1011110000: data <= 22'h00022d; 
        10'b1011110001: data <= 22'h0003dc; 
        10'b1011110010: data <= 22'h3ffc57; 
        10'b1011110011: data <= 22'h000222; 
        10'b1011110100: data <= 22'h3ffda9; 
        10'b1011110101: data <= 22'h000476; 
        10'b1011110110: data <= 22'h3ffbfa; 
        10'b1011110111: data <= 22'h000bd2; 
        10'b1011111000: data <= 22'h0006c9; 
        10'b1011111001: data <= 22'h0003c0; 
        10'b1011111010: data <= 22'h3ffe53; 
        10'b1011111011: data <= 22'h000b7d; 
        10'b1011111100: data <= 22'h0009b6; 
        10'b1011111101: data <= 22'h0006a4; 
        10'b1011111110: data <= 22'h3ffddc; 
        10'b1011111111: data <= 22'h3ffd9a; 
        10'b1100000000: data <= 22'h000248; 
        10'b1100000001: data <= 22'h3ffdde; 
        10'b1100000010: data <= 22'h00027a; 
        10'b1100000011: data <= 22'h000760; 
        10'b1100000100: data <= 22'h0000ae; 
        10'b1100000101: data <= 22'h000406; 
        10'b1100000110: data <= 22'h000d1e; 
        10'b1100000111: data <= 22'h000baf; 
        10'b1100001000: data <= 22'h000695; 
        10'b1100001001: data <= 22'h000405; 
        10'b1100001010: data <= 22'h3ffcbe; 
        10'b1100001011: data <= 22'h000cf7; 
        10'b1100001100: data <= 22'h00070b; 
        10'b1100001101: data <= 22'h3ffd9b; 
        10'b1100001110: data <= 22'h0000e6; 
        10'b1100001111: data <= 22'h3ffeb1; 
      endcase 
    end 
  end 
endgenerate 
assign dout = data; 
endmodule
