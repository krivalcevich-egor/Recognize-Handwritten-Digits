`timescale 1ns / 1ps 
 
////////////////////////////////////////////////////////////////////////////////// 
// WEIGHT MEMORY (ROM) 
////////////////////////////////////////////////////////////////////////////////// 
module ROM_weights_1 #( 
    parameter int WGHT_INT = 6, // integer part 
    parameter int WGHT_FRC = 16 // fractional part 
)( 
    input logic clk, // clock 
    input logic [9:0] address,
    output [WGHT_INT + WGHT_FRC-1:0] dout 
); 

(* rom_style = "block" *) reg [WGHT_INT + WGHT_FRC-1:0] data;
generate 
  if (WGHT_FRC == 1) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 7'h00; 
        10'b0000000001: data <= 7'h00; 
        10'b0000000010: data <= 7'h00; 
        10'b0000000011: data <= 7'h00; 
        10'b0000000100: data <= 7'h00; 
        10'b0000000101: data <= 7'h00; 
        10'b0000000110: data <= 7'h00; 
        10'b0000000111: data <= 7'h00; 
        10'b0000001000: data <= 7'h00; 
        10'b0000001001: data <= 7'h00; 
        10'b0000001010: data <= 7'h00; 
        10'b0000001011: data <= 7'h00; 
        10'b0000001100: data <= 7'h00; 
        10'b0000001101: data <= 7'h00; 
        10'b0000001110: data <= 7'h00; 
        10'b0000001111: data <= 7'h00; 
        10'b0000010000: data <= 7'h00; 
        10'b0000010001: data <= 7'h00; 
        10'b0000010010: data <= 7'h00; 
        10'b0000010011: data <= 7'h00; 
        10'b0000010100: data <= 7'h00; 
        10'b0000010101: data <= 7'h00; 
        10'b0000010110: data <= 7'h00; 
        10'b0000010111: data <= 7'h00; 
        10'b0000011000: data <= 7'h00; 
        10'b0000011001: data <= 7'h00; 
        10'b0000011010: data <= 7'h00; 
        10'b0000011011: data <= 7'h00; 
        10'b0000011100: data <= 7'h00; 
        10'b0000011101: data <= 7'h00; 
        10'b0000011110: data <= 7'h00; 
        10'b0000011111: data <= 7'h00; 
        10'b0000100000: data <= 7'h00; 
        10'b0000100001: data <= 7'h00; 
        10'b0000100010: data <= 7'h00; 
        10'b0000100011: data <= 7'h00; 
        10'b0000100100: data <= 7'h00; 
        10'b0000100101: data <= 7'h00; 
        10'b0000100110: data <= 7'h00; 
        10'b0000100111: data <= 7'h00; 
        10'b0000101000: data <= 7'h00; 
        10'b0000101001: data <= 7'h00; 
        10'b0000101010: data <= 7'h00; 
        10'b0000101011: data <= 7'h00; 
        10'b0000101100: data <= 7'h00; 
        10'b0000101101: data <= 7'h00; 
        10'b0000101110: data <= 7'h00; 
        10'b0000101111: data <= 7'h00; 
        10'b0000110000: data <= 7'h00; 
        10'b0000110001: data <= 7'h00; 
        10'b0000110010: data <= 7'h00; 
        10'b0000110011: data <= 7'h00; 
        10'b0000110100: data <= 7'h00; 
        10'b0000110101: data <= 7'h00; 
        10'b0000110110: data <= 7'h00; 
        10'b0000110111: data <= 7'h00; 
        10'b0000111000: data <= 7'h00; 
        10'b0000111001: data <= 7'h00; 
        10'b0000111010: data <= 7'h00; 
        10'b0000111011: data <= 7'h00; 
        10'b0000111100: data <= 7'h00; 
        10'b0000111101: data <= 7'h00; 
        10'b0000111110: data <= 7'h00; 
        10'b0000111111: data <= 7'h00; 
        10'b0001000000: data <= 7'h00; 
        10'b0001000001: data <= 7'h00; 
        10'b0001000010: data <= 7'h00; 
        10'b0001000011: data <= 7'h00; 
        10'b0001000100: data <= 7'h00; 
        10'b0001000101: data <= 7'h00; 
        10'b0001000110: data <= 7'h00; 
        10'b0001000111: data <= 7'h00; 
        10'b0001001000: data <= 7'h00; 
        10'b0001001001: data <= 7'h00; 
        10'b0001001010: data <= 7'h00; 
        10'b0001001011: data <= 7'h00; 
        10'b0001001100: data <= 7'h00; 
        10'b0001001101: data <= 7'h00; 
        10'b0001001110: data <= 7'h00; 
        10'b0001001111: data <= 7'h00; 
        10'b0001010000: data <= 7'h00; 
        10'b0001010001: data <= 7'h00; 
        10'b0001010010: data <= 7'h00; 
        10'b0001010011: data <= 7'h00; 
        10'b0001010100: data <= 7'h00; 
        10'b0001010101: data <= 7'h00; 
        10'b0001010110: data <= 7'h00; 
        10'b0001010111: data <= 7'h00; 
        10'b0001011000: data <= 7'h00; 
        10'b0001011001: data <= 7'h00; 
        10'b0001011010: data <= 7'h00; 
        10'b0001011011: data <= 7'h00; 
        10'b0001011100: data <= 7'h00; 
        10'b0001011101: data <= 7'h00; 
        10'b0001011110: data <= 7'h00; 
        10'b0001011111: data <= 7'h00; 
        10'b0001100000: data <= 7'h00; 
        10'b0001100001: data <= 7'h00; 
        10'b0001100010: data <= 7'h00; 
        10'b0001100011: data <= 7'h00; 
        10'b0001100100: data <= 7'h00; 
        10'b0001100101: data <= 7'h00; 
        10'b0001100110: data <= 7'h00; 
        10'b0001100111: data <= 7'h00; 
        10'b0001101000: data <= 7'h00; 
        10'b0001101001: data <= 7'h00; 
        10'b0001101010: data <= 7'h00; 
        10'b0001101011: data <= 7'h00; 
        10'b0001101100: data <= 7'h00; 
        10'b0001101101: data <= 7'h00; 
        10'b0001101110: data <= 7'h00; 
        10'b0001101111: data <= 7'h00; 
        10'b0001110000: data <= 7'h00; 
        10'b0001110001: data <= 7'h00; 
        10'b0001110010: data <= 7'h00; 
        10'b0001110011: data <= 7'h00; 
        10'b0001110100: data <= 7'h00; 
        10'b0001110101: data <= 7'h00; 
        10'b0001110110: data <= 7'h00; 
        10'b0001110111: data <= 7'h00; 
        10'b0001111000: data <= 7'h00; 
        10'b0001111001: data <= 7'h00; 
        10'b0001111010: data <= 7'h00; 
        10'b0001111011: data <= 7'h00; 
        10'b0001111100: data <= 7'h00; 
        10'b0001111101: data <= 7'h00; 
        10'b0001111110: data <= 7'h00; 
        10'b0001111111: data <= 7'h00; 
        10'b0010000000: data <= 7'h00; 
        10'b0010000001: data <= 7'h00; 
        10'b0010000010: data <= 7'h00; 
        10'b0010000011: data <= 7'h00; 
        10'b0010000100: data <= 7'h00; 
        10'b0010000101: data <= 7'h00; 
        10'b0010000110: data <= 7'h00; 
        10'b0010000111: data <= 7'h00; 
        10'b0010001000: data <= 7'h00; 
        10'b0010001001: data <= 7'h00; 
        10'b0010001010: data <= 7'h00; 
        10'b0010001011: data <= 7'h00; 
        10'b0010001100: data <= 7'h00; 
        10'b0010001101: data <= 7'h00; 
        10'b0010001110: data <= 7'h00; 
        10'b0010001111: data <= 7'h00; 
        10'b0010010000: data <= 7'h00; 
        10'b0010010001: data <= 7'h00; 
        10'b0010010010: data <= 7'h00; 
        10'b0010010011: data <= 7'h00; 
        10'b0010010100: data <= 7'h00; 
        10'b0010010101: data <= 7'h00; 
        10'b0010010110: data <= 7'h00; 
        10'b0010010111: data <= 7'h00; 
        10'b0010011000: data <= 7'h00; 
        10'b0010011001: data <= 7'h00; 
        10'b0010011010: data <= 7'h00; 
        10'b0010011011: data <= 7'h00; 
        10'b0010011100: data <= 7'h00; 
        10'b0010011101: data <= 7'h00; 
        10'b0010011110: data <= 7'h00; 
        10'b0010011111: data <= 7'h00; 
        10'b0010100000: data <= 7'h00; 
        10'b0010100001: data <= 7'h00; 
        10'b0010100010: data <= 7'h00; 
        10'b0010100011: data <= 7'h00; 
        10'b0010100100: data <= 7'h00; 
        10'b0010100101: data <= 7'h00; 
        10'b0010100110: data <= 7'h00; 
        10'b0010100111: data <= 7'h00; 
        10'b0010101000: data <= 7'h00; 
        10'b0010101001: data <= 7'h00; 
        10'b0010101010: data <= 7'h00; 
        10'b0010101011: data <= 7'h00; 
        10'b0010101100: data <= 7'h00; 
        10'b0010101101: data <= 7'h00; 
        10'b0010101110: data <= 7'h00; 
        10'b0010101111: data <= 7'h00; 
        10'b0010110000: data <= 7'h00; 
        10'b0010110001: data <= 7'h00; 
        10'b0010110010: data <= 7'h00; 
        10'b0010110011: data <= 7'h00; 
        10'b0010110100: data <= 7'h00; 
        10'b0010110101: data <= 7'h00; 
        10'b0010110110: data <= 7'h00; 
        10'b0010110111: data <= 7'h00; 
        10'b0010111000: data <= 7'h00; 
        10'b0010111001: data <= 7'h00; 
        10'b0010111010: data <= 7'h00; 
        10'b0010111011: data <= 7'h00; 
        10'b0010111100: data <= 7'h00; 
        10'b0010111101: data <= 7'h00; 
        10'b0010111110: data <= 7'h00; 
        10'b0010111111: data <= 7'h00; 
        10'b0011000000: data <= 7'h00; 
        10'b0011000001: data <= 7'h00; 
        10'b0011000010: data <= 7'h00; 
        10'b0011000011: data <= 7'h00; 
        10'b0011000100: data <= 7'h00; 
        10'b0011000101: data <= 7'h00; 
        10'b0011000110: data <= 7'h00; 
        10'b0011000111: data <= 7'h00; 
        10'b0011001000: data <= 7'h00; 
        10'b0011001001: data <= 7'h00; 
        10'b0011001010: data <= 7'h00; 
        10'b0011001011: data <= 7'h00; 
        10'b0011001100: data <= 7'h00; 
        10'b0011001101: data <= 7'h7f; 
        10'b0011001110: data <= 7'h00; 
        10'b0011001111: data <= 7'h00; 
        10'b0011010000: data <= 7'h00; 
        10'b0011010001: data <= 7'h00; 
        10'b0011010010: data <= 7'h00; 
        10'b0011010011: data <= 7'h00; 
        10'b0011010100: data <= 7'h00; 
        10'b0011010101: data <= 7'h00; 
        10'b0011010110: data <= 7'h00; 
        10'b0011010111: data <= 7'h00; 
        10'b0011011000: data <= 7'h00; 
        10'b0011011001: data <= 7'h00; 
        10'b0011011010: data <= 7'h00; 
        10'b0011011011: data <= 7'h00; 
        10'b0011011100: data <= 7'h00; 
        10'b0011011101: data <= 7'h00; 
        10'b0011011110: data <= 7'h00; 
        10'b0011011111: data <= 7'h00; 
        10'b0011100000: data <= 7'h00; 
        10'b0011100001: data <= 7'h00; 
        10'b0011100010: data <= 7'h00; 
        10'b0011100011: data <= 7'h00; 
        10'b0011100100: data <= 7'h00; 
        10'b0011100101: data <= 7'h00; 
        10'b0011100110: data <= 7'h00; 
        10'b0011100111: data <= 7'h00; 
        10'b0011101000: data <= 7'h7f; 
        10'b0011101001: data <= 7'h7f; 
        10'b0011101010: data <= 7'h7f; 
        10'b0011101011: data <= 7'h00; 
        10'b0011101100: data <= 7'h00; 
        10'b0011101101: data <= 7'h00; 
        10'b0011101110: data <= 7'h00; 
        10'b0011101111: data <= 7'h00; 
        10'b0011110000: data <= 7'h00; 
        10'b0011110001: data <= 7'h00; 
        10'b0011110010: data <= 7'h00; 
        10'b0011110011: data <= 7'h00; 
        10'b0011110100: data <= 7'h00; 
        10'b0011110101: data <= 7'h00; 
        10'b0011110110: data <= 7'h00; 
        10'b0011110111: data <= 7'h00; 
        10'b0011111000: data <= 7'h00; 
        10'b0011111001: data <= 7'h00; 
        10'b0011111010: data <= 7'h00; 
        10'b0011111011: data <= 7'h00; 
        10'b0011111100: data <= 7'h00; 
        10'b0011111101: data <= 7'h00; 
        10'b0011111110: data <= 7'h00; 
        10'b0011111111: data <= 7'h00; 
        10'b0100000000: data <= 7'h00; 
        10'b0100000001: data <= 7'h00; 
        10'b0100000010: data <= 7'h00; 
        10'b0100000011: data <= 7'h00; 
        10'b0100000100: data <= 7'h00; 
        10'b0100000101: data <= 7'h7f; 
        10'b0100000110: data <= 7'h7f; 
        10'b0100000111: data <= 7'h00; 
        10'b0100001000: data <= 7'h00; 
        10'b0100001001: data <= 7'h00; 
        10'b0100001010: data <= 7'h00; 
        10'b0100001011: data <= 7'h01; 
        10'b0100001100: data <= 7'h00; 
        10'b0100001101: data <= 7'h00; 
        10'b0100001110: data <= 7'h00; 
        10'b0100001111: data <= 7'h00; 
        10'b0100010000: data <= 7'h00; 
        10'b0100010001: data <= 7'h00; 
        10'b0100010010: data <= 7'h7f; 
        10'b0100010011: data <= 7'h00; 
        10'b0100010100: data <= 7'h00; 
        10'b0100010101: data <= 7'h00; 
        10'b0100010110: data <= 7'h00; 
        10'b0100010111: data <= 7'h00; 
        10'b0100011000: data <= 7'h00; 
        10'b0100011001: data <= 7'h00; 
        10'b0100011010: data <= 7'h00; 
        10'b0100011011: data <= 7'h00; 
        10'b0100011100: data <= 7'h00; 
        10'b0100011101: data <= 7'h00; 
        10'b0100011110: data <= 7'h00; 
        10'b0100011111: data <= 7'h00; 
        10'b0100100000: data <= 7'h00; 
        10'b0100100001: data <= 7'h00; 
        10'b0100100010: data <= 7'h00; 
        10'b0100100011: data <= 7'h00; 
        10'b0100100100: data <= 7'h00; 
        10'b0100100101: data <= 7'h00; 
        10'b0100100110: data <= 7'h01; 
        10'b0100100111: data <= 7'h01; 
        10'b0100101000: data <= 7'h00; 
        10'b0100101001: data <= 7'h00; 
        10'b0100101010: data <= 7'h00; 
        10'b0100101011: data <= 7'h00; 
        10'b0100101100: data <= 7'h00; 
        10'b0100101101: data <= 7'h00; 
        10'b0100101110: data <= 7'h00; 
        10'b0100101111: data <= 7'h00; 
        10'b0100110000: data <= 7'h00; 
        10'b0100110001: data <= 7'h00; 
        10'b0100110010: data <= 7'h00; 
        10'b0100110011: data <= 7'h00; 
        10'b0100110100: data <= 7'h00; 
        10'b0100110101: data <= 7'h00; 
        10'b0100110110: data <= 7'h00; 
        10'b0100110111: data <= 7'h00; 
        10'b0100111000: data <= 7'h00; 
        10'b0100111001: data <= 7'h00; 
        10'b0100111010: data <= 7'h00; 
        10'b0100111011: data <= 7'h00; 
        10'b0100111100: data <= 7'h00; 
        10'b0100111101: data <= 7'h00; 
        10'b0100111110: data <= 7'h00; 
        10'b0100111111: data <= 7'h00; 
        10'b0101000000: data <= 7'h00; 
        10'b0101000001: data <= 7'h01; 
        10'b0101000010: data <= 7'h01; 
        10'b0101000011: data <= 7'h01; 
        10'b0101000100: data <= 7'h00; 
        10'b0101000101: data <= 7'h00; 
        10'b0101000110: data <= 7'h00; 
        10'b0101000111: data <= 7'h00; 
        10'b0101001000: data <= 7'h00; 
        10'b0101001001: data <= 7'h00; 
        10'b0101001010: data <= 7'h00; 
        10'b0101001011: data <= 7'h00; 
        10'b0101001100: data <= 7'h00; 
        10'b0101001101: data <= 7'h00; 
        10'b0101001110: data <= 7'h00; 
        10'b0101001111: data <= 7'h00; 
        10'b0101010000: data <= 7'h00; 
        10'b0101010001: data <= 7'h00; 
        10'b0101010010: data <= 7'h00; 
        10'b0101010011: data <= 7'h00; 
        10'b0101010100: data <= 7'h00; 
        10'b0101010101: data <= 7'h00; 
        10'b0101010110: data <= 7'h00; 
        10'b0101010111: data <= 7'h00; 
        10'b0101011000: data <= 7'h00; 
        10'b0101011001: data <= 7'h00; 
        10'b0101011010: data <= 7'h00; 
        10'b0101011011: data <= 7'h7f; 
        10'b0101011100: data <= 7'h00; 
        10'b0101011101: data <= 7'h01; 
        10'b0101011110: data <= 7'h01; 
        10'b0101011111: data <= 7'h01; 
        10'b0101100000: data <= 7'h00; 
        10'b0101100001: data <= 7'h00; 
        10'b0101100010: data <= 7'h00; 
        10'b0101100011: data <= 7'h00; 
        10'b0101100100: data <= 7'h00; 
        10'b0101100101: data <= 7'h00; 
        10'b0101100110: data <= 7'h00; 
        10'b0101100111: data <= 7'h00; 
        10'b0101101000: data <= 7'h00; 
        10'b0101101001: data <= 7'h00; 
        10'b0101101010: data <= 7'h00; 
        10'b0101101011: data <= 7'h00; 
        10'b0101101100: data <= 7'h00; 
        10'b0101101101: data <= 7'h00; 
        10'b0101101110: data <= 7'h00; 
        10'b0101101111: data <= 7'h00; 
        10'b0101110000: data <= 7'h00; 
        10'b0101110001: data <= 7'h00; 
        10'b0101110010: data <= 7'h00; 
        10'b0101110011: data <= 7'h00; 
        10'b0101110100: data <= 7'h00; 
        10'b0101110101: data <= 7'h00; 
        10'b0101110110: data <= 7'h7f; 
        10'b0101110111: data <= 7'h7f; 
        10'b0101111000: data <= 7'h00; 
        10'b0101111001: data <= 7'h00; 
        10'b0101111010: data <= 7'h01; 
        10'b0101111011: data <= 7'h01; 
        10'b0101111100: data <= 7'h00; 
        10'b0101111101: data <= 7'h00; 
        10'b0101111110: data <= 7'h00; 
        10'b0101111111: data <= 7'h00; 
        10'b0110000000: data <= 7'h00; 
        10'b0110000001: data <= 7'h00; 
        10'b0110000010: data <= 7'h00; 
        10'b0110000011: data <= 7'h00; 
        10'b0110000100: data <= 7'h00; 
        10'b0110000101: data <= 7'h00; 
        10'b0110000110: data <= 7'h00; 
        10'b0110000111: data <= 7'h00; 
        10'b0110001000: data <= 7'h00; 
        10'b0110001001: data <= 7'h00; 
        10'b0110001010: data <= 7'h00; 
        10'b0110001011: data <= 7'h00; 
        10'b0110001100: data <= 7'h00; 
        10'b0110001101: data <= 7'h00; 
        10'b0110001110: data <= 7'h00; 
        10'b0110001111: data <= 7'h00; 
        10'b0110010000: data <= 7'h00; 
        10'b0110010001: data <= 7'h00; 
        10'b0110010010: data <= 7'h7f; 
        10'b0110010011: data <= 7'h7f; 
        10'b0110010100: data <= 7'h00; 
        10'b0110010101: data <= 7'h00; 
        10'b0110010110: data <= 7'h01; 
        10'b0110010111: data <= 7'h01; 
        10'b0110011000: data <= 7'h00; 
        10'b0110011001: data <= 7'h00; 
        10'b0110011010: data <= 7'h00; 
        10'b0110011011: data <= 7'h00; 
        10'b0110011100: data <= 7'h00; 
        10'b0110011101: data <= 7'h00; 
        10'b0110011110: data <= 7'h00; 
        10'b0110011111: data <= 7'h00; 
        10'b0110100000: data <= 7'h00; 
        10'b0110100001: data <= 7'h00; 
        10'b0110100010: data <= 7'h00; 
        10'b0110100011: data <= 7'h00; 
        10'b0110100100: data <= 7'h00; 
        10'b0110100101: data <= 7'h00; 
        10'b0110100110: data <= 7'h00; 
        10'b0110100111: data <= 7'h00; 
        10'b0110101000: data <= 7'h00; 
        10'b0110101001: data <= 7'h00; 
        10'b0110101010: data <= 7'h00; 
        10'b0110101011: data <= 7'h00; 
        10'b0110101100: data <= 7'h00; 
        10'b0110101101: data <= 7'h00; 
        10'b0110101110: data <= 7'h7f; 
        10'b0110101111: data <= 7'h00; 
        10'b0110110000: data <= 7'h00; 
        10'b0110110001: data <= 7'h01; 
        10'b0110110010: data <= 7'h01; 
        10'b0110110011: data <= 7'h00; 
        10'b0110110100: data <= 7'h00; 
        10'b0110110101: data <= 7'h7f; 
        10'b0110110110: data <= 7'h7f; 
        10'b0110110111: data <= 7'h00; 
        10'b0110111000: data <= 7'h00; 
        10'b0110111001: data <= 7'h00; 
        10'b0110111010: data <= 7'h00; 
        10'b0110111011: data <= 7'h00; 
        10'b0110111100: data <= 7'h00; 
        10'b0110111101: data <= 7'h00; 
        10'b0110111110: data <= 7'h00; 
        10'b0110111111: data <= 7'h00; 
        10'b0111000000: data <= 7'h00; 
        10'b0111000001: data <= 7'h00; 
        10'b0111000010: data <= 7'h00; 
        10'b0111000011: data <= 7'h00; 
        10'b0111000100: data <= 7'h00; 
        10'b0111000101: data <= 7'h00; 
        10'b0111000110: data <= 7'h00; 
        10'b0111000111: data <= 7'h00; 
        10'b0111001000: data <= 7'h00; 
        10'b0111001001: data <= 7'h00; 
        10'b0111001010: data <= 7'h00; 
        10'b0111001011: data <= 7'h00; 
        10'b0111001100: data <= 7'h00; 
        10'b0111001101: data <= 7'h01; 
        10'b0111001110: data <= 7'h01; 
        10'b0111001111: data <= 7'h00; 
        10'b0111010000: data <= 7'h00; 
        10'b0111010001: data <= 7'h7f; 
        10'b0111010010: data <= 7'h7f; 
        10'b0111010011: data <= 7'h00; 
        10'b0111010100: data <= 7'h00; 
        10'b0111010101: data <= 7'h00; 
        10'b0111010110: data <= 7'h00; 
        10'b0111010111: data <= 7'h00; 
        10'b0111011000: data <= 7'h00; 
        10'b0111011001: data <= 7'h00; 
        10'b0111011010: data <= 7'h00; 
        10'b0111011011: data <= 7'h00; 
        10'b0111011100: data <= 7'h00; 
        10'b0111011101: data <= 7'h00; 
        10'b0111011110: data <= 7'h00; 
        10'b0111011111: data <= 7'h00; 
        10'b0111100000: data <= 7'h00; 
        10'b0111100001: data <= 7'h00; 
        10'b0111100010: data <= 7'h00; 
        10'b0111100011: data <= 7'h00; 
        10'b0111100100: data <= 7'h00; 
        10'b0111100101: data <= 7'h00; 
        10'b0111100110: data <= 7'h00; 
        10'b0111100111: data <= 7'h00; 
        10'b0111101000: data <= 7'h00; 
        10'b0111101001: data <= 7'h01; 
        10'b0111101010: data <= 7'h01; 
        10'b0111101011: data <= 7'h00; 
        10'b0111101100: data <= 7'h7f; 
        10'b0111101101: data <= 7'h7f; 
        10'b0111101110: data <= 7'h7f; 
        10'b0111101111: data <= 7'h00; 
        10'b0111110000: data <= 7'h00; 
        10'b0111110001: data <= 7'h00; 
        10'b0111110010: data <= 7'h00; 
        10'b0111110011: data <= 7'h00; 
        10'b0111110100: data <= 7'h00; 
        10'b0111110101: data <= 7'h00; 
        10'b0111110110: data <= 7'h00; 
        10'b0111110111: data <= 7'h00; 
        10'b0111111000: data <= 7'h00; 
        10'b0111111001: data <= 7'h00; 
        10'b0111111010: data <= 7'h00; 
        10'b0111111011: data <= 7'h00; 
        10'b0111111100: data <= 7'h00; 
        10'b0111111101: data <= 7'h00; 
        10'b0111111110: data <= 7'h00; 
        10'b0111111111: data <= 7'h00; 
        10'b1000000000: data <= 7'h00; 
        10'b1000000001: data <= 7'h00; 
        10'b1000000010: data <= 7'h00; 
        10'b1000000011: data <= 7'h00; 
        10'b1000000100: data <= 7'h00; 
        10'b1000000101: data <= 7'h01; 
        10'b1000000110: data <= 7'h00; 
        10'b1000000111: data <= 7'h00; 
        10'b1000001000: data <= 7'h7f; 
        10'b1000001001: data <= 7'h00; 
        10'b1000001010: data <= 7'h00; 
        10'b1000001011: data <= 7'h00; 
        10'b1000001100: data <= 7'h00; 
        10'b1000001101: data <= 7'h00; 
        10'b1000001110: data <= 7'h00; 
        10'b1000001111: data <= 7'h00; 
        10'b1000010000: data <= 7'h00; 
        10'b1000010001: data <= 7'h00; 
        10'b1000010010: data <= 7'h00; 
        10'b1000010011: data <= 7'h00; 
        10'b1000010100: data <= 7'h00; 
        10'b1000010101: data <= 7'h00; 
        10'b1000010110: data <= 7'h00; 
        10'b1000010111: data <= 7'h00; 
        10'b1000011000: data <= 7'h00; 
        10'b1000011001: data <= 7'h00; 
        10'b1000011010: data <= 7'h00; 
        10'b1000011011: data <= 7'h00; 
        10'b1000011100: data <= 7'h00; 
        10'b1000011101: data <= 7'h00; 
        10'b1000011110: data <= 7'h00; 
        10'b1000011111: data <= 7'h00; 
        10'b1000100000: data <= 7'h00; 
        10'b1000100001: data <= 7'h00; 
        10'b1000100010: data <= 7'h00; 
        10'b1000100011: data <= 7'h00; 
        10'b1000100100: data <= 7'h00; 
        10'b1000100101: data <= 7'h00; 
        10'b1000100110: data <= 7'h00; 
        10'b1000100111: data <= 7'h00; 
        10'b1000101000: data <= 7'h00; 
        10'b1000101001: data <= 7'h00; 
        10'b1000101010: data <= 7'h00; 
        10'b1000101011: data <= 7'h00; 
        10'b1000101100: data <= 7'h00; 
        10'b1000101101: data <= 7'h00; 
        10'b1000101110: data <= 7'h00; 
        10'b1000101111: data <= 7'h00; 
        10'b1000110000: data <= 7'h00; 
        10'b1000110001: data <= 7'h00; 
        10'b1000110010: data <= 7'h00; 
        10'b1000110011: data <= 7'h00; 
        10'b1000110100: data <= 7'h00; 
        10'b1000110101: data <= 7'h00; 
        10'b1000110110: data <= 7'h00; 
        10'b1000110111: data <= 7'h00; 
        10'b1000111000: data <= 7'h00; 
        10'b1000111001: data <= 7'h00; 
        10'b1000111010: data <= 7'h00; 
        10'b1000111011: data <= 7'h00; 
        10'b1000111100: data <= 7'h00; 
        10'b1000111101: data <= 7'h00; 
        10'b1000111110: data <= 7'h00; 
        10'b1000111111: data <= 7'h00; 
        10'b1001000000: data <= 7'h00; 
        10'b1001000001: data <= 7'h00; 
        10'b1001000010: data <= 7'h00; 
        10'b1001000011: data <= 7'h00; 
        10'b1001000100: data <= 7'h00; 
        10'b1001000101: data <= 7'h00; 
        10'b1001000110: data <= 7'h00; 
        10'b1001000111: data <= 7'h00; 
        10'b1001001000: data <= 7'h00; 
        10'b1001001001: data <= 7'h00; 
        10'b1001001010: data <= 7'h00; 
        10'b1001001011: data <= 7'h00; 
        10'b1001001100: data <= 7'h00; 
        10'b1001001101: data <= 7'h00; 
        10'b1001001110: data <= 7'h00; 
        10'b1001001111: data <= 7'h00; 
        10'b1001010000: data <= 7'h00; 
        10'b1001010001: data <= 7'h00; 
        10'b1001010010: data <= 7'h00; 
        10'b1001010011: data <= 7'h00; 
        10'b1001010100: data <= 7'h00; 
        10'b1001010101: data <= 7'h00; 
        10'b1001010110: data <= 7'h00; 
        10'b1001010111: data <= 7'h00; 
        10'b1001011000: data <= 7'h00; 
        10'b1001011001: data <= 7'h00; 
        10'b1001011010: data <= 7'h00; 
        10'b1001011011: data <= 7'h00; 
        10'b1001011100: data <= 7'h00; 
        10'b1001011101: data <= 7'h00; 
        10'b1001011110: data <= 7'h00; 
        10'b1001011111: data <= 7'h00; 
        10'b1001100000: data <= 7'h00; 
        10'b1001100001: data <= 7'h00; 
        10'b1001100010: data <= 7'h00; 
        10'b1001100011: data <= 7'h00; 
        10'b1001100100: data <= 7'h00; 
        10'b1001100101: data <= 7'h00; 
        10'b1001100110: data <= 7'h00; 
        10'b1001100111: data <= 7'h00; 
        10'b1001101000: data <= 7'h00; 
        10'b1001101001: data <= 7'h00; 
        10'b1001101010: data <= 7'h00; 
        10'b1001101011: data <= 7'h00; 
        10'b1001101100: data <= 7'h00; 
        10'b1001101101: data <= 7'h00; 
        10'b1001101110: data <= 7'h00; 
        10'b1001101111: data <= 7'h00; 
        10'b1001110000: data <= 7'h00; 
        10'b1001110001: data <= 7'h00; 
        10'b1001110010: data <= 7'h00; 
        10'b1001110011: data <= 7'h00; 
        10'b1001110100: data <= 7'h7f; 
        10'b1001110101: data <= 7'h7f; 
        10'b1001110110: data <= 7'h00; 
        10'b1001110111: data <= 7'h00; 
        10'b1001111000: data <= 7'h00; 
        10'b1001111001: data <= 7'h01; 
        10'b1001111010: data <= 7'h00; 
        10'b1001111011: data <= 7'h00; 
        10'b1001111100: data <= 7'h00; 
        10'b1001111101: data <= 7'h00; 
        10'b1001111110: data <= 7'h00; 
        10'b1001111111: data <= 7'h00; 
        10'b1010000000: data <= 7'h00; 
        10'b1010000001: data <= 7'h00; 
        10'b1010000010: data <= 7'h00; 
        10'b1010000011: data <= 7'h00; 
        10'b1010000100: data <= 7'h00; 
        10'b1010000101: data <= 7'h00; 
        10'b1010000110: data <= 7'h00; 
        10'b1010000111: data <= 7'h00; 
        10'b1010001000: data <= 7'h00; 
        10'b1010001001: data <= 7'h00; 
        10'b1010001010: data <= 7'h00; 
        10'b1010001011: data <= 7'h00; 
        10'b1010001100: data <= 7'h00; 
        10'b1010001101: data <= 7'h00; 
        10'b1010001110: data <= 7'h00; 
        10'b1010001111: data <= 7'h00; 
        10'b1010010000: data <= 7'h00; 
        10'b1010010001: data <= 7'h00; 
        10'b1010010010: data <= 7'h00; 
        10'b1010010011: data <= 7'h00; 
        10'b1010010100: data <= 7'h00; 
        10'b1010010101: data <= 7'h01; 
        10'b1010010110: data <= 7'h00; 
        10'b1010010111: data <= 7'h00; 
        10'b1010011000: data <= 7'h00; 
        10'b1010011001: data <= 7'h00; 
        10'b1010011010: data <= 7'h00; 
        10'b1010011011: data <= 7'h00; 
        10'b1010011100: data <= 7'h00; 
        10'b1010011101: data <= 7'h00; 
        10'b1010011110: data <= 7'h00; 
        10'b1010011111: data <= 7'h00; 
        10'b1010100000: data <= 7'h00; 
        10'b1010100001: data <= 7'h00; 
        10'b1010100010: data <= 7'h00; 
        10'b1010100011: data <= 7'h00; 
        10'b1010100100: data <= 7'h00; 
        10'b1010100101: data <= 7'h00; 
        10'b1010100110: data <= 7'h00; 
        10'b1010100111: data <= 7'h00; 
        10'b1010101000: data <= 7'h00; 
        10'b1010101001: data <= 7'h00; 
        10'b1010101010: data <= 7'h00; 
        10'b1010101011: data <= 7'h00; 
        10'b1010101100: data <= 7'h00; 
        10'b1010101101: data <= 7'h00; 
        10'b1010101110: data <= 7'h00; 
        10'b1010101111: data <= 7'h00; 
        10'b1010110000: data <= 7'h00; 
        10'b1010110001: data <= 7'h00; 
        10'b1010110010: data <= 7'h00; 
        10'b1010110011: data <= 7'h00; 
        10'b1010110100: data <= 7'h00; 
        10'b1010110101: data <= 7'h00; 
        10'b1010110110: data <= 7'h00; 
        10'b1010110111: data <= 7'h00; 
        10'b1010111000: data <= 7'h00; 
        10'b1010111001: data <= 7'h00; 
        10'b1010111010: data <= 7'h00; 
        10'b1010111011: data <= 7'h00; 
        10'b1010111100: data <= 7'h00; 
        10'b1010111101: data <= 7'h00; 
        10'b1010111110: data <= 7'h00; 
        10'b1010111111: data <= 7'h00; 
        10'b1011000000: data <= 7'h00; 
        10'b1011000001: data <= 7'h00; 
        10'b1011000010: data <= 7'h00; 
        10'b1011000011: data <= 7'h00; 
        10'b1011000100: data <= 7'h00; 
        10'b1011000101: data <= 7'h00; 
        10'b1011000110: data <= 7'h00; 
        10'b1011000111: data <= 7'h00; 
        10'b1011001000: data <= 7'h00; 
        10'b1011001001: data <= 7'h00; 
        10'b1011001010: data <= 7'h00; 
        10'b1011001011: data <= 7'h00; 
        10'b1011001100: data <= 7'h00; 
        10'b1011001101: data <= 7'h00; 
        10'b1011001110: data <= 7'h00; 
        10'b1011001111: data <= 7'h00; 
        10'b1011010000: data <= 7'h00; 
        10'b1011010001: data <= 7'h00; 
        10'b1011010010: data <= 7'h00; 
        10'b1011010011: data <= 7'h00; 
        10'b1011010100: data <= 7'h00; 
        10'b1011010101: data <= 7'h00; 
        10'b1011010110: data <= 7'h00; 
        10'b1011010111: data <= 7'h00; 
        10'b1011011000: data <= 7'h00; 
        10'b1011011001: data <= 7'h00; 
        10'b1011011010: data <= 7'h00; 
        10'b1011011011: data <= 7'h00; 
        10'b1011011100: data <= 7'h00; 
        10'b1011011101: data <= 7'h00; 
        10'b1011011110: data <= 7'h00; 
        10'b1011011111: data <= 7'h00; 
        10'b1011100000: data <= 7'h00; 
        10'b1011100001: data <= 7'h00; 
        10'b1011100010: data <= 7'h00; 
        10'b1011100011: data <= 7'h00; 
        10'b1011100100: data <= 7'h00; 
        10'b1011100101: data <= 7'h00; 
        10'b1011100110: data <= 7'h00; 
        10'b1011100111: data <= 7'h00; 
        10'b1011101000: data <= 7'h00; 
        10'b1011101001: data <= 7'h00; 
        10'b1011101010: data <= 7'h00; 
        10'b1011101011: data <= 7'h00; 
        10'b1011101100: data <= 7'h00; 
        10'b1011101101: data <= 7'h00; 
        10'b1011101110: data <= 7'h00; 
        10'b1011101111: data <= 7'h00; 
        10'b1011110000: data <= 7'h00; 
        10'b1011110001: data <= 7'h00; 
        10'b1011110010: data <= 7'h00; 
        10'b1011110011: data <= 7'h00; 
        10'b1011110100: data <= 7'h00; 
        10'b1011110101: data <= 7'h00; 
        10'b1011110110: data <= 7'h00; 
        10'b1011110111: data <= 7'h00; 
        10'b1011111000: data <= 7'h00; 
        10'b1011111001: data <= 7'h00; 
        10'b1011111010: data <= 7'h00; 
        10'b1011111011: data <= 7'h00; 
        10'b1011111100: data <= 7'h00; 
        10'b1011111101: data <= 7'h00; 
        10'b1011111110: data <= 7'h00; 
        10'b1011111111: data <= 7'h00; 
        10'b1100000000: data <= 7'h00; 
        10'b1100000001: data <= 7'h00; 
        10'b1100000010: data <= 7'h00; 
        10'b1100000011: data <= 7'h00; 
        10'b1100000100: data <= 7'h00; 
        10'b1100000101: data <= 7'h00; 
        10'b1100000110: data <= 7'h00; 
        10'b1100000111: data <= 7'h00; 
        10'b1100001000: data <= 7'h00; 
        10'b1100001001: data <= 7'h00; 
        10'b1100001010: data <= 7'h00; 
        10'b1100001011: data <= 7'h00; 
        10'b1100001100: data <= 7'h00; 
        10'b1100001101: data <= 7'h00; 
        10'b1100001110: data <= 7'h00; 
        10'b1100001111: data <= 7'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 2) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 8'h00; 
        10'b0000000001: data <= 8'h00; 
        10'b0000000010: data <= 8'h00; 
        10'b0000000011: data <= 8'h00; 
        10'b0000000100: data <= 8'h00; 
        10'b0000000101: data <= 8'h00; 
        10'b0000000110: data <= 8'h00; 
        10'b0000000111: data <= 8'h00; 
        10'b0000001000: data <= 8'h00; 
        10'b0000001001: data <= 8'h00; 
        10'b0000001010: data <= 8'h00; 
        10'b0000001011: data <= 8'h00; 
        10'b0000001100: data <= 8'h00; 
        10'b0000001101: data <= 8'h00; 
        10'b0000001110: data <= 8'h00; 
        10'b0000001111: data <= 8'h00; 
        10'b0000010000: data <= 8'h00; 
        10'b0000010001: data <= 8'h00; 
        10'b0000010010: data <= 8'h00; 
        10'b0000010011: data <= 8'h00; 
        10'b0000010100: data <= 8'h00; 
        10'b0000010101: data <= 8'h00; 
        10'b0000010110: data <= 8'h00; 
        10'b0000010111: data <= 8'h00; 
        10'b0000011000: data <= 8'h00; 
        10'b0000011001: data <= 8'h00; 
        10'b0000011010: data <= 8'h00; 
        10'b0000011011: data <= 8'h00; 
        10'b0000011100: data <= 8'h00; 
        10'b0000011101: data <= 8'h00; 
        10'b0000011110: data <= 8'h00; 
        10'b0000011111: data <= 8'h00; 
        10'b0000100000: data <= 8'h00; 
        10'b0000100001: data <= 8'h00; 
        10'b0000100010: data <= 8'h00; 
        10'b0000100011: data <= 8'h00; 
        10'b0000100100: data <= 8'h00; 
        10'b0000100101: data <= 8'h00; 
        10'b0000100110: data <= 8'h00; 
        10'b0000100111: data <= 8'h00; 
        10'b0000101000: data <= 8'h00; 
        10'b0000101001: data <= 8'h00; 
        10'b0000101010: data <= 8'h00; 
        10'b0000101011: data <= 8'h00; 
        10'b0000101100: data <= 8'h00; 
        10'b0000101101: data <= 8'h00; 
        10'b0000101110: data <= 8'h00; 
        10'b0000101111: data <= 8'h00; 
        10'b0000110000: data <= 8'h00; 
        10'b0000110001: data <= 8'h00; 
        10'b0000110010: data <= 8'h00; 
        10'b0000110011: data <= 8'h00; 
        10'b0000110100: data <= 8'h00; 
        10'b0000110101: data <= 8'h00; 
        10'b0000110110: data <= 8'h00; 
        10'b0000110111: data <= 8'h00; 
        10'b0000111000: data <= 8'h00; 
        10'b0000111001: data <= 8'h00; 
        10'b0000111010: data <= 8'h00; 
        10'b0000111011: data <= 8'h00; 
        10'b0000111100: data <= 8'h00; 
        10'b0000111101: data <= 8'h00; 
        10'b0000111110: data <= 8'h00; 
        10'b0000111111: data <= 8'h00; 
        10'b0001000000: data <= 8'h00; 
        10'b0001000001: data <= 8'h00; 
        10'b0001000010: data <= 8'h00; 
        10'b0001000011: data <= 8'h00; 
        10'b0001000100: data <= 8'h00; 
        10'b0001000101: data <= 8'h00; 
        10'b0001000110: data <= 8'h00; 
        10'b0001000111: data <= 8'h00; 
        10'b0001001000: data <= 8'h00; 
        10'b0001001001: data <= 8'h00; 
        10'b0001001010: data <= 8'h00; 
        10'b0001001011: data <= 8'h00; 
        10'b0001001100: data <= 8'h00; 
        10'b0001001101: data <= 8'h00; 
        10'b0001001110: data <= 8'h00; 
        10'b0001001111: data <= 8'h00; 
        10'b0001010000: data <= 8'h00; 
        10'b0001010001: data <= 8'h00; 
        10'b0001010010: data <= 8'h00; 
        10'b0001010011: data <= 8'h00; 
        10'b0001010100: data <= 8'h00; 
        10'b0001010101: data <= 8'h00; 
        10'b0001010110: data <= 8'h00; 
        10'b0001010111: data <= 8'h00; 
        10'b0001011000: data <= 8'h00; 
        10'b0001011001: data <= 8'h00; 
        10'b0001011010: data <= 8'h00; 
        10'b0001011011: data <= 8'h00; 
        10'b0001011100: data <= 8'h00; 
        10'b0001011101: data <= 8'h00; 
        10'b0001011110: data <= 8'h00; 
        10'b0001011111: data <= 8'h00; 
        10'b0001100000: data <= 8'h00; 
        10'b0001100001: data <= 8'h00; 
        10'b0001100010: data <= 8'h00; 
        10'b0001100011: data <= 8'h00; 
        10'b0001100100: data <= 8'h00; 
        10'b0001100101: data <= 8'h00; 
        10'b0001100110: data <= 8'h00; 
        10'b0001100111: data <= 8'h00; 
        10'b0001101000: data <= 8'h00; 
        10'b0001101001: data <= 8'h00; 
        10'b0001101010: data <= 8'h00; 
        10'b0001101011: data <= 8'h00; 
        10'b0001101100: data <= 8'h00; 
        10'b0001101101: data <= 8'h00; 
        10'b0001101110: data <= 8'h00; 
        10'b0001101111: data <= 8'h00; 
        10'b0001110000: data <= 8'h00; 
        10'b0001110001: data <= 8'h00; 
        10'b0001110010: data <= 8'h00; 
        10'b0001110011: data <= 8'h00; 
        10'b0001110100: data <= 8'h00; 
        10'b0001110101: data <= 8'h00; 
        10'b0001110110: data <= 8'h00; 
        10'b0001110111: data <= 8'h00; 
        10'b0001111000: data <= 8'h00; 
        10'b0001111001: data <= 8'h00; 
        10'b0001111010: data <= 8'h00; 
        10'b0001111011: data <= 8'h00; 
        10'b0001111100: data <= 8'h00; 
        10'b0001111101: data <= 8'h00; 
        10'b0001111110: data <= 8'h00; 
        10'b0001111111: data <= 8'h01; 
        10'b0010000000: data <= 8'h00; 
        10'b0010000001: data <= 8'h00; 
        10'b0010000010: data <= 8'h00; 
        10'b0010000011: data <= 8'h00; 
        10'b0010000100: data <= 8'h00; 
        10'b0010000101: data <= 8'h00; 
        10'b0010000110: data <= 8'h00; 
        10'b0010000111: data <= 8'h00; 
        10'b0010001000: data <= 8'h00; 
        10'b0010001001: data <= 8'h00; 
        10'b0010001010: data <= 8'h00; 
        10'b0010001011: data <= 8'h00; 
        10'b0010001100: data <= 8'h00; 
        10'b0010001101: data <= 8'h00; 
        10'b0010001110: data <= 8'h00; 
        10'b0010001111: data <= 8'h00; 
        10'b0010010000: data <= 8'h00; 
        10'b0010010001: data <= 8'h00; 
        10'b0010010010: data <= 8'h00; 
        10'b0010010011: data <= 8'h00; 
        10'b0010010100: data <= 8'hff; 
        10'b0010010101: data <= 8'hff; 
        10'b0010010110: data <= 8'h00; 
        10'b0010010111: data <= 8'h00; 
        10'b0010011000: data <= 8'h00; 
        10'b0010011001: data <= 8'h00; 
        10'b0010011010: data <= 8'h00; 
        10'b0010011011: data <= 8'h00; 
        10'b0010011100: data <= 8'h00; 
        10'b0010011101: data <= 8'h00; 
        10'b0010011110: data <= 8'h00; 
        10'b0010011111: data <= 8'h00; 
        10'b0010100000: data <= 8'h00; 
        10'b0010100001: data <= 8'h00; 
        10'b0010100010: data <= 8'h01; 
        10'b0010100011: data <= 8'h01; 
        10'b0010100100: data <= 8'h00; 
        10'b0010100101: data <= 8'h00; 
        10'b0010100110: data <= 8'h00; 
        10'b0010100111: data <= 8'h00; 
        10'b0010101000: data <= 8'h00; 
        10'b0010101001: data <= 8'h00; 
        10'b0010101010: data <= 8'h00; 
        10'b0010101011: data <= 8'h00; 
        10'b0010101100: data <= 8'h00; 
        10'b0010101101: data <= 8'h00; 
        10'b0010101110: data <= 8'h00; 
        10'b0010101111: data <= 8'h00; 
        10'b0010110000: data <= 8'hff; 
        10'b0010110001: data <= 8'hff; 
        10'b0010110010: data <= 8'hff; 
        10'b0010110011: data <= 8'h00; 
        10'b0010110100: data <= 8'h00; 
        10'b0010110101: data <= 8'h00; 
        10'b0010110110: data <= 8'h00; 
        10'b0010110111: data <= 8'hff; 
        10'b0010111000: data <= 8'hff; 
        10'b0010111001: data <= 8'hff; 
        10'b0010111010: data <= 8'h00; 
        10'b0010111011: data <= 8'h00; 
        10'b0010111100: data <= 8'h00; 
        10'b0010111101: data <= 8'h01; 
        10'b0010111110: data <= 8'h00; 
        10'b0010111111: data <= 8'h00; 
        10'b0011000000: data <= 8'h00; 
        10'b0011000001: data <= 8'h00; 
        10'b0011000010: data <= 8'h00; 
        10'b0011000011: data <= 8'h00; 
        10'b0011000100: data <= 8'h00; 
        10'b0011000101: data <= 8'h00; 
        10'b0011000110: data <= 8'h00; 
        10'b0011000111: data <= 8'h00; 
        10'b0011001000: data <= 8'h00; 
        10'b0011001001: data <= 8'h00; 
        10'b0011001010: data <= 8'h00; 
        10'b0011001011: data <= 8'hff; 
        10'b0011001100: data <= 8'hff; 
        10'b0011001101: data <= 8'hff; 
        10'b0011001110: data <= 8'hff; 
        10'b0011001111: data <= 8'h00; 
        10'b0011010000: data <= 8'h00; 
        10'b0011010001: data <= 8'h00; 
        10'b0011010010: data <= 8'hff; 
        10'b0011010011: data <= 8'hff; 
        10'b0011010100: data <= 8'hff; 
        10'b0011010101: data <= 8'hff; 
        10'b0011010110: data <= 8'hff; 
        10'b0011010111: data <= 8'h00; 
        10'b0011011000: data <= 8'h00; 
        10'b0011011001: data <= 8'h00; 
        10'b0011011010: data <= 8'h00; 
        10'b0011011011: data <= 8'h00; 
        10'b0011011100: data <= 8'h00; 
        10'b0011011101: data <= 8'h00; 
        10'b0011011110: data <= 8'h00; 
        10'b0011011111: data <= 8'h00; 
        10'b0011100000: data <= 8'h00; 
        10'b0011100001: data <= 8'h00; 
        10'b0011100010: data <= 8'h00; 
        10'b0011100011: data <= 8'h00; 
        10'b0011100100: data <= 8'h00; 
        10'b0011100101: data <= 8'h00; 
        10'b0011100110: data <= 8'h00; 
        10'b0011100111: data <= 8'hff; 
        10'b0011101000: data <= 8'hff; 
        10'b0011101001: data <= 8'hff; 
        10'b0011101010: data <= 8'hff; 
        10'b0011101011: data <= 8'hff; 
        10'b0011101100: data <= 8'h00; 
        10'b0011101101: data <= 8'h00; 
        10'b0011101110: data <= 8'h00; 
        10'b0011101111: data <= 8'h00; 
        10'b0011110000: data <= 8'h00; 
        10'b0011110001: data <= 8'h00; 
        10'b0011110010: data <= 8'h00; 
        10'b0011110011: data <= 8'h00; 
        10'b0011110100: data <= 8'h00; 
        10'b0011110101: data <= 8'h00; 
        10'b0011110110: data <= 8'hff; 
        10'b0011110111: data <= 8'hff; 
        10'b0011111000: data <= 8'hff; 
        10'b0011111001: data <= 8'h00; 
        10'b0011111010: data <= 8'h00; 
        10'b0011111011: data <= 8'h00; 
        10'b0011111100: data <= 8'h00; 
        10'b0011111101: data <= 8'h00; 
        10'b0011111110: data <= 8'h00; 
        10'b0011111111: data <= 8'h00; 
        10'b0100000000: data <= 8'h00; 
        10'b0100000001: data <= 8'h00; 
        10'b0100000010: data <= 8'h00; 
        10'b0100000011: data <= 8'h00; 
        10'b0100000100: data <= 8'hff; 
        10'b0100000101: data <= 8'hff; 
        10'b0100000110: data <= 8'hff; 
        10'b0100000111: data <= 8'h00; 
        10'b0100001000: data <= 8'h00; 
        10'b0100001001: data <= 8'h00; 
        10'b0100001010: data <= 8'h01; 
        10'b0100001011: data <= 8'h01; 
        10'b0100001100: data <= 8'h00; 
        10'b0100001101: data <= 8'h00; 
        10'b0100001110: data <= 8'h00; 
        10'b0100001111: data <= 8'hff; 
        10'b0100010000: data <= 8'hff; 
        10'b0100010001: data <= 8'hff; 
        10'b0100010010: data <= 8'hff; 
        10'b0100010011: data <= 8'hff; 
        10'b0100010100: data <= 8'hff; 
        10'b0100010101: data <= 8'h00; 
        10'b0100010110: data <= 8'h00; 
        10'b0100010111: data <= 8'h00; 
        10'b0100011000: data <= 8'h00; 
        10'b0100011001: data <= 8'h00; 
        10'b0100011010: data <= 8'h00; 
        10'b0100011011: data <= 8'h00; 
        10'b0100011100: data <= 8'h00; 
        10'b0100011101: data <= 8'h00; 
        10'b0100011110: data <= 8'h00; 
        10'b0100011111: data <= 8'h00; 
        10'b0100100000: data <= 8'hff; 
        10'b0100100001: data <= 8'hff; 
        10'b0100100010: data <= 8'h00; 
        10'b0100100011: data <= 8'h00; 
        10'b0100100100: data <= 8'h00; 
        10'b0100100101: data <= 8'h01; 
        10'b0100100110: data <= 8'h02; 
        10'b0100100111: data <= 8'h02; 
        10'b0100101000: data <= 8'h01; 
        10'b0100101001: data <= 8'h00; 
        10'b0100101010: data <= 8'hff; 
        10'b0100101011: data <= 8'hff; 
        10'b0100101100: data <= 8'hff; 
        10'b0100101101: data <= 8'hff; 
        10'b0100101110: data <= 8'hff; 
        10'b0100101111: data <= 8'h00; 
        10'b0100110000: data <= 8'h00; 
        10'b0100110001: data <= 8'h00; 
        10'b0100110010: data <= 8'h00; 
        10'b0100110011: data <= 8'h00; 
        10'b0100110100: data <= 8'h00; 
        10'b0100110101: data <= 8'h00; 
        10'b0100110110: data <= 8'h00; 
        10'b0100110111: data <= 8'h00; 
        10'b0100111000: data <= 8'h00; 
        10'b0100111001: data <= 8'h00; 
        10'b0100111010: data <= 8'h00; 
        10'b0100111011: data <= 8'h00; 
        10'b0100111100: data <= 8'h00; 
        10'b0100111101: data <= 8'h00; 
        10'b0100111110: data <= 8'hff; 
        10'b0100111111: data <= 8'hff; 
        10'b0101000000: data <= 8'h00; 
        10'b0101000001: data <= 8'h01; 
        10'b0101000010: data <= 8'h02; 
        10'b0101000011: data <= 8'h02; 
        10'b0101000100: data <= 8'h01; 
        10'b0101000101: data <= 8'h00; 
        10'b0101000110: data <= 8'h00; 
        10'b0101000111: data <= 8'h00; 
        10'b0101001000: data <= 8'hff; 
        10'b0101001001: data <= 8'h00; 
        10'b0101001010: data <= 8'h00; 
        10'b0101001011: data <= 8'h00; 
        10'b0101001100: data <= 8'h00; 
        10'b0101001101: data <= 8'h00; 
        10'b0101001110: data <= 8'h00; 
        10'b0101001111: data <= 8'h00; 
        10'b0101010000: data <= 8'h00; 
        10'b0101010001: data <= 8'h00; 
        10'b0101010010: data <= 8'h00; 
        10'b0101010011: data <= 8'h00; 
        10'b0101010100: data <= 8'h00; 
        10'b0101010101: data <= 8'h00; 
        10'b0101010110: data <= 8'h00; 
        10'b0101010111: data <= 8'h00; 
        10'b0101011000: data <= 8'h00; 
        10'b0101011001: data <= 8'h00; 
        10'b0101011010: data <= 8'hff; 
        10'b0101011011: data <= 8'hff; 
        10'b0101011100: data <= 8'h00; 
        10'b0101011101: data <= 8'h01; 
        10'b0101011110: data <= 8'h03; 
        10'b0101011111: data <= 8'h02; 
        10'b0101100000: data <= 8'h00; 
        10'b0101100001: data <= 8'h00; 
        10'b0101100010: data <= 8'h00; 
        10'b0101100011: data <= 8'hff; 
        10'b0101100100: data <= 8'h00; 
        10'b0101100101: data <= 8'h00; 
        10'b0101100110: data <= 8'h00; 
        10'b0101100111: data <= 8'h00; 
        10'b0101101000: data <= 8'h00; 
        10'b0101101001: data <= 8'h00; 
        10'b0101101010: data <= 8'h00; 
        10'b0101101011: data <= 8'h00; 
        10'b0101101100: data <= 8'h00; 
        10'b0101101101: data <= 8'h00; 
        10'b0101101110: data <= 8'h00; 
        10'b0101101111: data <= 8'h00; 
        10'b0101110000: data <= 8'h00; 
        10'b0101110001: data <= 8'h00; 
        10'b0101110010: data <= 8'h00; 
        10'b0101110011: data <= 8'h00; 
        10'b0101110100: data <= 8'h00; 
        10'b0101110101: data <= 8'hff; 
        10'b0101110110: data <= 8'hfe; 
        10'b0101110111: data <= 8'hfe; 
        10'b0101111000: data <= 8'h00; 
        10'b0101111001: data <= 8'h01; 
        10'b0101111010: data <= 8'h02; 
        10'b0101111011: data <= 8'h01; 
        10'b0101111100: data <= 8'h00; 
        10'b0101111101: data <= 8'h00; 
        10'b0101111110: data <= 8'hff; 
        10'b0101111111: data <= 8'hff; 
        10'b0110000000: data <= 8'h00; 
        10'b0110000001: data <= 8'h00; 
        10'b0110000010: data <= 8'h00; 
        10'b0110000011: data <= 8'h00; 
        10'b0110000100: data <= 8'h00; 
        10'b0110000101: data <= 8'h00; 
        10'b0110000110: data <= 8'h00; 
        10'b0110000111: data <= 8'h00; 
        10'b0110001000: data <= 8'h00; 
        10'b0110001001: data <= 8'h00; 
        10'b0110001010: data <= 8'h00; 
        10'b0110001011: data <= 8'h00; 
        10'b0110001100: data <= 8'h00; 
        10'b0110001101: data <= 8'h00; 
        10'b0110001110: data <= 8'h00; 
        10'b0110001111: data <= 8'h00; 
        10'b0110010000: data <= 8'hff; 
        10'b0110010001: data <= 8'hff; 
        10'b0110010010: data <= 8'hfe; 
        10'b0110010011: data <= 8'hff; 
        10'b0110010100: data <= 8'h00; 
        10'b0110010101: data <= 8'h01; 
        10'b0110010110: data <= 8'h02; 
        10'b0110010111: data <= 8'h01; 
        10'b0110011000: data <= 8'h00; 
        10'b0110011001: data <= 8'hff; 
        10'b0110011010: data <= 8'hff; 
        10'b0110011011: data <= 8'hff; 
        10'b0110011100: data <= 8'h00; 
        10'b0110011101: data <= 8'h00; 
        10'b0110011110: data <= 8'h00; 
        10'b0110011111: data <= 8'h00; 
        10'b0110100000: data <= 8'h00; 
        10'b0110100001: data <= 8'h00; 
        10'b0110100010: data <= 8'h00; 
        10'b0110100011: data <= 8'h00; 
        10'b0110100100: data <= 8'h00; 
        10'b0110100101: data <= 8'h00; 
        10'b0110100110: data <= 8'h00; 
        10'b0110100111: data <= 8'h00; 
        10'b0110101000: data <= 8'h00; 
        10'b0110101001: data <= 8'h00; 
        10'b0110101010: data <= 8'h00; 
        10'b0110101011: data <= 8'h00; 
        10'b0110101100: data <= 8'h00; 
        10'b0110101101: data <= 8'hff; 
        10'b0110101110: data <= 8'hff; 
        10'b0110101111: data <= 8'h00; 
        10'b0110110000: data <= 8'h00; 
        10'b0110110001: data <= 8'h01; 
        10'b0110110010: data <= 8'h02; 
        10'b0110110011: data <= 8'h01; 
        10'b0110110100: data <= 8'h00; 
        10'b0110110101: data <= 8'hff; 
        10'b0110110110: data <= 8'hff; 
        10'b0110110111: data <= 8'hff; 
        10'b0110111000: data <= 8'h00; 
        10'b0110111001: data <= 8'h00; 
        10'b0110111010: data <= 8'h00; 
        10'b0110111011: data <= 8'h00; 
        10'b0110111100: data <= 8'h00; 
        10'b0110111101: data <= 8'h00; 
        10'b0110111110: data <= 8'h00; 
        10'b0110111111: data <= 8'h00; 
        10'b0111000000: data <= 8'h00; 
        10'b0111000001: data <= 8'h00; 
        10'b0111000010: data <= 8'h00; 
        10'b0111000011: data <= 8'h00; 
        10'b0111000100: data <= 8'h00; 
        10'b0111000101: data <= 8'h00; 
        10'b0111000110: data <= 8'h00; 
        10'b0111000111: data <= 8'h00; 
        10'b0111001000: data <= 8'hff; 
        10'b0111001001: data <= 8'h00; 
        10'b0111001010: data <= 8'h00; 
        10'b0111001011: data <= 8'h00; 
        10'b0111001100: data <= 8'h00; 
        10'b0111001101: data <= 8'h02; 
        10'b0111001110: data <= 8'h02; 
        10'b0111001111: data <= 8'h00; 
        10'b0111010000: data <= 8'hff; 
        10'b0111010001: data <= 8'hff; 
        10'b0111010010: data <= 8'hff; 
        10'b0111010011: data <= 8'hff; 
        10'b0111010100: data <= 8'hff; 
        10'b0111010101: data <= 8'h00; 
        10'b0111010110: data <= 8'h00; 
        10'b0111010111: data <= 8'h00; 
        10'b0111011000: data <= 8'h00; 
        10'b0111011001: data <= 8'h00; 
        10'b0111011010: data <= 8'h00; 
        10'b0111011011: data <= 8'h00; 
        10'b0111011100: data <= 8'h00; 
        10'b0111011101: data <= 8'h00; 
        10'b0111011110: data <= 8'h00; 
        10'b0111011111: data <= 8'h00; 
        10'b0111100000: data <= 8'h00; 
        10'b0111100001: data <= 8'h00; 
        10'b0111100010: data <= 8'hff; 
        10'b0111100011: data <= 8'hff; 
        10'b0111100100: data <= 8'h00; 
        10'b0111100101: data <= 8'h00; 
        10'b0111100110: data <= 8'h00; 
        10'b0111100111: data <= 8'h00; 
        10'b0111101000: data <= 8'h01; 
        10'b0111101001: data <= 8'h02; 
        10'b0111101010: data <= 8'h02; 
        10'b0111101011: data <= 8'h00; 
        10'b0111101100: data <= 8'hff; 
        10'b0111101101: data <= 8'hff; 
        10'b0111101110: data <= 8'hff; 
        10'b0111101111: data <= 8'hff; 
        10'b0111110000: data <= 8'h00; 
        10'b0111110001: data <= 8'h00; 
        10'b0111110010: data <= 8'h00; 
        10'b0111110011: data <= 8'h00; 
        10'b0111110100: data <= 8'h00; 
        10'b0111110101: data <= 8'h00; 
        10'b0111110110: data <= 8'h00; 
        10'b0111110111: data <= 8'h00; 
        10'b0111111000: data <= 8'h00; 
        10'b0111111001: data <= 8'h00; 
        10'b0111111010: data <= 8'h00; 
        10'b0111111011: data <= 8'h00; 
        10'b0111111100: data <= 8'h00; 
        10'b0111111101: data <= 8'h00; 
        10'b0111111110: data <= 8'hff; 
        10'b0111111111: data <= 8'hff; 
        10'b1000000000: data <= 8'h00; 
        10'b1000000001: data <= 8'h00; 
        10'b1000000010: data <= 8'h00; 
        10'b1000000011: data <= 8'h00; 
        10'b1000000100: data <= 8'h01; 
        10'b1000000101: data <= 8'h01; 
        10'b1000000110: data <= 8'h01; 
        10'b1000000111: data <= 8'hff; 
        10'b1000001000: data <= 8'hff; 
        10'b1000001001: data <= 8'hff; 
        10'b1000001010: data <= 8'hff; 
        10'b1000001011: data <= 8'hff; 
        10'b1000001100: data <= 8'h00; 
        10'b1000001101: data <= 8'h00; 
        10'b1000001110: data <= 8'h00; 
        10'b1000001111: data <= 8'h00; 
        10'b1000010000: data <= 8'h00; 
        10'b1000010001: data <= 8'h00; 
        10'b1000010010: data <= 8'h00; 
        10'b1000010011: data <= 8'h00; 
        10'b1000010100: data <= 8'h00; 
        10'b1000010101: data <= 8'h00; 
        10'b1000010110: data <= 8'h00; 
        10'b1000010111: data <= 8'h00; 
        10'b1000011000: data <= 8'h00; 
        10'b1000011001: data <= 8'h00; 
        10'b1000011010: data <= 8'hff; 
        10'b1000011011: data <= 8'hff; 
        10'b1000011100: data <= 8'h00; 
        10'b1000011101: data <= 8'h00; 
        10'b1000011110: data <= 8'h00; 
        10'b1000011111: data <= 8'h00; 
        10'b1000100000: data <= 8'h00; 
        10'b1000100001: data <= 8'h01; 
        10'b1000100010: data <= 8'h00; 
        10'b1000100011: data <= 8'hff; 
        10'b1000100100: data <= 8'h00; 
        10'b1000100101: data <= 8'h00; 
        10'b1000100110: data <= 8'h00; 
        10'b1000100111: data <= 8'h00; 
        10'b1000101000: data <= 8'hff; 
        10'b1000101001: data <= 8'h00; 
        10'b1000101010: data <= 8'h00; 
        10'b1000101011: data <= 8'h00; 
        10'b1000101100: data <= 8'h00; 
        10'b1000101101: data <= 8'h00; 
        10'b1000101110: data <= 8'h00; 
        10'b1000101111: data <= 8'h00; 
        10'b1000110000: data <= 8'h00; 
        10'b1000110001: data <= 8'h00; 
        10'b1000110010: data <= 8'h00; 
        10'b1000110011: data <= 8'h00; 
        10'b1000110100: data <= 8'h00; 
        10'b1000110101: data <= 8'h00; 
        10'b1000110110: data <= 8'h00; 
        10'b1000110111: data <= 8'h00; 
        10'b1000111000: data <= 8'h00; 
        10'b1000111001: data <= 8'h00; 
        10'b1000111010: data <= 8'h00; 
        10'b1000111011: data <= 8'h00; 
        10'b1000111100: data <= 8'h00; 
        10'b1000111101: data <= 8'h00; 
        10'b1000111110: data <= 8'h00; 
        10'b1000111111: data <= 8'h00; 
        10'b1001000000: data <= 8'h00; 
        10'b1001000001: data <= 8'h00; 
        10'b1001000010: data <= 8'h00; 
        10'b1001000011: data <= 8'h00; 
        10'b1001000100: data <= 8'hff; 
        10'b1001000101: data <= 8'h00; 
        10'b1001000110: data <= 8'h00; 
        10'b1001000111: data <= 8'h00; 
        10'b1001001000: data <= 8'h00; 
        10'b1001001001: data <= 8'h00; 
        10'b1001001010: data <= 8'h00; 
        10'b1001001011: data <= 8'h00; 
        10'b1001001100: data <= 8'h00; 
        10'b1001001101: data <= 8'h00; 
        10'b1001001110: data <= 8'h00; 
        10'b1001001111: data <= 8'h00; 
        10'b1001010000: data <= 8'h00; 
        10'b1001010001: data <= 8'h00; 
        10'b1001010010: data <= 8'h00; 
        10'b1001010011: data <= 8'h00; 
        10'b1001010100: data <= 8'h00; 
        10'b1001010101: data <= 8'h00; 
        10'b1001010110: data <= 8'h00; 
        10'b1001010111: data <= 8'h00; 
        10'b1001011000: data <= 8'hff; 
        10'b1001011001: data <= 8'hff; 
        10'b1001011010: data <= 8'h00; 
        10'b1001011011: data <= 8'h00; 
        10'b1001011100: data <= 8'h00; 
        10'b1001011101: data <= 8'h00; 
        10'b1001011110: data <= 8'h00; 
        10'b1001011111: data <= 8'h00; 
        10'b1001100000: data <= 8'h00; 
        10'b1001100001: data <= 8'h00; 
        10'b1001100010: data <= 8'h00; 
        10'b1001100011: data <= 8'h00; 
        10'b1001100100: data <= 8'h00; 
        10'b1001100101: data <= 8'h00; 
        10'b1001100110: data <= 8'h00; 
        10'b1001100111: data <= 8'h00; 
        10'b1001101000: data <= 8'h00; 
        10'b1001101001: data <= 8'h00; 
        10'b1001101010: data <= 8'h00; 
        10'b1001101011: data <= 8'h00; 
        10'b1001101100: data <= 8'h00; 
        10'b1001101101: data <= 8'h01; 
        10'b1001101110: data <= 8'h01; 
        10'b1001101111: data <= 8'h01; 
        10'b1001110000: data <= 8'h00; 
        10'b1001110001: data <= 8'h00; 
        10'b1001110010: data <= 8'h00; 
        10'b1001110011: data <= 8'hff; 
        10'b1001110100: data <= 8'hff; 
        10'b1001110101: data <= 8'hff; 
        10'b1001110110: data <= 8'h00; 
        10'b1001110111: data <= 8'h00; 
        10'b1001111000: data <= 8'h01; 
        10'b1001111001: data <= 8'h01; 
        10'b1001111010: data <= 8'h01; 
        10'b1001111011: data <= 8'h00; 
        10'b1001111100: data <= 8'h00; 
        10'b1001111101: data <= 8'h00; 
        10'b1001111110: data <= 8'h00; 
        10'b1001111111: data <= 8'h00; 
        10'b1010000000: data <= 8'h00; 
        10'b1010000001: data <= 8'h00; 
        10'b1010000010: data <= 8'h00; 
        10'b1010000011: data <= 8'h00; 
        10'b1010000100: data <= 8'h00; 
        10'b1010000101: data <= 8'h00; 
        10'b1010000110: data <= 8'h00; 
        10'b1010000111: data <= 8'h00; 
        10'b1010001000: data <= 8'h00; 
        10'b1010001001: data <= 8'h01; 
        10'b1010001010: data <= 8'h01; 
        10'b1010001011: data <= 8'h00; 
        10'b1010001100: data <= 8'h00; 
        10'b1010001101: data <= 8'h00; 
        10'b1010001110: data <= 8'h00; 
        10'b1010001111: data <= 8'h00; 
        10'b1010010000: data <= 8'h00; 
        10'b1010010001: data <= 8'h00; 
        10'b1010010010: data <= 8'h00; 
        10'b1010010011: data <= 8'h00; 
        10'b1010010100: data <= 8'h01; 
        10'b1010010101: data <= 8'h01; 
        10'b1010010110: data <= 8'h01; 
        10'b1010010111: data <= 8'h00; 
        10'b1010011000: data <= 8'h00; 
        10'b1010011001: data <= 8'h00; 
        10'b1010011010: data <= 8'h00; 
        10'b1010011011: data <= 8'h00; 
        10'b1010011100: data <= 8'h00; 
        10'b1010011101: data <= 8'h00; 
        10'b1010011110: data <= 8'h00; 
        10'b1010011111: data <= 8'h00; 
        10'b1010100000: data <= 8'h00; 
        10'b1010100001: data <= 8'h00; 
        10'b1010100010: data <= 8'h00; 
        10'b1010100011: data <= 8'h00; 
        10'b1010100100: data <= 8'h00; 
        10'b1010100101: data <= 8'h00; 
        10'b1010100110: data <= 8'h00; 
        10'b1010100111: data <= 8'h00; 
        10'b1010101000: data <= 8'hff; 
        10'b1010101001: data <= 8'hff; 
        10'b1010101010: data <= 8'hff; 
        10'b1010101011: data <= 8'hff; 
        10'b1010101100: data <= 8'hff; 
        10'b1010101101: data <= 8'hff; 
        10'b1010101110: data <= 8'hff; 
        10'b1010101111: data <= 8'hff; 
        10'b1010110000: data <= 8'h00; 
        10'b1010110001: data <= 8'h00; 
        10'b1010110010: data <= 8'h00; 
        10'b1010110011: data <= 8'h00; 
        10'b1010110100: data <= 8'h00; 
        10'b1010110101: data <= 8'h00; 
        10'b1010110110: data <= 8'h00; 
        10'b1010110111: data <= 8'h00; 
        10'b1010111000: data <= 8'h00; 
        10'b1010111001: data <= 8'h00; 
        10'b1010111010: data <= 8'h00; 
        10'b1010111011: data <= 8'h00; 
        10'b1010111100: data <= 8'h00; 
        10'b1010111101: data <= 8'h00; 
        10'b1010111110: data <= 8'h00; 
        10'b1010111111: data <= 8'h00; 
        10'b1011000000: data <= 8'h00; 
        10'b1011000001: data <= 8'h00; 
        10'b1011000010: data <= 8'h00; 
        10'b1011000011: data <= 8'h00; 
        10'b1011000100: data <= 8'h00; 
        10'b1011000101: data <= 8'h00; 
        10'b1011000110: data <= 8'h00; 
        10'b1011000111: data <= 8'hff; 
        10'b1011001000: data <= 8'h00; 
        10'b1011001001: data <= 8'hff; 
        10'b1011001010: data <= 8'h00; 
        10'b1011001011: data <= 8'h00; 
        10'b1011001100: data <= 8'h00; 
        10'b1011001101: data <= 8'h00; 
        10'b1011001110: data <= 8'h00; 
        10'b1011001111: data <= 8'h00; 
        10'b1011010000: data <= 8'h00; 
        10'b1011010001: data <= 8'h00; 
        10'b1011010010: data <= 8'h00; 
        10'b1011010011: data <= 8'h00; 
        10'b1011010100: data <= 8'h00; 
        10'b1011010101: data <= 8'h00; 
        10'b1011010110: data <= 8'h00; 
        10'b1011010111: data <= 8'h00; 
        10'b1011011000: data <= 8'h00; 
        10'b1011011001: data <= 8'h00; 
        10'b1011011010: data <= 8'h00; 
        10'b1011011011: data <= 8'h00; 
        10'b1011011100: data <= 8'h00; 
        10'b1011011101: data <= 8'h00; 
        10'b1011011110: data <= 8'h00; 
        10'b1011011111: data <= 8'h00; 
        10'b1011100000: data <= 8'h00; 
        10'b1011100001: data <= 8'h00; 
        10'b1011100010: data <= 8'h00; 
        10'b1011100011: data <= 8'h00; 
        10'b1011100100: data <= 8'h00; 
        10'b1011100101: data <= 8'h00; 
        10'b1011100110: data <= 8'h00; 
        10'b1011100111: data <= 8'h00; 
        10'b1011101000: data <= 8'h00; 
        10'b1011101001: data <= 8'h00; 
        10'b1011101010: data <= 8'h00; 
        10'b1011101011: data <= 8'h00; 
        10'b1011101100: data <= 8'h00; 
        10'b1011101101: data <= 8'h00; 
        10'b1011101110: data <= 8'h00; 
        10'b1011101111: data <= 8'h00; 
        10'b1011110000: data <= 8'h00; 
        10'b1011110001: data <= 8'h00; 
        10'b1011110010: data <= 8'h00; 
        10'b1011110011: data <= 8'h00; 
        10'b1011110100: data <= 8'h00; 
        10'b1011110101: data <= 8'h00; 
        10'b1011110110: data <= 8'h00; 
        10'b1011110111: data <= 8'h00; 
        10'b1011111000: data <= 8'h00; 
        10'b1011111001: data <= 8'h00; 
        10'b1011111010: data <= 8'h00; 
        10'b1011111011: data <= 8'h00; 
        10'b1011111100: data <= 8'h00; 
        10'b1011111101: data <= 8'h00; 
        10'b1011111110: data <= 8'h00; 
        10'b1011111111: data <= 8'h00; 
        10'b1100000000: data <= 8'h00; 
        10'b1100000001: data <= 8'h00; 
        10'b1100000010: data <= 8'h00; 
        10'b1100000011: data <= 8'h00; 
        10'b1100000100: data <= 8'h00; 
        10'b1100000101: data <= 8'h00; 
        10'b1100000110: data <= 8'h00; 
        10'b1100000111: data <= 8'h00; 
        10'b1100001000: data <= 8'h00; 
        10'b1100001001: data <= 8'h00; 
        10'b1100001010: data <= 8'h00; 
        10'b1100001011: data <= 8'h00; 
        10'b1100001100: data <= 8'h00; 
        10'b1100001101: data <= 8'h00; 
        10'b1100001110: data <= 8'h00; 
        10'b1100001111: data <= 8'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 3) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 9'h000; 
        10'b0000000001: data <= 9'h000; 
        10'b0000000010: data <= 9'h000; 
        10'b0000000011: data <= 9'h000; 
        10'b0000000100: data <= 9'h000; 
        10'b0000000101: data <= 9'h000; 
        10'b0000000110: data <= 9'h000; 
        10'b0000000111: data <= 9'h000; 
        10'b0000001000: data <= 9'h000; 
        10'b0000001001: data <= 9'h000; 
        10'b0000001010: data <= 9'h000; 
        10'b0000001011: data <= 9'h000; 
        10'b0000001100: data <= 9'h000; 
        10'b0000001101: data <= 9'h001; 
        10'b0000001110: data <= 9'h000; 
        10'b0000001111: data <= 9'h000; 
        10'b0000010000: data <= 9'h000; 
        10'b0000010001: data <= 9'h000; 
        10'b0000010010: data <= 9'h001; 
        10'b0000010011: data <= 9'h001; 
        10'b0000010100: data <= 9'h000; 
        10'b0000010101: data <= 9'h000; 
        10'b0000010110: data <= 9'h000; 
        10'b0000010111: data <= 9'h001; 
        10'b0000011000: data <= 9'h000; 
        10'b0000011001: data <= 9'h001; 
        10'b0000011010: data <= 9'h000; 
        10'b0000011011: data <= 9'h000; 
        10'b0000011100: data <= 9'h000; 
        10'b0000011101: data <= 9'h001; 
        10'b0000011110: data <= 9'h000; 
        10'b0000011111: data <= 9'h000; 
        10'b0000100000: data <= 9'h000; 
        10'b0000100001: data <= 9'h000; 
        10'b0000100010: data <= 9'h000; 
        10'b0000100011: data <= 9'h000; 
        10'b0000100100: data <= 9'h000; 
        10'b0000100101: data <= 9'h000; 
        10'b0000100110: data <= 9'h000; 
        10'b0000100111: data <= 9'h000; 
        10'b0000101000: data <= 9'h000; 
        10'b0000101001: data <= 9'h000; 
        10'b0000101010: data <= 9'h001; 
        10'b0000101011: data <= 9'h000; 
        10'b0000101100: data <= 9'h000; 
        10'b0000101101: data <= 9'h001; 
        10'b0000101110: data <= 9'h000; 
        10'b0000101111: data <= 9'h000; 
        10'b0000110000: data <= 9'h001; 
        10'b0000110001: data <= 9'h001; 
        10'b0000110010: data <= 9'h000; 
        10'b0000110011: data <= 9'h001; 
        10'b0000110100: data <= 9'h001; 
        10'b0000110101: data <= 9'h000; 
        10'b0000110110: data <= 9'h001; 
        10'b0000110111: data <= 9'h000; 
        10'b0000111000: data <= 9'h001; 
        10'b0000111001: data <= 9'h000; 
        10'b0000111010: data <= 9'h001; 
        10'b0000111011: data <= 9'h000; 
        10'b0000111100: data <= 9'h000; 
        10'b0000111101: data <= 9'h000; 
        10'b0000111110: data <= 9'h000; 
        10'b0000111111: data <= 9'h000; 
        10'b0001000000: data <= 9'h000; 
        10'b0001000001: data <= 9'h000; 
        10'b0001000010: data <= 9'h000; 
        10'b0001000011: data <= 9'h000; 
        10'b0001000100: data <= 9'h000; 
        10'b0001000101: data <= 9'h000; 
        10'b0001000110: data <= 9'h000; 
        10'b0001000111: data <= 9'h000; 
        10'b0001001000: data <= 9'h000; 
        10'b0001001001: data <= 9'h000; 
        10'b0001001010: data <= 9'h000; 
        10'b0001001011: data <= 9'h000; 
        10'b0001001100: data <= 9'h000; 
        10'b0001001101: data <= 9'h000; 
        10'b0001001110: data <= 9'h001; 
        10'b0001001111: data <= 9'h000; 
        10'b0001010000: data <= 9'h000; 
        10'b0001010001: data <= 9'h000; 
        10'b0001010010: data <= 9'h000; 
        10'b0001010011: data <= 9'h000; 
        10'b0001010100: data <= 9'h000; 
        10'b0001010101: data <= 9'h000; 
        10'b0001010110: data <= 9'h000; 
        10'b0001010111: data <= 9'h000; 
        10'b0001011000: data <= 9'h001; 
        10'b0001011001: data <= 9'h000; 
        10'b0001011010: data <= 9'h000; 
        10'b0001011011: data <= 9'h001; 
        10'b0001011100: data <= 9'h000; 
        10'b0001011101: data <= 9'h000; 
        10'b0001011110: data <= 9'h000; 
        10'b0001011111: data <= 9'h000; 
        10'b0001100000: data <= 9'h000; 
        10'b0001100001: data <= 9'h000; 
        10'b0001100010: data <= 9'h000; 
        10'b0001100011: data <= 9'h000; 
        10'b0001100100: data <= 9'h000; 
        10'b0001100101: data <= 9'h000; 
        10'b0001100110: data <= 9'h000; 
        10'b0001100111: data <= 9'h000; 
        10'b0001101000: data <= 9'h000; 
        10'b0001101001: data <= 9'h000; 
        10'b0001101010: data <= 9'h000; 
        10'b0001101011: data <= 9'h000; 
        10'b0001101100: data <= 9'h000; 
        10'b0001101101: data <= 9'h001; 
        10'b0001101110: data <= 9'h000; 
        10'b0001101111: data <= 9'h001; 
        10'b0001110000: data <= 9'h000; 
        10'b0001110001: data <= 9'h000; 
        10'b0001110010: data <= 9'h001; 
        10'b0001110011: data <= 9'h001; 
        10'b0001110100: data <= 9'h000; 
        10'b0001110101: data <= 9'h000; 
        10'b0001110110: data <= 9'h001; 
        10'b0001110111: data <= 9'h000; 
        10'b0001111000: data <= 9'h000; 
        10'b0001111001: data <= 9'h1ff; 
        10'b0001111010: data <= 9'h000; 
        10'b0001111011: data <= 9'h000; 
        10'b0001111100: data <= 9'h000; 
        10'b0001111101: data <= 9'h001; 
        10'b0001111110: data <= 9'h001; 
        10'b0001111111: data <= 9'h001; 
        10'b0010000000: data <= 9'h000; 
        10'b0010000001: data <= 9'h000; 
        10'b0010000010: data <= 9'h000; 
        10'b0010000011: data <= 9'h000; 
        10'b0010000100: data <= 9'h001; 
        10'b0010000101: data <= 9'h001; 
        10'b0010000110: data <= 9'h001; 
        10'b0010000111: data <= 9'h001; 
        10'b0010001000: data <= 9'h000; 
        10'b0010001001: data <= 9'h000; 
        10'b0010001010: data <= 9'h000; 
        10'b0010001011: data <= 9'h000; 
        10'b0010001100: data <= 9'h000; 
        10'b0010001101: data <= 9'h000; 
        10'b0010001110: data <= 9'h000; 
        10'b0010001111: data <= 9'h000; 
        10'b0010010000: data <= 9'h000; 
        10'b0010010001: data <= 9'h000; 
        10'b0010010010: data <= 9'h000; 
        10'b0010010011: data <= 9'h000; 
        10'b0010010100: data <= 9'h1ff; 
        10'b0010010101: data <= 9'h1ff; 
        10'b0010010110: data <= 9'h1ff; 
        10'b0010010111: data <= 9'h000; 
        10'b0010011000: data <= 9'h000; 
        10'b0010011001: data <= 9'h000; 
        10'b0010011010: data <= 9'h001; 
        10'b0010011011: data <= 9'h001; 
        10'b0010011100: data <= 9'h000; 
        10'b0010011101: data <= 9'h1ff; 
        10'b0010011110: data <= 9'h000; 
        10'b0010011111: data <= 9'h000; 
        10'b0010100000: data <= 9'h001; 
        10'b0010100001: data <= 9'h001; 
        10'b0010100010: data <= 9'h002; 
        10'b0010100011: data <= 9'h001; 
        10'b0010100100: data <= 9'h001; 
        10'b0010100101: data <= 9'h000; 
        10'b0010100110: data <= 9'h000; 
        10'b0010100111: data <= 9'h000; 
        10'b0010101000: data <= 9'h000; 
        10'b0010101001: data <= 9'h000; 
        10'b0010101010: data <= 9'h000; 
        10'b0010101011: data <= 9'h000; 
        10'b0010101100: data <= 9'h000; 
        10'b0010101101: data <= 9'h000; 
        10'b0010101110: data <= 9'h1ff; 
        10'b0010101111: data <= 9'h1ff; 
        10'b0010110000: data <= 9'h1ff; 
        10'b0010110001: data <= 9'h1fe; 
        10'b0010110010: data <= 9'h1ff; 
        10'b0010110011: data <= 9'h000; 
        10'b0010110100: data <= 9'h000; 
        10'b0010110101: data <= 9'h1ff; 
        10'b0010110110: data <= 9'h000; 
        10'b0010110111: data <= 9'h1ff; 
        10'b0010111000: data <= 9'h1ff; 
        10'b0010111001: data <= 9'h1ff; 
        10'b0010111010: data <= 9'h1ff; 
        10'b0010111011: data <= 9'h000; 
        10'b0010111100: data <= 9'h001; 
        10'b0010111101: data <= 9'h001; 
        10'b0010111110: data <= 9'h001; 
        10'b0010111111: data <= 9'h001; 
        10'b0011000000: data <= 9'h000; 
        10'b0011000001: data <= 9'h000; 
        10'b0011000010: data <= 9'h000; 
        10'b0011000011: data <= 9'h000; 
        10'b0011000100: data <= 9'h000; 
        10'b0011000101: data <= 9'h000; 
        10'b0011000110: data <= 9'h000; 
        10'b0011000111: data <= 9'h000; 
        10'b0011001000: data <= 9'h000; 
        10'b0011001001: data <= 9'h000; 
        10'b0011001010: data <= 9'h1ff; 
        10'b0011001011: data <= 9'h1ff; 
        10'b0011001100: data <= 9'h1fe; 
        10'b0011001101: data <= 9'h1fe; 
        10'b0011001110: data <= 9'h1fe; 
        10'b0011001111: data <= 9'h1ff; 
        10'b0011010000: data <= 9'h1ff; 
        10'b0011010001: data <= 9'h1ff; 
        10'b0011010010: data <= 9'h1ff; 
        10'b0011010011: data <= 9'h1fe; 
        10'b0011010100: data <= 9'h1fe; 
        10'b0011010101: data <= 9'h1ff; 
        10'b0011010110: data <= 9'h1ff; 
        10'b0011010111: data <= 9'h000; 
        10'b0011011000: data <= 9'h000; 
        10'b0011011001: data <= 9'h000; 
        10'b0011011010: data <= 9'h000; 
        10'b0011011011: data <= 9'h1ff; 
        10'b0011011100: data <= 9'h1ff; 
        10'b0011011101: data <= 9'h000; 
        10'b0011011110: data <= 9'h000; 
        10'b0011011111: data <= 9'h000; 
        10'b0011100000: data <= 9'h000; 
        10'b0011100001: data <= 9'h000; 
        10'b0011100010: data <= 9'h000; 
        10'b0011100011: data <= 9'h001; 
        10'b0011100100: data <= 9'h000; 
        10'b0011100101: data <= 9'h000; 
        10'b0011100110: data <= 9'h1ff; 
        10'b0011100111: data <= 9'h1ff; 
        10'b0011101000: data <= 9'h1fe; 
        10'b0011101001: data <= 9'h1fe; 
        10'b0011101010: data <= 9'h1fe; 
        10'b0011101011: data <= 9'h1ff; 
        10'b0011101100: data <= 9'h1ff; 
        10'b0011101101: data <= 9'h1ff; 
        10'b0011101110: data <= 9'h1ff; 
        10'b0011101111: data <= 9'h000; 
        10'b0011110000: data <= 9'h1ff; 
        10'b0011110001: data <= 9'h000; 
        10'b0011110010: data <= 9'h000; 
        10'b0011110011: data <= 9'h000; 
        10'b0011110100: data <= 9'h1ff; 
        10'b0011110101: data <= 9'h1ff; 
        10'b0011110110: data <= 9'h1ff; 
        10'b0011110111: data <= 9'h1fe; 
        10'b0011111000: data <= 9'h1ff; 
        10'b0011111001: data <= 9'h000; 
        10'b0011111010: data <= 9'h000; 
        10'b0011111011: data <= 9'h001; 
        10'b0011111100: data <= 9'h001; 
        10'b0011111101: data <= 9'h000; 
        10'b0011111110: data <= 9'h000; 
        10'b0011111111: data <= 9'h000; 
        10'b0100000000: data <= 9'h000; 
        10'b0100000001: data <= 9'h000; 
        10'b0100000010: data <= 9'h1ff; 
        10'b0100000011: data <= 9'h1ff; 
        10'b0100000100: data <= 9'h1fe; 
        10'b0100000101: data <= 9'h1fe; 
        10'b0100000110: data <= 9'h1fe; 
        10'b0100000111: data <= 9'h1ff; 
        10'b0100001000: data <= 9'h1ff; 
        10'b0100001001: data <= 9'h000; 
        10'b0100001010: data <= 9'h001; 
        10'b0100001011: data <= 9'h002; 
        10'b0100001100: data <= 9'h001; 
        10'b0100001101: data <= 9'h000; 
        10'b0100001110: data <= 9'h000; 
        10'b0100001111: data <= 9'h1ff; 
        10'b0100010000: data <= 9'h1fe; 
        10'b0100010001: data <= 9'h1fe; 
        10'b0100010010: data <= 9'h1fe; 
        10'b0100010011: data <= 9'h1fe; 
        10'b0100010100: data <= 9'h1ff; 
        10'b0100010101: data <= 9'h000; 
        10'b0100010110: data <= 9'h000; 
        10'b0100010111: data <= 9'h000; 
        10'b0100011000: data <= 9'h001; 
        10'b0100011001: data <= 9'h001; 
        10'b0100011010: data <= 9'h001; 
        10'b0100011011: data <= 9'h000; 
        10'b0100011100: data <= 9'h000; 
        10'b0100011101: data <= 9'h000; 
        10'b0100011110: data <= 9'h1ff; 
        10'b0100011111: data <= 9'h000; 
        10'b0100100000: data <= 9'h1ff; 
        10'b0100100001: data <= 9'h1ff; 
        10'b0100100010: data <= 9'h1ff; 
        10'b0100100011: data <= 9'h1ff; 
        10'b0100100100: data <= 9'h000; 
        10'b0100100101: data <= 9'h001; 
        10'b0100100110: data <= 9'h004; 
        10'b0100100111: data <= 9'h004; 
        10'b0100101000: data <= 9'h002; 
        10'b0100101001: data <= 9'h000; 
        10'b0100101010: data <= 9'h1ff; 
        10'b0100101011: data <= 9'h1ff; 
        10'b0100101100: data <= 9'h1fe; 
        10'b0100101101: data <= 9'h1fe; 
        10'b0100101110: data <= 9'h1ff; 
        10'b0100101111: data <= 9'h1ff; 
        10'b0100110000: data <= 9'h000; 
        10'b0100110001: data <= 9'h000; 
        10'b0100110010: data <= 9'h001; 
        10'b0100110011: data <= 9'h000; 
        10'b0100110100: data <= 9'h000; 
        10'b0100110101: data <= 9'h000; 
        10'b0100110110: data <= 9'h000; 
        10'b0100110111: data <= 9'h000; 
        10'b0100111000: data <= 9'h000; 
        10'b0100111001: data <= 9'h000; 
        10'b0100111010: data <= 9'h000; 
        10'b0100111011: data <= 9'h1ff; 
        10'b0100111100: data <= 9'h000; 
        10'b0100111101: data <= 9'h1ff; 
        10'b0100111110: data <= 9'h1ff; 
        10'b0100111111: data <= 9'h1fe; 
        10'b0101000000: data <= 9'h000; 
        10'b0101000001: data <= 9'h002; 
        10'b0101000010: data <= 9'h005; 
        10'b0101000011: data <= 9'h005; 
        10'b0101000100: data <= 9'h002; 
        10'b0101000101: data <= 9'h000; 
        10'b0101000110: data <= 9'h000; 
        10'b0101000111: data <= 9'h1ff; 
        10'b0101001000: data <= 9'h1ff; 
        10'b0101001001: data <= 9'h1ff; 
        10'b0101001010: data <= 9'h1ff; 
        10'b0101001011: data <= 9'h000; 
        10'b0101001100: data <= 9'h000; 
        10'b0101001101: data <= 9'h000; 
        10'b0101001110: data <= 9'h001; 
        10'b0101001111: data <= 9'h000; 
        10'b0101010000: data <= 9'h000; 
        10'b0101010001: data <= 9'h001; 
        10'b0101010010: data <= 9'h000; 
        10'b0101010011: data <= 9'h000; 
        10'b0101010100: data <= 9'h001; 
        10'b0101010101: data <= 9'h000; 
        10'b0101010110: data <= 9'h000; 
        10'b0101010111: data <= 9'h000; 
        10'b0101011000: data <= 9'h1ff; 
        10'b0101011001: data <= 9'h1ff; 
        10'b0101011010: data <= 9'h1fe; 
        10'b0101011011: data <= 9'h1fd; 
        10'b0101011100: data <= 9'h000; 
        10'b0101011101: data <= 9'h002; 
        10'b0101011110: data <= 9'h005; 
        10'b0101011111: data <= 9'h004; 
        10'b0101100000: data <= 9'h001; 
        10'b0101100001: data <= 9'h000; 
        10'b0101100010: data <= 9'h000; 
        10'b0101100011: data <= 9'h1ff; 
        10'b0101100100: data <= 9'h1ff; 
        10'b0101100101: data <= 9'h000; 
        10'b0101100110: data <= 9'h000; 
        10'b0101100111: data <= 9'h000; 
        10'b0101101000: data <= 9'h000; 
        10'b0101101001: data <= 9'h001; 
        10'b0101101010: data <= 9'h000; 
        10'b0101101011: data <= 9'h000; 
        10'b0101101100: data <= 9'h000; 
        10'b0101101101: data <= 9'h000; 
        10'b0101101110: data <= 9'h000; 
        10'b0101101111: data <= 9'h000; 
        10'b0101110000: data <= 9'h001; 
        10'b0101110001: data <= 9'h000; 
        10'b0101110010: data <= 9'h000; 
        10'b0101110011: data <= 9'h000; 
        10'b0101110100: data <= 9'h000; 
        10'b0101110101: data <= 9'h1fe; 
        10'b0101110110: data <= 9'h1fd; 
        10'b0101110111: data <= 9'h1fd; 
        10'b0101111000: data <= 9'h000; 
        10'b0101111001: data <= 9'h002; 
        10'b0101111010: data <= 9'h004; 
        10'b0101111011: data <= 9'h003; 
        10'b0101111100: data <= 9'h001; 
        10'b0101111101: data <= 9'h000; 
        10'b0101111110: data <= 9'h1ff; 
        10'b0101111111: data <= 9'h1ff; 
        10'b0110000000: data <= 9'h1ff; 
        10'b0110000001: data <= 9'h000; 
        10'b0110000010: data <= 9'h000; 
        10'b0110000011: data <= 9'h000; 
        10'b0110000100: data <= 9'h000; 
        10'b0110000101: data <= 9'h000; 
        10'b0110000110: data <= 9'h001; 
        10'b0110000111: data <= 9'h000; 
        10'b0110001000: data <= 9'h000; 
        10'b0110001001: data <= 9'h001; 
        10'b0110001010: data <= 9'h000; 
        10'b0110001011: data <= 9'h000; 
        10'b0110001100: data <= 9'h000; 
        10'b0110001101: data <= 9'h000; 
        10'b0110001110: data <= 9'h000; 
        10'b0110001111: data <= 9'h000; 
        10'b0110010000: data <= 9'h1ff; 
        10'b0110010001: data <= 9'h1fe; 
        10'b0110010010: data <= 9'h1fd; 
        10'b0110010011: data <= 9'h1fe; 
        10'b0110010100: data <= 9'h000; 
        10'b0110010101: data <= 9'h002; 
        10'b0110010110: data <= 9'h004; 
        10'b0110010111: data <= 9'h002; 
        10'b0110011000: data <= 9'h001; 
        10'b0110011001: data <= 9'h1ff; 
        10'b0110011010: data <= 9'h1fe; 
        10'b0110011011: data <= 9'h1ff; 
        10'b0110011100: data <= 9'h1ff; 
        10'b0110011101: data <= 9'h000; 
        10'b0110011110: data <= 9'h000; 
        10'b0110011111: data <= 9'h000; 
        10'b0110100000: data <= 9'h000; 
        10'b0110100001: data <= 9'h000; 
        10'b0110100010: data <= 9'h000; 
        10'b0110100011: data <= 9'h000; 
        10'b0110100100: data <= 9'h001; 
        10'b0110100101: data <= 9'h000; 
        10'b0110100110: data <= 9'h000; 
        10'b0110100111: data <= 9'h000; 
        10'b0110101000: data <= 9'h000; 
        10'b0110101001: data <= 9'h000; 
        10'b0110101010: data <= 9'h000; 
        10'b0110101011: data <= 9'h000; 
        10'b0110101100: data <= 9'h1ff; 
        10'b0110101101: data <= 9'h1fe; 
        10'b0110101110: data <= 9'h1fe; 
        10'b0110101111: data <= 9'h1ff; 
        10'b0110110000: data <= 9'h001; 
        10'b0110110001: data <= 9'h002; 
        10'b0110110010: data <= 9'h004; 
        10'b0110110011: data <= 9'h001; 
        10'b0110110100: data <= 9'h000; 
        10'b0110110101: data <= 9'h1fd; 
        10'b0110110110: data <= 9'h1fe; 
        10'b0110110111: data <= 9'h1ff; 
        10'b0110111000: data <= 9'h1ff; 
        10'b0110111001: data <= 9'h1ff; 
        10'b0110111010: data <= 9'h000; 
        10'b0110111011: data <= 9'h000; 
        10'b0110111100: data <= 9'h000; 
        10'b0110111101: data <= 9'h000; 
        10'b0110111110: data <= 9'h001; 
        10'b0110111111: data <= 9'h000; 
        10'b0111000000: data <= 9'h001; 
        10'b0111000001: data <= 9'h000; 
        10'b0111000010: data <= 9'h001; 
        10'b0111000011: data <= 9'h000; 
        10'b0111000100: data <= 9'h000; 
        10'b0111000101: data <= 9'h000; 
        10'b0111000110: data <= 9'h1ff; 
        10'b0111000111: data <= 9'h1ff; 
        10'b0111001000: data <= 9'h1ff; 
        10'b0111001001: data <= 9'h1ff; 
        10'b0111001010: data <= 9'h1ff; 
        10'b0111001011: data <= 9'h000; 
        10'b0111001100: data <= 9'h000; 
        10'b0111001101: data <= 9'h003; 
        10'b0111001110: data <= 9'h004; 
        10'b0111001111: data <= 9'h000; 
        10'b0111010000: data <= 9'h1ff; 
        10'b0111010001: data <= 9'h1fd; 
        10'b0111010010: data <= 9'h1fe; 
        10'b0111010011: data <= 9'h1ff; 
        10'b0111010100: data <= 9'h1ff; 
        10'b0111010101: data <= 9'h000; 
        10'b0111010110: data <= 9'h000; 
        10'b0111010111: data <= 9'h000; 
        10'b0111011000: data <= 9'h000; 
        10'b0111011001: data <= 9'h000; 
        10'b0111011010: data <= 9'h000; 
        10'b0111011011: data <= 9'h000; 
        10'b0111011100: data <= 9'h000; 
        10'b0111011101: data <= 9'h001; 
        10'b0111011110: data <= 9'h000; 
        10'b0111011111: data <= 9'h001; 
        10'b0111100000: data <= 9'h000; 
        10'b0111100001: data <= 9'h000; 
        10'b0111100010: data <= 9'h1ff; 
        10'b0111100011: data <= 9'h1ff; 
        10'b0111100100: data <= 9'h1ff; 
        10'b0111100101: data <= 9'h1ff; 
        10'b0111100110: data <= 9'h000; 
        10'b0111100111: data <= 9'h000; 
        10'b0111101000: data <= 9'h001; 
        10'b0111101001: data <= 9'h004; 
        10'b0111101010: data <= 9'h003; 
        10'b0111101011: data <= 9'h1ff; 
        10'b0111101100: data <= 9'h1fe; 
        10'b0111101101: data <= 9'h1fd; 
        10'b0111101110: data <= 9'h1fe; 
        10'b0111101111: data <= 9'h1ff; 
        10'b0111110000: data <= 9'h1ff; 
        10'b0111110001: data <= 9'h000; 
        10'b0111110010: data <= 9'h000; 
        10'b0111110011: data <= 9'h000; 
        10'b0111110100: data <= 9'h000; 
        10'b0111110101: data <= 9'h000; 
        10'b0111110110: data <= 9'h000; 
        10'b0111110111: data <= 9'h000; 
        10'b0111111000: data <= 9'h000; 
        10'b0111111001: data <= 9'h000; 
        10'b0111111010: data <= 9'h000; 
        10'b0111111011: data <= 9'h000; 
        10'b0111111100: data <= 9'h000; 
        10'b0111111101: data <= 9'h000; 
        10'b0111111110: data <= 9'h1ff; 
        10'b0111111111: data <= 9'h1ff; 
        10'b1000000000: data <= 9'h000; 
        10'b1000000001: data <= 9'h000; 
        10'b1000000010: data <= 9'h000; 
        10'b1000000011: data <= 9'h001; 
        10'b1000000100: data <= 9'h002; 
        10'b1000000101: data <= 9'h003; 
        10'b1000000110: data <= 9'h002; 
        10'b1000000111: data <= 9'h1ff; 
        10'b1000001000: data <= 9'h1fe; 
        10'b1000001001: data <= 9'h1fe; 
        10'b1000001010: data <= 9'h1fe; 
        10'b1000001011: data <= 9'h1ff; 
        10'b1000001100: data <= 9'h000; 
        10'b1000001101: data <= 9'h1ff; 
        10'b1000001110: data <= 9'h000; 
        10'b1000001111: data <= 9'h1ff; 
        10'b1000010000: data <= 9'h000; 
        10'b1000010001: data <= 9'h000; 
        10'b1000010010: data <= 9'h001; 
        10'b1000010011: data <= 9'h001; 
        10'b1000010100: data <= 9'h001; 
        10'b1000010101: data <= 9'h000; 
        10'b1000010110: data <= 9'h000; 
        10'b1000010111: data <= 9'h000; 
        10'b1000011000: data <= 9'h000; 
        10'b1000011001: data <= 9'h1ff; 
        10'b1000011010: data <= 9'h1fe; 
        10'b1000011011: data <= 9'h1ff; 
        10'b1000011100: data <= 9'h000; 
        10'b1000011101: data <= 9'h000; 
        10'b1000011110: data <= 9'h000; 
        10'b1000011111: data <= 9'h000; 
        10'b1000100000: data <= 9'h000; 
        10'b1000100001: data <= 9'h001; 
        10'b1000100010: data <= 9'h000; 
        10'b1000100011: data <= 9'h1ff; 
        10'b1000100100: data <= 9'h1ff; 
        10'b1000100101: data <= 9'h1ff; 
        10'b1000100110: data <= 9'h1ff; 
        10'b1000100111: data <= 9'h1ff; 
        10'b1000101000: data <= 9'h1ff; 
        10'b1000101001: data <= 9'h1ff; 
        10'b1000101010: data <= 9'h1ff; 
        10'b1000101011: data <= 9'h000; 
        10'b1000101100: data <= 9'h000; 
        10'b1000101101: data <= 9'h000; 
        10'b1000101110: data <= 9'h000; 
        10'b1000101111: data <= 9'h000; 
        10'b1000110000: data <= 9'h000; 
        10'b1000110001: data <= 9'h001; 
        10'b1000110010: data <= 9'h000; 
        10'b1000110011: data <= 9'h000; 
        10'b1000110100: data <= 9'h000; 
        10'b1000110101: data <= 9'h1ff; 
        10'b1000110110: data <= 9'h000; 
        10'b1000110111: data <= 9'h000; 
        10'b1000111000: data <= 9'h000; 
        10'b1000111001: data <= 9'h000; 
        10'b1000111010: data <= 9'h000; 
        10'b1000111011: data <= 9'h000; 
        10'b1000111100: data <= 9'h1ff; 
        10'b1000111101: data <= 9'h000; 
        10'b1000111110: data <= 9'h000; 
        10'b1000111111: data <= 9'h000; 
        10'b1001000000: data <= 9'h001; 
        10'b1001000001: data <= 9'h000; 
        10'b1001000010: data <= 9'h000; 
        10'b1001000011: data <= 9'h1ff; 
        10'b1001000100: data <= 9'h1ff; 
        10'b1001000101: data <= 9'h1ff; 
        10'b1001000110: data <= 9'h1ff; 
        10'b1001000111: data <= 9'h000; 
        10'b1001001000: data <= 9'h000; 
        10'b1001001001: data <= 9'h000; 
        10'b1001001010: data <= 9'h000; 
        10'b1001001011: data <= 9'h001; 
        10'b1001001100: data <= 9'h000; 
        10'b1001001101: data <= 9'h000; 
        10'b1001001110: data <= 9'h000; 
        10'b1001001111: data <= 9'h000; 
        10'b1001010000: data <= 9'h000; 
        10'b1001010001: data <= 9'h001; 
        10'b1001010010: data <= 9'h001; 
        10'b1001010011: data <= 9'h000; 
        10'b1001010100: data <= 9'h000; 
        10'b1001010101: data <= 9'h000; 
        10'b1001010110: data <= 9'h000; 
        10'b1001010111: data <= 9'h1ff; 
        10'b1001011000: data <= 9'h1ff; 
        10'b1001011001: data <= 9'h1ff; 
        10'b1001011010: data <= 9'h000; 
        10'b1001011011: data <= 9'h000; 
        10'b1001011100: data <= 9'h001; 
        10'b1001011101: data <= 9'h001; 
        10'b1001011110: data <= 9'h001; 
        10'b1001011111: data <= 9'h1ff; 
        10'b1001100000: data <= 9'h1ff; 
        10'b1001100001: data <= 9'h1ff; 
        10'b1001100010: data <= 9'h1ff; 
        10'b1001100011: data <= 9'h000; 
        10'b1001100100: data <= 9'h000; 
        10'b1001100101: data <= 9'h000; 
        10'b1001100110: data <= 9'h000; 
        10'b1001100111: data <= 9'h000; 
        10'b1001101000: data <= 9'h000; 
        10'b1001101001: data <= 9'h000; 
        10'b1001101010: data <= 9'h000; 
        10'b1001101011: data <= 9'h000; 
        10'b1001101100: data <= 9'h001; 
        10'b1001101101: data <= 9'h002; 
        10'b1001101110: data <= 9'h002; 
        10'b1001101111: data <= 9'h001; 
        10'b1001110000: data <= 9'h000; 
        10'b1001110001: data <= 9'h000; 
        10'b1001110010: data <= 9'h000; 
        10'b1001110011: data <= 9'h1fe; 
        10'b1001110100: data <= 9'h1fd; 
        10'b1001110101: data <= 9'h1fe; 
        10'b1001110110: data <= 9'h000; 
        10'b1001110111: data <= 9'h000; 
        10'b1001111000: data <= 9'h002; 
        10'b1001111001: data <= 9'h003; 
        10'b1001111010: data <= 9'h001; 
        10'b1001111011: data <= 9'h000; 
        10'b1001111100: data <= 9'h1ff; 
        10'b1001111101: data <= 9'h000; 
        10'b1001111110: data <= 9'h000; 
        10'b1001111111: data <= 9'h000; 
        10'b1010000000: data <= 9'h000; 
        10'b1010000001: data <= 9'h000; 
        10'b1010000010: data <= 9'h001; 
        10'b1010000011: data <= 9'h000; 
        10'b1010000100: data <= 9'h001; 
        10'b1010000101: data <= 9'h000; 
        10'b1010000110: data <= 9'h000; 
        10'b1010000111: data <= 9'h000; 
        10'b1010001000: data <= 9'h001; 
        10'b1010001001: data <= 9'h002; 
        10'b1010001010: data <= 9'h002; 
        10'b1010001011: data <= 9'h001; 
        10'b1010001100: data <= 9'h000; 
        10'b1010001101: data <= 9'h000; 
        10'b1010001110: data <= 9'h000; 
        10'b1010001111: data <= 9'h1ff; 
        10'b1010010000: data <= 9'h1ff; 
        10'b1010010001: data <= 9'h1ff; 
        10'b1010010010: data <= 9'h1ff; 
        10'b1010010011: data <= 9'h000; 
        10'b1010010100: data <= 9'h002; 
        10'b1010010101: data <= 9'h002; 
        10'b1010010110: data <= 9'h001; 
        10'b1010010111: data <= 9'h000; 
        10'b1010011000: data <= 9'h000; 
        10'b1010011001: data <= 9'h1ff; 
        10'b1010011010: data <= 9'h000; 
        10'b1010011011: data <= 9'h000; 
        10'b1010011100: data <= 9'h000; 
        10'b1010011101: data <= 9'h000; 
        10'b1010011110: data <= 9'h000; 
        10'b1010011111: data <= 9'h000; 
        10'b1010100000: data <= 9'h000; 
        10'b1010100001: data <= 9'h000; 
        10'b1010100010: data <= 9'h000; 
        10'b1010100011: data <= 9'h000; 
        10'b1010100100: data <= 9'h000; 
        10'b1010100101: data <= 9'h001; 
        10'b1010100110: data <= 9'h001; 
        10'b1010100111: data <= 9'h000; 
        10'b1010101000: data <= 9'h1ff; 
        10'b1010101001: data <= 9'h1ff; 
        10'b1010101010: data <= 9'h1fe; 
        10'b1010101011: data <= 9'h1fe; 
        10'b1010101100: data <= 9'h1fe; 
        10'b1010101101: data <= 9'h1ff; 
        10'b1010101110: data <= 9'h1ff; 
        10'b1010101111: data <= 9'h1ff; 
        10'b1010110000: data <= 9'h000; 
        10'b1010110001: data <= 9'h000; 
        10'b1010110010: data <= 9'h000; 
        10'b1010110011: data <= 9'h000; 
        10'b1010110100: data <= 9'h000; 
        10'b1010110101: data <= 9'h000; 
        10'b1010110110: data <= 9'h000; 
        10'b1010110111: data <= 9'h000; 
        10'b1010111000: data <= 9'h000; 
        10'b1010111001: data <= 9'h000; 
        10'b1010111010: data <= 9'h000; 
        10'b1010111011: data <= 9'h000; 
        10'b1010111100: data <= 9'h001; 
        10'b1010111101: data <= 9'h000; 
        10'b1010111110: data <= 9'h000; 
        10'b1010111111: data <= 9'h000; 
        10'b1011000000: data <= 9'h000; 
        10'b1011000001: data <= 9'h000; 
        10'b1011000010: data <= 9'h000; 
        10'b1011000011: data <= 9'h000; 
        10'b1011000100: data <= 9'h000; 
        10'b1011000101: data <= 9'h000; 
        10'b1011000110: data <= 9'h1ff; 
        10'b1011000111: data <= 9'h1ff; 
        10'b1011001000: data <= 9'h1ff; 
        10'b1011001001: data <= 9'h1ff; 
        10'b1011001010: data <= 9'h1ff; 
        10'b1011001011: data <= 9'h1ff; 
        10'b1011001100: data <= 9'h1ff; 
        10'b1011001101: data <= 9'h000; 
        10'b1011001110: data <= 9'h000; 
        10'b1011001111: data <= 9'h000; 
        10'b1011010000: data <= 9'h000; 
        10'b1011010001: data <= 9'h000; 
        10'b1011010010: data <= 9'h000; 
        10'b1011010011: data <= 9'h001; 
        10'b1011010100: data <= 9'h000; 
        10'b1011010101: data <= 9'h000; 
        10'b1011010110: data <= 9'h000; 
        10'b1011010111: data <= 9'h000; 
        10'b1011011000: data <= 9'h000; 
        10'b1011011001: data <= 9'h000; 
        10'b1011011010: data <= 9'h000; 
        10'b1011011011: data <= 9'h000; 
        10'b1011011100: data <= 9'h000; 
        10'b1011011101: data <= 9'h001; 
        10'b1011011110: data <= 9'h000; 
        10'b1011011111: data <= 9'h000; 
        10'b1011100000: data <= 9'h000; 
        10'b1011100001: data <= 9'h000; 
        10'b1011100010: data <= 9'h000; 
        10'b1011100011: data <= 9'h000; 
        10'b1011100100: data <= 9'h000; 
        10'b1011100101: data <= 9'h000; 
        10'b1011100110: data <= 9'h000; 
        10'b1011100111: data <= 9'h000; 
        10'b1011101000: data <= 9'h000; 
        10'b1011101001: data <= 9'h001; 
        10'b1011101010: data <= 9'h000; 
        10'b1011101011: data <= 9'h000; 
        10'b1011101100: data <= 9'h000; 
        10'b1011101101: data <= 9'h000; 
        10'b1011101110: data <= 9'h000; 
        10'b1011101111: data <= 9'h000; 
        10'b1011110000: data <= 9'h000; 
        10'b1011110001: data <= 9'h000; 
        10'b1011110010: data <= 9'h001; 
        10'b1011110011: data <= 9'h000; 
        10'b1011110100: data <= 9'h000; 
        10'b1011110101: data <= 9'h001; 
        10'b1011110110: data <= 9'h000; 
        10'b1011110111: data <= 9'h000; 
        10'b1011111000: data <= 9'h001; 
        10'b1011111001: data <= 9'h000; 
        10'b1011111010: data <= 9'h001; 
        10'b1011111011: data <= 9'h000; 
        10'b1011111100: data <= 9'h001; 
        10'b1011111101: data <= 9'h000; 
        10'b1011111110: data <= 9'h000; 
        10'b1011111111: data <= 9'h000; 
        10'b1100000000: data <= 9'h000; 
        10'b1100000001: data <= 9'h000; 
        10'b1100000010: data <= 9'h001; 
        10'b1100000011: data <= 9'h000; 
        10'b1100000100: data <= 9'h000; 
        10'b1100000101: data <= 9'h000; 
        10'b1100000110: data <= 9'h000; 
        10'b1100000111: data <= 9'h000; 
        10'b1100001000: data <= 9'h000; 
        10'b1100001001: data <= 9'h000; 
        10'b1100001010: data <= 9'h000; 
        10'b1100001011: data <= 9'h000; 
        10'b1100001100: data <= 9'h001; 
        10'b1100001101: data <= 9'h001; 
        10'b1100001110: data <= 9'h001; 
        10'b1100001111: data <= 9'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 4) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 10'h001; 
        10'b0000000001: data <= 10'h000; 
        10'b0000000010: data <= 10'h001; 
        10'b0000000011: data <= 10'h000; 
        10'b0000000100: data <= 10'h001; 
        10'b0000000101: data <= 10'h001; 
        10'b0000000110: data <= 10'h001; 
        10'b0000000111: data <= 10'h000; 
        10'b0000001000: data <= 10'h001; 
        10'b0000001001: data <= 10'h000; 
        10'b0000001010: data <= 10'h001; 
        10'b0000001011: data <= 10'h001; 
        10'b0000001100: data <= 10'h001; 
        10'b0000001101: data <= 10'h001; 
        10'b0000001110: data <= 10'h001; 
        10'b0000001111: data <= 10'h001; 
        10'b0000010000: data <= 10'h001; 
        10'b0000010001: data <= 10'h000; 
        10'b0000010010: data <= 10'h001; 
        10'b0000010011: data <= 10'h001; 
        10'b0000010100: data <= 10'h001; 
        10'b0000010101: data <= 10'h001; 
        10'b0000010110: data <= 10'h001; 
        10'b0000010111: data <= 10'h001; 
        10'b0000011000: data <= 10'h000; 
        10'b0000011001: data <= 10'h001; 
        10'b0000011010: data <= 10'h001; 
        10'b0000011011: data <= 10'h001; 
        10'b0000011100: data <= 10'h000; 
        10'b0000011101: data <= 10'h001; 
        10'b0000011110: data <= 10'h000; 
        10'b0000011111: data <= 10'h001; 
        10'b0000100000: data <= 10'h001; 
        10'b0000100001: data <= 10'h000; 
        10'b0000100010: data <= 10'h000; 
        10'b0000100011: data <= 10'h001; 
        10'b0000100100: data <= 10'h001; 
        10'b0000100101: data <= 10'h001; 
        10'b0000100110: data <= 10'h001; 
        10'b0000100111: data <= 10'h001; 
        10'b0000101000: data <= 10'h001; 
        10'b0000101001: data <= 10'h001; 
        10'b0000101010: data <= 10'h001; 
        10'b0000101011: data <= 10'h001; 
        10'b0000101100: data <= 10'h001; 
        10'b0000101101: data <= 10'h001; 
        10'b0000101110: data <= 10'h001; 
        10'b0000101111: data <= 10'h000; 
        10'b0000110000: data <= 10'h001; 
        10'b0000110001: data <= 10'h001; 
        10'b0000110010: data <= 10'h000; 
        10'b0000110011: data <= 10'h001; 
        10'b0000110100: data <= 10'h001; 
        10'b0000110101: data <= 10'h001; 
        10'b0000110110: data <= 10'h001; 
        10'b0000110111: data <= 10'h001; 
        10'b0000111000: data <= 10'h001; 
        10'b0000111001: data <= 10'h001; 
        10'b0000111010: data <= 10'h001; 
        10'b0000111011: data <= 10'h000; 
        10'b0000111100: data <= 10'h000; 
        10'b0000111101: data <= 10'h001; 
        10'b0000111110: data <= 10'h001; 
        10'b0000111111: data <= 10'h001; 
        10'b0001000000: data <= 10'h000; 
        10'b0001000001: data <= 10'h001; 
        10'b0001000010: data <= 10'h000; 
        10'b0001000011: data <= 10'h000; 
        10'b0001000100: data <= 10'h000; 
        10'b0001000101: data <= 10'h000; 
        10'b0001000110: data <= 10'h001; 
        10'b0001000111: data <= 10'h001; 
        10'b0001001000: data <= 10'h001; 
        10'b0001001001: data <= 10'h000; 
        10'b0001001010: data <= 10'h001; 
        10'b0001001011: data <= 10'h000; 
        10'b0001001100: data <= 10'h001; 
        10'b0001001101: data <= 10'h000; 
        10'b0001001110: data <= 10'h001; 
        10'b0001001111: data <= 10'h001; 
        10'b0001010000: data <= 10'h001; 
        10'b0001010001: data <= 10'h000; 
        10'b0001010010: data <= 10'h001; 
        10'b0001010011: data <= 10'h001; 
        10'b0001010100: data <= 10'h000; 
        10'b0001010101: data <= 10'h000; 
        10'b0001010110: data <= 10'h001; 
        10'b0001010111: data <= 10'h001; 
        10'b0001011000: data <= 10'h001; 
        10'b0001011001: data <= 10'h001; 
        10'b0001011010: data <= 10'h000; 
        10'b0001011011: data <= 10'h001; 
        10'b0001011100: data <= 10'h000; 
        10'b0001011101: data <= 10'h000; 
        10'b0001011110: data <= 10'h000; 
        10'b0001011111: data <= 10'h3ff; 
        10'b0001100000: data <= 10'h000; 
        10'b0001100001: data <= 10'h000; 
        10'b0001100010: data <= 10'h000; 
        10'b0001100011: data <= 10'h001; 
        10'b0001100100: data <= 10'h000; 
        10'b0001100101: data <= 10'h000; 
        10'b0001100110: data <= 10'h000; 
        10'b0001100111: data <= 10'h3ff; 
        10'b0001101000: data <= 10'h000; 
        10'b0001101001: data <= 10'h000; 
        10'b0001101010: data <= 10'h001; 
        10'b0001101011: data <= 10'h001; 
        10'b0001101100: data <= 10'h000; 
        10'b0001101101: data <= 10'h001; 
        10'b0001101110: data <= 10'h000; 
        10'b0001101111: data <= 10'h001; 
        10'b0001110000: data <= 10'h001; 
        10'b0001110001: data <= 10'h001; 
        10'b0001110010: data <= 10'h001; 
        10'b0001110011: data <= 10'h001; 
        10'b0001110100: data <= 10'h000; 
        10'b0001110101: data <= 10'h000; 
        10'b0001110110: data <= 10'h001; 
        10'b0001110111: data <= 10'h001; 
        10'b0001111000: data <= 10'h000; 
        10'b0001111001: data <= 10'h3ff; 
        10'b0001111010: data <= 10'h000; 
        10'b0001111011: data <= 10'h000; 
        10'b0001111100: data <= 10'h001; 
        10'b0001111101: data <= 10'h001; 
        10'b0001111110: data <= 10'h001; 
        10'b0001111111: data <= 10'h002; 
        10'b0010000000: data <= 10'h001; 
        10'b0010000001: data <= 10'h3ff; 
        10'b0010000010: data <= 10'h3ff; 
        10'b0010000011: data <= 10'h000; 
        10'b0010000100: data <= 10'h001; 
        10'b0010000101: data <= 10'h002; 
        10'b0010000110: data <= 10'h002; 
        10'b0010000111: data <= 10'h002; 
        10'b0010001000: data <= 10'h001; 
        10'b0010001001: data <= 10'h000; 
        10'b0010001010: data <= 10'h000; 
        10'b0010001011: data <= 10'h000; 
        10'b0010001100: data <= 10'h000; 
        10'b0010001101: data <= 10'h001; 
        10'b0010001110: data <= 10'h000; 
        10'b0010001111: data <= 10'h001; 
        10'b0010010000: data <= 10'h000; 
        10'b0010010001: data <= 10'h001; 
        10'b0010010010: data <= 10'h000; 
        10'b0010010011: data <= 10'h000; 
        10'b0010010100: data <= 10'h3fe; 
        10'b0010010101: data <= 10'h3fe; 
        10'b0010010110: data <= 10'h3ff; 
        10'b0010010111: data <= 10'h000; 
        10'b0010011000: data <= 10'h001; 
        10'b0010011001: data <= 10'h001; 
        10'b0010011010: data <= 10'h002; 
        10'b0010011011: data <= 10'h001; 
        10'b0010011100: data <= 10'h001; 
        10'b0010011101: data <= 10'h3ff; 
        10'b0010011110: data <= 10'h000; 
        10'b0010011111: data <= 10'h000; 
        10'b0010100000: data <= 10'h001; 
        10'b0010100001: data <= 10'h002; 
        10'b0010100010: data <= 10'h003; 
        10'b0010100011: data <= 10'h002; 
        10'b0010100100: data <= 10'h002; 
        10'b0010100101: data <= 10'h000; 
        10'b0010100110: data <= 10'h000; 
        10'b0010100111: data <= 10'h000; 
        10'b0010101000: data <= 10'h000; 
        10'b0010101001: data <= 10'h001; 
        10'b0010101010: data <= 10'h000; 
        10'b0010101011: data <= 10'h001; 
        10'b0010101100: data <= 10'h000; 
        10'b0010101101: data <= 10'h000; 
        10'b0010101110: data <= 10'h3ff; 
        10'b0010101111: data <= 10'h3ff; 
        10'b0010110000: data <= 10'h3fd; 
        10'b0010110001: data <= 10'h3fd; 
        10'b0010110010: data <= 10'h3fe; 
        10'b0010110011: data <= 10'h000; 
        10'b0010110100: data <= 10'h3ff; 
        10'b0010110101: data <= 10'h3ff; 
        10'b0010110110: data <= 10'h000; 
        10'b0010110111: data <= 10'h3fe; 
        10'b0010111000: data <= 10'h3fd; 
        10'b0010111001: data <= 10'h3fd; 
        10'b0010111010: data <= 10'h3ff; 
        10'b0010111011: data <= 10'h3ff; 
        10'b0010111100: data <= 10'h001; 
        10'b0010111101: data <= 10'h002; 
        10'b0010111110: data <= 10'h002; 
        10'b0010111111: data <= 10'h002; 
        10'b0011000000: data <= 10'h000; 
        10'b0011000001: data <= 10'h000; 
        10'b0011000010: data <= 10'h000; 
        10'b0011000011: data <= 10'h001; 
        10'b0011000100: data <= 10'h000; 
        10'b0011000101: data <= 10'h000; 
        10'b0011000110: data <= 10'h000; 
        10'b0011000111: data <= 10'h000; 
        10'b0011001000: data <= 10'h001; 
        10'b0011001001: data <= 10'h000; 
        10'b0011001010: data <= 10'h3ff; 
        10'b0011001011: data <= 10'h3fe; 
        10'b0011001100: data <= 10'h3fc; 
        10'b0011001101: data <= 10'h3fb; 
        10'b0011001110: data <= 10'h3fd; 
        10'b0011001111: data <= 10'h3ff; 
        10'b0011010000: data <= 10'h3ff; 
        10'b0011010001: data <= 10'h3fe; 
        10'b0011010010: data <= 10'h3fe; 
        10'b0011010011: data <= 10'h3fc; 
        10'b0011010100: data <= 10'h3fd; 
        10'b0011010101: data <= 10'h3fd; 
        10'b0011010110: data <= 10'h3fd; 
        10'b0011010111: data <= 10'h000; 
        10'b0011011000: data <= 10'h001; 
        10'b0011011001: data <= 10'h000; 
        10'b0011011010: data <= 10'h000; 
        10'b0011011011: data <= 10'h3ff; 
        10'b0011011100: data <= 10'h3ff; 
        10'b0011011101: data <= 10'h3ff; 
        10'b0011011110: data <= 10'h000; 
        10'b0011011111: data <= 10'h001; 
        10'b0011100000: data <= 10'h001; 
        10'b0011100001: data <= 10'h000; 
        10'b0011100010: data <= 10'h000; 
        10'b0011100011: data <= 10'h001; 
        10'b0011100100: data <= 10'h000; 
        10'b0011100101: data <= 10'h000; 
        10'b0011100110: data <= 10'h3ff; 
        10'b0011100111: data <= 10'h3fe; 
        10'b0011101000: data <= 10'h3fc; 
        10'b0011101001: data <= 10'h3fb; 
        10'b0011101010: data <= 10'h3fb; 
        10'b0011101011: data <= 10'h3fe; 
        10'b0011101100: data <= 10'h3ff; 
        10'b0011101101: data <= 10'h3ff; 
        10'b0011101110: data <= 10'h3ff; 
        10'b0011101111: data <= 10'h000; 
        10'b0011110000: data <= 10'h3fe; 
        10'b0011110001: data <= 10'h3ff; 
        10'b0011110010: data <= 10'h000; 
        10'b0011110011: data <= 10'h000; 
        10'b0011110100: data <= 10'h3ff; 
        10'b0011110101: data <= 10'h3ff; 
        10'b0011110110: data <= 10'h3fe; 
        10'b0011110111: data <= 10'h3fd; 
        10'b0011111000: data <= 10'h3fe; 
        10'b0011111001: data <= 10'h3ff; 
        10'b0011111010: data <= 10'h001; 
        10'b0011111011: data <= 10'h001; 
        10'b0011111100: data <= 10'h001; 
        10'b0011111101: data <= 10'h000; 
        10'b0011111110: data <= 10'h000; 
        10'b0011111111: data <= 10'h000; 
        10'b0100000000: data <= 10'h000; 
        10'b0100000001: data <= 10'h000; 
        10'b0100000010: data <= 10'h3fe; 
        10'b0100000011: data <= 10'h3fe; 
        10'b0100000100: data <= 10'h3fd; 
        10'b0100000101: data <= 10'h3fb; 
        10'b0100000110: data <= 10'h3fc; 
        10'b0100000111: data <= 10'h3fe; 
        10'b0100001000: data <= 10'h3ff; 
        10'b0100001001: data <= 10'h001; 
        10'b0100001010: data <= 10'h003; 
        10'b0100001011: data <= 10'h004; 
        10'b0100001100: data <= 10'h002; 
        10'b0100001101: data <= 10'h000; 
        10'b0100001110: data <= 10'h3ff; 
        10'b0100001111: data <= 10'h3fd; 
        10'b0100010000: data <= 10'h3fc; 
        10'b0100010001: data <= 10'h3fc; 
        10'b0100010010: data <= 10'h3fc; 
        10'b0100010011: data <= 10'h3fc; 
        10'b0100010100: data <= 10'h3fe; 
        10'b0100010101: data <= 10'h000; 
        10'b0100010110: data <= 10'h001; 
        10'b0100010111: data <= 10'h001; 
        10'b0100011000: data <= 10'h001; 
        10'b0100011001: data <= 10'h001; 
        10'b0100011010: data <= 10'h001; 
        10'b0100011011: data <= 10'h000; 
        10'b0100011100: data <= 10'h001; 
        10'b0100011101: data <= 10'h3ff; 
        10'b0100011110: data <= 10'h3fe; 
        10'b0100011111: data <= 10'h3ff; 
        10'b0100100000: data <= 10'h3fe; 
        10'b0100100001: data <= 10'h3fe; 
        10'b0100100010: data <= 10'h3fe; 
        10'b0100100011: data <= 10'h3ff; 
        10'b0100100100: data <= 10'h3ff; 
        10'b0100100101: data <= 10'h002; 
        10'b0100100110: data <= 10'h008; 
        10'b0100100111: data <= 10'h008; 
        10'b0100101000: data <= 10'h004; 
        10'b0100101001: data <= 10'h000; 
        10'b0100101010: data <= 10'h3fe; 
        10'b0100101011: data <= 10'h3fd; 
        10'b0100101100: data <= 10'h3fd; 
        10'b0100101101: data <= 10'h3fd; 
        10'b0100101110: data <= 10'h3fd; 
        10'b0100101111: data <= 10'h3fe; 
        10'b0100110000: data <= 10'h3ff; 
        10'b0100110001: data <= 10'h000; 
        10'b0100110010: data <= 10'h001; 
        10'b0100110011: data <= 10'h000; 
        10'b0100110100: data <= 10'h000; 
        10'b0100110101: data <= 10'h000; 
        10'b0100110110: data <= 10'h001; 
        10'b0100110111: data <= 10'h001; 
        10'b0100111000: data <= 10'h000; 
        10'b0100111001: data <= 10'h000; 
        10'b0100111010: data <= 10'h000; 
        10'b0100111011: data <= 10'h3ff; 
        10'b0100111100: data <= 10'h3ff; 
        10'b0100111101: data <= 10'h3ff; 
        10'b0100111110: data <= 10'h3fe; 
        10'b0100111111: data <= 10'h3fd; 
        10'b0101000000: data <= 10'h000; 
        10'b0101000001: data <= 10'h004; 
        10'b0101000010: data <= 10'h009; 
        10'b0101000011: data <= 10'h00a; 
        10'b0101000100: data <= 10'h004; 
        10'b0101000101: data <= 10'h3ff; 
        10'b0101000110: data <= 10'h3ff; 
        10'b0101000111: data <= 10'h3fe; 
        10'b0101001000: data <= 10'h3fe; 
        10'b0101001001: data <= 10'h3fe; 
        10'b0101001010: data <= 10'h3fe; 
        10'b0101001011: data <= 10'h3ff; 
        10'b0101001100: data <= 10'h000; 
        10'b0101001101: data <= 10'h001; 
        10'b0101001110: data <= 10'h001; 
        10'b0101001111: data <= 10'h001; 
        10'b0101010000: data <= 10'h000; 
        10'b0101010001: data <= 10'h001; 
        10'b0101010010: data <= 10'h001; 
        10'b0101010011: data <= 10'h000; 
        10'b0101010100: data <= 10'h001; 
        10'b0101010101: data <= 10'h000; 
        10'b0101010110: data <= 10'h000; 
        10'b0101010111: data <= 10'h000; 
        10'b0101011000: data <= 10'h3ff; 
        10'b0101011001: data <= 10'h3fe; 
        10'b0101011010: data <= 10'h3fc; 
        10'b0101011011: data <= 10'h3fb; 
        10'b0101011100: data <= 10'h000; 
        10'b0101011101: data <= 10'h004; 
        10'b0101011110: data <= 10'h00b; 
        10'b0101011111: data <= 10'h008; 
        10'b0101100000: data <= 10'h001; 
        10'b0101100001: data <= 10'h001; 
        10'b0101100010: data <= 10'h000; 
        10'b0101100011: data <= 10'h3fe; 
        10'b0101100100: data <= 10'h3ff; 
        10'b0101100101: data <= 10'h3ff; 
        10'b0101100110: data <= 10'h000; 
        10'b0101100111: data <= 10'h000; 
        10'b0101101000: data <= 10'h000; 
        10'b0101101001: data <= 10'h001; 
        10'b0101101010: data <= 10'h000; 
        10'b0101101011: data <= 10'h001; 
        10'b0101101100: data <= 10'h000; 
        10'b0101101101: data <= 10'h001; 
        10'b0101101110: data <= 10'h001; 
        10'b0101101111: data <= 10'h001; 
        10'b0101110000: data <= 10'h001; 
        10'b0101110001: data <= 10'h000; 
        10'b0101110010: data <= 10'h000; 
        10'b0101110011: data <= 10'h3ff; 
        10'b0101110100: data <= 10'h3ff; 
        10'b0101110101: data <= 10'h3fd; 
        10'b0101110110: data <= 10'h3fa; 
        10'b0101110111: data <= 10'h3f9; 
        10'b0101111000: data <= 10'h000; 
        10'b0101111001: data <= 10'h003; 
        10'b0101111010: data <= 10'h009; 
        10'b0101111011: data <= 10'h005; 
        10'b0101111100: data <= 10'h001; 
        10'b0101111101: data <= 10'h001; 
        10'b0101111110: data <= 10'h3fe; 
        10'b0101111111: data <= 10'h3fd; 
        10'b0110000000: data <= 10'h3ff; 
        10'b0110000001: data <= 10'h000; 
        10'b0110000010: data <= 10'h000; 
        10'b0110000011: data <= 10'h000; 
        10'b0110000100: data <= 10'h001; 
        10'b0110000101: data <= 10'h001; 
        10'b0110000110: data <= 10'h001; 
        10'b0110000111: data <= 10'h001; 
        10'b0110001000: data <= 10'h001; 
        10'b0110001001: data <= 10'h001; 
        10'b0110001010: data <= 10'h001; 
        10'b0110001011: data <= 10'h001; 
        10'b0110001100: data <= 10'h001; 
        10'b0110001101: data <= 10'h000; 
        10'b0110001110: data <= 10'h000; 
        10'b0110001111: data <= 10'h000; 
        10'b0110010000: data <= 10'h3fe; 
        10'b0110010001: data <= 10'h3fd; 
        10'b0110010010: data <= 10'h3fa; 
        10'b0110010011: data <= 10'h3fb; 
        10'b0110010100: data <= 10'h000; 
        10'b0110010101: data <= 10'h003; 
        10'b0110010110: data <= 10'h008; 
        10'b0110010111: data <= 10'h005; 
        10'b0110011000: data <= 10'h001; 
        10'b0110011001: data <= 10'h3fd; 
        10'b0110011010: data <= 10'h3fc; 
        10'b0110011011: data <= 10'h3fd; 
        10'b0110011100: data <= 10'h3fe; 
        10'b0110011101: data <= 10'h000; 
        10'b0110011110: data <= 10'h3ff; 
        10'b0110011111: data <= 10'h000; 
        10'b0110100000: data <= 10'h001; 
        10'b0110100001: data <= 10'h000; 
        10'b0110100010: data <= 10'h000; 
        10'b0110100011: data <= 10'h001; 
        10'b0110100100: data <= 10'h001; 
        10'b0110100101: data <= 10'h000; 
        10'b0110100110: data <= 10'h001; 
        10'b0110100111: data <= 10'h001; 
        10'b0110101000: data <= 10'h000; 
        10'b0110101001: data <= 10'h001; 
        10'b0110101010: data <= 10'h3ff; 
        10'b0110101011: data <= 10'h3ff; 
        10'b0110101100: data <= 10'h3ff; 
        10'b0110101101: data <= 10'h3fc; 
        10'b0110101110: data <= 10'h3fc; 
        10'b0110101111: data <= 10'h3ff; 
        10'b0110110000: data <= 10'h002; 
        10'b0110110001: data <= 10'h005; 
        10'b0110110010: data <= 10'h008; 
        10'b0110110011: data <= 10'h003; 
        10'b0110110100: data <= 10'h001; 
        10'b0110110101: data <= 10'h3fb; 
        10'b0110110110: data <= 10'h3fb; 
        10'b0110110111: data <= 10'h3fd; 
        10'b0110111000: data <= 10'h3fe; 
        10'b0110111001: data <= 10'h3ff; 
        10'b0110111010: data <= 10'h000; 
        10'b0110111011: data <= 10'h000; 
        10'b0110111100: data <= 10'h000; 
        10'b0110111101: data <= 10'h001; 
        10'b0110111110: data <= 10'h001; 
        10'b0110111111: data <= 10'h000; 
        10'b0111000000: data <= 10'h001; 
        10'b0111000001: data <= 10'h001; 
        10'b0111000010: data <= 10'h001; 
        10'b0111000011: data <= 10'h001; 
        10'b0111000100: data <= 10'h000; 
        10'b0111000101: data <= 10'h000; 
        10'b0111000110: data <= 10'h3ff; 
        10'b0111000111: data <= 10'h3ff; 
        10'b0111001000: data <= 10'h3fd; 
        10'b0111001001: data <= 10'h3fe; 
        10'b0111001010: data <= 10'h3ff; 
        10'b0111001011: data <= 10'h3ff; 
        10'b0111001100: data <= 10'h000; 
        10'b0111001101: data <= 10'h006; 
        10'b0111001110: data <= 10'h008; 
        10'b0111001111: data <= 10'h000; 
        10'b0111010000: data <= 10'h3fe; 
        10'b0111010001: data <= 10'h3fa; 
        10'b0111010010: data <= 10'h3fb; 
        10'b0111010011: data <= 10'h3fd; 
        10'b0111010100: data <= 10'h3fe; 
        10'b0111010101: data <= 10'h3ff; 
        10'b0111010110: data <= 10'h3ff; 
        10'b0111010111: data <= 10'h000; 
        10'b0111011000: data <= 10'h000; 
        10'b0111011001: data <= 10'h000; 
        10'b0111011010: data <= 10'h000; 
        10'b0111011011: data <= 10'h001; 
        10'b0111011100: data <= 10'h000; 
        10'b0111011101: data <= 10'h001; 
        10'b0111011110: data <= 10'h000; 
        10'b0111011111: data <= 10'h001; 
        10'b0111100000: data <= 10'h001; 
        10'b0111100001: data <= 10'h3ff; 
        10'b0111100010: data <= 10'h3fe; 
        10'b0111100011: data <= 10'h3fd; 
        10'b0111100100: data <= 10'h3fe; 
        10'b0111100101: data <= 10'h3ff; 
        10'b0111100110: data <= 10'h001; 
        10'b0111100111: data <= 10'h000; 
        10'b0111101000: data <= 10'h002; 
        10'b0111101001: data <= 10'h007; 
        10'b0111101010: data <= 10'h006; 
        10'b0111101011: data <= 10'h3ff; 
        10'b0111101100: data <= 10'h3fc; 
        10'b0111101101: data <= 10'h3fa; 
        10'b0111101110: data <= 10'h3fb; 
        10'b0111101111: data <= 10'h3fd; 
        10'b0111110000: data <= 10'h3ff; 
        10'b0111110001: data <= 10'h3ff; 
        10'b0111110010: data <= 10'h000; 
        10'b0111110011: data <= 10'h3ff; 
        10'b0111110100: data <= 10'h3ff; 
        10'b0111110101: data <= 10'h000; 
        10'b0111110110: data <= 10'h001; 
        10'b0111110111: data <= 10'h001; 
        10'b0111111000: data <= 10'h001; 
        10'b0111111001: data <= 10'h001; 
        10'b0111111010: data <= 10'h000; 
        10'b0111111011: data <= 10'h001; 
        10'b0111111100: data <= 10'h001; 
        10'b0111111101: data <= 10'h3ff; 
        10'b0111111110: data <= 10'h3fd; 
        10'b0111111111: data <= 10'h3fd; 
        10'b1000000000: data <= 10'h3ff; 
        10'b1000000001: data <= 10'h001; 
        10'b1000000010: data <= 10'h001; 
        10'b1000000011: data <= 10'h001; 
        10'b1000000100: data <= 10'h003; 
        10'b1000000101: data <= 10'h006; 
        10'b1000000110: data <= 10'h004; 
        10'b1000000111: data <= 10'h3fd; 
        10'b1000001000: data <= 10'h3fc; 
        10'b1000001001: data <= 10'h3fc; 
        10'b1000001010: data <= 10'h3fd; 
        10'b1000001011: data <= 10'h3fe; 
        10'b1000001100: data <= 10'h3ff; 
        10'b1000001101: data <= 10'h3fe; 
        10'b1000001110: data <= 10'h3ff; 
        10'b1000001111: data <= 10'h3ff; 
        10'b1000010000: data <= 10'h3ff; 
        10'b1000010001: data <= 10'h001; 
        10'b1000010010: data <= 10'h001; 
        10'b1000010011: data <= 10'h001; 
        10'b1000010100: data <= 10'h001; 
        10'b1000010101: data <= 10'h001; 
        10'b1000010110: data <= 10'h001; 
        10'b1000010111: data <= 10'h001; 
        10'b1000011000: data <= 10'h000; 
        10'b1000011001: data <= 10'h3ff; 
        10'b1000011010: data <= 10'h3fd; 
        10'b1000011011: data <= 10'h3fe; 
        10'b1000011100: data <= 10'h3ff; 
        10'b1000011101: data <= 10'h001; 
        10'b1000011110: data <= 10'h000; 
        10'b1000011111: data <= 10'h000; 
        10'b1000100000: data <= 10'h000; 
        10'b1000100001: data <= 10'h003; 
        10'b1000100010: data <= 10'h001; 
        10'b1000100011: data <= 10'h3fe; 
        10'b1000100100: data <= 10'h3fe; 
        10'b1000100101: data <= 10'h3fe; 
        10'b1000100110: data <= 10'h3fe; 
        10'b1000100111: data <= 10'h3ff; 
        10'b1000101000: data <= 10'h3fe; 
        10'b1000101001: data <= 10'h3fe; 
        10'b1000101010: data <= 10'h3ff; 
        10'b1000101011: data <= 10'h3ff; 
        10'b1000101100: data <= 10'h000; 
        10'b1000101101: data <= 10'h000; 
        10'b1000101110: data <= 10'h000; 
        10'b1000101111: data <= 10'h000; 
        10'b1000110000: data <= 10'h000; 
        10'b1000110001: data <= 10'h001; 
        10'b1000110010: data <= 10'h001; 
        10'b1000110011: data <= 10'h000; 
        10'b1000110100: data <= 10'h000; 
        10'b1000110101: data <= 10'h3ff; 
        10'b1000110110: data <= 10'h000; 
        10'b1000110111: data <= 10'h3ff; 
        10'b1000111000: data <= 10'h000; 
        10'b1000111001: data <= 10'h000; 
        10'b1000111010: data <= 10'h3ff; 
        10'b1000111011: data <= 10'h000; 
        10'b1000111100: data <= 10'h3ff; 
        10'b1000111101: data <= 10'h000; 
        10'b1000111110: data <= 10'h000; 
        10'b1000111111: data <= 10'h000; 
        10'b1001000000: data <= 10'h001; 
        10'b1001000001: data <= 10'h000; 
        10'b1001000010: data <= 10'h000; 
        10'b1001000011: data <= 10'h3fe; 
        10'b1001000100: data <= 10'h3fe; 
        10'b1001000101: data <= 10'h3fe; 
        10'b1001000110: data <= 10'h3fe; 
        10'b1001000111: data <= 10'h000; 
        10'b1001001000: data <= 10'h000; 
        10'b1001001001: data <= 10'h001; 
        10'b1001001010: data <= 10'h000; 
        10'b1001001011: data <= 10'h001; 
        10'b1001001100: data <= 10'h001; 
        10'b1001001101: data <= 10'h000; 
        10'b1001001110: data <= 10'h001; 
        10'b1001001111: data <= 10'h001; 
        10'b1001010000: data <= 10'h001; 
        10'b1001010001: data <= 10'h002; 
        10'b1001010010: data <= 10'h001; 
        10'b1001010011: data <= 10'h001; 
        10'b1001010100: data <= 10'h000; 
        10'b1001010101: data <= 10'h3ff; 
        10'b1001010110: data <= 10'h000; 
        10'b1001010111: data <= 10'h3ff; 
        10'b1001011000: data <= 10'h3fe; 
        10'b1001011001: data <= 10'h3fd; 
        10'b1001011010: data <= 10'h000; 
        10'b1001011011: data <= 10'h001; 
        10'b1001011100: data <= 10'h001; 
        10'b1001011101: data <= 10'h001; 
        10'b1001011110: data <= 10'h001; 
        10'b1001011111: data <= 10'h3fe; 
        10'b1001100000: data <= 10'h3fe; 
        10'b1001100001: data <= 10'h3fe; 
        10'b1001100010: data <= 10'h3ff; 
        10'b1001100011: data <= 10'h3ff; 
        10'b1001100100: data <= 10'h000; 
        10'b1001100101: data <= 10'h001; 
        10'b1001100110: data <= 10'h000; 
        10'b1001100111: data <= 10'h000; 
        10'b1001101000: data <= 10'h001; 
        10'b1001101001: data <= 10'h001; 
        10'b1001101010: data <= 10'h001; 
        10'b1001101011: data <= 10'h000; 
        10'b1001101100: data <= 10'h002; 
        10'b1001101101: data <= 10'h004; 
        10'b1001101110: data <= 10'h004; 
        10'b1001101111: data <= 10'h002; 
        10'b1001110000: data <= 10'h000; 
        10'b1001110001: data <= 10'h000; 
        10'b1001110010: data <= 10'h3ff; 
        10'b1001110011: data <= 10'h3fd; 
        10'b1001110100: data <= 10'h3fa; 
        10'b1001110101: data <= 10'h3fc; 
        10'b1001110110: data <= 10'h000; 
        10'b1001110111: data <= 10'h001; 
        10'b1001111000: data <= 10'h003; 
        10'b1001111001: data <= 10'h005; 
        10'b1001111010: data <= 10'h002; 
        10'b1001111011: data <= 10'h000; 
        10'b1001111100: data <= 10'h3ff; 
        10'b1001111101: data <= 10'h3ff; 
        10'b1001111110: data <= 10'h000; 
        10'b1001111111: data <= 10'h000; 
        10'b1010000000: data <= 10'h000; 
        10'b1010000001: data <= 10'h001; 
        10'b1010000010: data <= 10'h001; 
        10'b1010000011: data <= 10'h001; 
        10'b1010000100: data <= 10'h001; 
        10'b1010000101: data <= 10'h001; 
        10'b1010000110: data <= 10'h001; 
        10'b1010000111: data <= 10'h000; 
        10'b1010001000: data <= 10'h001; 
        10'b1010001001: data <= 10'h003; 
        10'b1010001010: data <= 10'h003; 
        10'b1010001011: data <= 10'h001; 
        10'b1010001100: data <= 10'h000; 
        10'b1010001101: data <= 10'h3ff; 
        10'b1010001110: data <= 10'h3ff; 
        10'b1010001111: data <= 10'h3fe; 
        10'b1010010000: data <= 10'h3ff; 
        10'b1010010001: data <= 10'h3ff; 
        10'b1010010010: data <= 10'h3fe; 
        10'b1010010011: data <= 10'h001; 
        10'b1010010100: data <= 10'h004; 
        10'b1010010101: data <= 10'h005; 
        10'b1010010110: data <= 10'h002; 
        10'b1010010111: data <= 10'h000; 
        10'b1010011000: data <= 10'h3ff; 
        10'b1010011001: data <= 10'h3ff; 
        10'b1010011010: data <= 10'h000; 
        10'b1010011011: data <= 10'h000; 
        10'b1010011100: data <= 10'h000; 
        10'b1010011101: data <= 10'h000; 
        10'b1010011110: data <= 10'h000; 
        10'b1010011111: data <= 10'h000; 
        10'b1010100000: data <= 10'h000; 
        10'b1010100001: data <= 10'h000; 
        10'b1010100010: data <= 10'h000; 
        10'b1010100011: data <= 10'h000; 
        10'b1010100100: data <= 10'h001; 
        10'b1010100101: data <= 10'h001; 
        10'b1010100110: data <= 10'h001; 
        10'b1010100111: data <= 10'h000; 
        10'b1010101000: data <= 10'h3fe; 
        10'b1010101001: data <= 10'h3fe; 
        10'b1010101010: data <= 10'h3fc; 
        10'b1010101011: data <= 10'h3fd; 
        10'b1010101100: data <= 10'h3fd; 
        10'b1010101101: data <= 10'h3fd; 
        10'b1010101110: data <= 10'h3fd; 
        10'b1010101111: data <= 10'h3fd; 
        10'b1010110000: data <= 10'h3ff; 
        10'b1010110001: data <= 10'h000; 
        10'b1010110010: data <= 10'h001; 
        10'b1010110011: data <= 10'h001; 
        10'b1010110100: data <= 10'h001; 
        10'b1010110101: data <= 10'h000; 
        10'b1010110110: data <= 10'h000; 
        10'b1010110111: data <= 10'h001; 
        10'b1010111000: data <= 10'h000; 
        10'b1010111001: data <= 10'h000; 
        10'b1010111010: data <= 10'h001; 
        10'b1010111011: data <= 10'h000; 
        10'b1010111100: data <= 10'h001; 
        10'b1010111101: data <= 10'h000; 
        10'b1010111110: data <= 10'h000; 
        10'b1010111111: data <= 10'h001; 
        10'b1011000000: data <= 10'h001; 
        10'b1011000001: data <= 10'h001; 
        10'b1011000010: data <= 10'h000; 
        10'b1011000011: data <= 10'h3ff; 
        10'b1011000100: data <= 10'h000; 
        10'b1011000101: data <= 10'h000; 
        10'b1011000110: data <= 10'h3fe; 
        10'b1011000111: data <= 10'h3fe; 
        10'b1011001000: data <= 10'h3fe; 
        10'b1011001001: data <= 10'h3fe; 
        10'b1011001010: data <= 10'h3fe; 
        10'b1011001011: data <= 10'h3fe; 
        10'b1011001100: data <= 10'h3ff; 
        10'b1011001101: data <= 10'h000; 
        10'b1011001110: data <= 10'h000; 
        10'b1011001111: data <= 10'h001; 
        10'b1011010000: data <= 10'h000; 
        10'b1011010001: data <= 10'h001; 
        10'b1011010010: data <= 10'h000; 
        10'b1011010011: data <= 10'h001; 
        10'b1011010100: data <= 10'h000; 
        10'b1011010101: data <= 10'h000; 
        10'b1011010110: data <= 10'h000; 
        10'b1011010111: data <= 10'h000; 
        10'b1011011000: data <= 10'h000; 
        10'b1011011001: data <= 10'h001; 
        10'b1011011010: data <= 10'h001; 
        10'b1011011011: data <= 10'h000; 
        10'b1011011100: data <= 10'h001; 
        10'b1011011101: data <= 10'h001; 
        10'b1011011110: data <= 10'h001; 
        10'b1011011111: data <= 10'h001; 
        10'b1011100000: data <= 10'h001; 
        10'b1011100001: data <= 10'h001; 
        10'b1011100010: data <= 10'h000; 
        10'b1011100011: data <= 10'h001; 
        10'b1011100100: data <= 10'h001; 
        10'b1011100101: data <= 10'h000; 
        10'b1011100110: data <= 10'h000; 
        10'b1011100111: data <= 10'h000; 
        10'b1011101000: data <= 10'h001; 
        10'b1011101001: data <= 10'h001; 
        10'b1011101010: data <= 10'h001; 
        10'b1011101011: data <= 10'h000; 
        10'b1011101100: data <= 10'h001; 
        10'b1011101101: data <= 10'h001; 
        10'b1011101110: data <= 10'h001; 
        10'b1011101111: data <= 10'h000; 
        10'b1011110000: data <= 10'h000; 
        10'b1011110001: data <= 10'h001; 
        10'b1011110010: data <= 10'h001; 
        10'b1011110011: data <= 10'h001; 
        10'b1011110100: data <= 10'h001; 
        10'b1011110101: data <= 10'h001; 
        10'b1011110110: data <= 10'h000; 
        10'b1011110111: data <= 10'h001; 
        10'b1011111000: data <= 10'h001; 
        10'b1011111001: data <= 10'h001; 
        10'b1011111010: data <= 10'h001; 
        10'b1011111011: data <= 10'h001; 
        10'b1011111100: data <= 10'h001; 
        10'b1011111101: data <= 10'h001; 
        10'b1011111110: data <= 10'h001; 
        10'b1011111111: data <= 10'h001; 
        10'b1100000000: data <= 10'h000; 
        10'b1100000001: data <= 10'h000; 
        10'b1100000010: data <= 10'h001; 
        10'b1100000011: data <= 10'h001; 
        10'b1100000100: data <= 10'h001; 
        10'b1100000101: data <= 10'h000; 
        10'b1100000110: data <= 10'h001; 
        10'b1100000111: data <= 10'h000; 
        10'b1100001000: data <= 10'h000; 
        10'b1100001001: data <= 10'h000; 
        10'b1100001010: data <= 10'h001; 
        10'b1100001011: data <= 10'h001; 
        10'b1100001100: data <= 10'h001; 
        10'b1100001101: data <= 10'h001; 
        10'b1100001110: data <= 10'h001; 
        10'b1100001111: data <= 10'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 5) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 11'h002; 
        10'b0000000001: data <= 11'h001; 
        10'b0000000010: data <= 11'h001; 
        10'b0000000011: data <= 11'h000; 
        10'b0000000100: data <= 11'h002; 
        10'b0000000101: data <= 11'h002; 
        10'b0000000110: data <= 11'h002; 
        10'b0000000111: data <= 11'h000; 
        10'b0000001000: data <= 11'h002; 
        10'b0000001001: data <= 11'h000; 
        10'b0000001010: data <= 11'h002; 
        10'b0000001011: data <= 11'h001; 
        10'b0000001100: data <= 11'h002; 
        10'b0000001101: data <= 11'h002; 
        10'b0000001110: data <= 11'h002; 
        10'b0000001111: data <= 11'h001; 
        10'b0000010000: data <= 11'h001; 
        10'b0000010001: data <= 11'h000; 
        10'b0000010010: data <= 11'h002; 
        10'b0000010011: data <= 11'h002; 
        10'b0000010100: data <= 11'h001; 
        10'b0000010101: data <= 11'h002; 
        10'b0000010110: data <= 11'h001; 
        10'b0000010111: data <= 11'h002; 
        10'b0000011000: data <= 11'h001; 
        10'b0000011001: data <= 11'h002; 
        10'b0000011010: data <= 11'h001; 
        10'b0000011011: data <= 11'h002; 
        10'b0000011100: data <= 11'h000; 
        10'b0000011101: data <= 11'h002; 
        10'b0000011110: data <= 11'h001; 
        10'b0000011111: data <= 11'h001; 
        10'b0000100000: data <= 11'h001; 
        10'b0000100001: data <= 11'h001; 
        10'b0000100010: data <= 11'h001; 
        10'b0000100011: data <= 11'h002; 
        10'b0000100100: data <= 11'h002; 
        10'b0000100101: data <= 11'h001; 
        10'b0000100110: data <= 11'h001; 
        10'b0000100111: data <= 11'h001; 
        10'b0000101000: data <= 11'h002; 
        10'b0000101001: data <= 11'h002; 
        10'b0000101010: data <= 11'h003; 
        10'b0000101011: data <= 11'h001; 
        10'b0000101100: data <= 11'h001; 
        10'b0000101101: data <= 11'h002; 
        10'b0000101110: data <= 11'h001; 
        10'b0000101111: data <= 11'h001; 
        10'b0000110000: data <= 11'h002; 
        10'b0000110001: data <= 11'h002; 
        10'b0000110010: data <= 11'h001; 
        10'b0000110011: data <= 11'h002; 
        10'b0000110100: data <= 11'h002; 
        10'b0000110101: data <= 11'h001; 
        10'b0000110110: data <= 11'h002; 
        10'b0000110111: data <= 11'h002; 
        10'b0000111000: data <= 11'h002; 
        10'b0000111001: data <= 11'h002; 
        10'b0000111010: data <= 11'h002; 
        10'b0000111011: data <= 11'h000; 
        10'b0000111100: data <= 11'h000; 
        10'b0000111101: data <= 11'h002; 
        10'b0000111110: data <= 11'h001; 
        10'b0000111111: data <= 11'h001; 
        10'b0001000000: data <= 11'h001; 
        10'b0001000001: data <= 11'h001; 
        10'b0001000010: data <= 11'h000; 
        10'b0001000011: data <= 11'h001; 
        10'b0001000100: data <= 11'h000; 
        10'b0001000101: data <= 11'h001; 
        10'b0001000110: data <= 11'h001; 
        10'b0001000111: data <= 11'h002; 
        10'b0001001000: data <= 11'h002; 
        10'b0001001001: data <= 11'h000; 
        10'b0001001010: data <= 11'h001; 
        10'b0001001011: data <= 11'h001; 
        10'b0001001100: data <= 11'h002; 
        10'b0001001101: data <= 11'h001; 
        10'b0001001110: data <= 11'h002; 
        10'b0001001111: data <= 11'h002; 
        10'b0001010000: data <= 11'h002; 
        10'b0001010001: data <= 11'h000; 
        10'b0001010010: data <= 11'h002; 
        10'b0001010011: data <= 11'h002; 
        10'b0001010100: data <= 11'h001; 
        10'b0001010101: data <= 11'h001; 
        10'b0001010110: data <= 11'h001; 
        10'b0001010111: data <= 11'h001; 
        10'b0001011000: data <= 11'h002; 
        10'b0001011001: data <= 11'h001; 
        10'b0001011010: data <= 11'h000; 
        10'b0001011011: data <= 11'h002; 
        10'b0001011100: data <= 11'h000; 
        10'b0001011101: data <= 11'h000; 
        10'b0001011110: data <= 11'h000; 
        10'b0001011111: data <= 11'h7ff; 
        10'b0001100000: data <= 11'h000; 
        10'b0001100001: data <= 11'h000; 
        10'b0001100010: data <= 11'h001; 
        10'b0001100011: data <= 11'h002; 
        10'b0001100100: data <= 11'h7ff; 
        10'b0001100101: data <= 11'h000; 
        10'b0001100110: data <= 11'h000; 
        10'b0001100111: data <= 11'h7ff; 
        10'b0001101000: data <= 11'h000; 
        10'b0001101001: data <= 11'h001; 
        10'b0001101010: data <= 11'h001; 
        10'b0001101011: data <= 11'h001; 
        10'b0001101100: data <= 11'h000; 
        10'b0001101101: data <= 11'h002; 
        10'b0001101110: data <= 11'h001; 
        10'b0001101111: data <= 11'h002; 
        10'b0001110000: data <= 11'h002; 
        10'b0001110001: data <= 11'h001; 
        10'b0001110010: data <= 11'h002; 
        10'b0001110011: data <= 11'h002; 
        10'b0001110100: data <= 11'h000; 
        10'b0001110101: data <= 11'h000; 
        10'b0001110110: data <= 11'h002; 
        10'b0001110111: data <= 11'h001; 
        10'b0001111000: data <= 11'h000; 
        10'b0001111001: data <= 11'h7fe; 
        10'b0001111010: data <= 11'h000; 
        10'b0001111011: data <= 11'h001; 
        10'b0001111100: data <= 11'h001; 
        10'b0001111101: data <= 11'h002; 
        10'b0001111110: data <= 11'h002; 
        10'b0001111111: data <= 11'h005; 
        10'b0010000000: data <= 11'h001; 
        10'b0010000001: data <= 11'h7ff; 
        10'b0010000010: data <= 11'h7ff; 
        10'b0010000011: data <= 11'h001; 
        10'b0010000100: data <= 11'h003; 
        10'b0010000101: data <= 11'h003; 
        10'b0010000110: data <= 11'h003; 
        10'b0010000111: data <= 11'h004; 
        10'b0010001000: data <= 11'h002; 
        10'b0010001001: data <= 11'h001; 
        10'b0010001010: data <= 11'h001; 
        10'b0010001011: data <= 11'h001; 
        10'b0010001100: data <= 11'h000; 
        10'b0010001101: data <= 11'h002; 
        10'b0010001110: data <= 11'h000; 
        10'b0010001111: data <= 11'h001; 
        10'b0010010000: data <= 11'h000; 
        10'b0010010001: data <= 11'h001; 
        10'b0010010010: data <= 11'h000; 
        10'b0010010011: data <= 11'h7ff; 
        10'b0010010100: data <= 11'h7fc; 
        10'b0010010101: data <= 11'h7fc; 
        10'b0010010110: data <= 11'h7fe; 
        10'b0010010111: data <= 11'h000; 
        10'b0010011000: data <= 11'h002; 
        10'b0010011001: data <= 11'h002; 
        10'b0010011010: data <= 11'h003; 
        10'b0010011011: data <= 11'h003; 
        10'b0010011100: data <= 11'h002; 
        10'b0010011101: data <= 11'h7fe; 
        10'b0010011110: data <= 11'h000; 
        10'b0010011111: data <= 11'h001; 
        10'b0010100000: data <= 11'h002; 
        10'b0010100001: data <= 11'h004; 
        10'b0010100010: data <= 11'h007; 
        10'b0010100011: data <= 11'h004; 
        10'b0010100100: data <= 11'h003; 
        10'b0010100101: data <= 11'h7ff; 
        10'b0010100110: data <= 11'h001; 
        10'b0010100111: data <= 11'h001; 
        10'b0010101000: data <= 11'h000; 
        10'b0010101001: data <= 11'h001; 
        10'b0010101010: data <= 11'h000; 
        10'b0010101011: data <= 11'h001; 
        10'b0010101100: data <= 11'h000; 
        10'b0010101101: data <= 11'h7ff; 
        10'b0010101110: data <= 11'h7fe; 
        10'b0010101111: data <= 11'h7fe; 
        10'b0010110000: data <= 11'h7fa; 
        10'b0010110001: data <= 11'h7f9; 
        10'b0010110010: data <= 11'h7fc; 
        10'b0010110011: data <= 11'h7ff; 
        10'b0010110100: data <= 11'h7ff; 
        10'b0010110101: data <= 11'h7fe; 
        10'b0010110110: data <= 11'h7ff; 
        10'b0010110111: data <= 11'h7fb; 
        10'b0010111000: data <= 11'h7fb; 
        10'b0010111001: data <= 11'h7fb; 
        10'b0010111010: data <= 11'h7fe; 
        10'b0010111011: data <= 11'h7fe; 
        10'b0010111100: data <= 11'h002; 
        10'b0010111101: data <= 11'h004; 
        10'b0010111110: data <= 11'h004; 
        10'b0010111111: data <= 11'h003; 
        10'b0011000000: data <= 11'h001; 
        10'b0011000001: data <= 11'h7ff; 
        10'b0011000010: data <= 11'h000; 
        10'b0011000011: data <= 11'h001; 
        10'b0011000100: data <= 11'h001; 
        10'b0011000101: data <= 11'h001; 
        10'b0011000110: data <= 11'h001; 
        10'b0011000111: data <= 11'h000; 
        10'b0011001000: data <= 11'h002; 
        10'b0011001001: data <= 11'h000; 
        10'b0011001010: data <= 11'h7fe; 
        10'b0011001011: data <= 11'h7fb; 
        10'b0011001100: data <= 11'h7f8; 
        10'b0011001101: data <= 11'h7f6; 
        10'b0011001110: data <= 11'h7fa; 
        10'b0011001111: data <= 11'h7fd; 
        10'b0011010000: data <= 11'h7fd; 
        10'b0011010001: data <= 11'h7fc; 
        10'b0011010010: data <= 11'h7fb; 
        10'b0011010011: data <= 11'h7f9; 
        10'b0011010100: data <= 11'h7fa; 
        10'b0011010101: data <= 11'h7fa; 
        10'b0011010110: data <= 11'h7fb; 
        10'b0011010111: data <= 11'h000; 
        10'b0011011000: data <= 11'h001; 
        10'b0011011001: data <= 11'h001; 
        10'b0011011010: data <= 11'h001; 
        10'b0011011011: data <= 11'h7fe; 
        10'b0011011100: data <= 11'h7fd; 
        10'b0011011101: data <= 11'h7ff; 
        10'b0011011110: data <= 11'h001; 
        10'b0011011111: data <= 11'h001; 
        10'b0011100000: data <= 11'h001; 
        10'b0011100001: data <= 11'h001; 
        10'b0011100010: data <= 11'h001; 
        10'b0011100011: data <= 11'h002; 
        10'b0011100100: data <= 11'h001; 
        10'b0011100101: data <= 11'h000; 
        10'b0011100110: data <= 11'h7fd; 
        10'b0011100111: data <= 11'h7fc; 
        10'b0011101000: data <= 11'h7f7; 
        10'b0011101001: data <= 11'h7f6; 
        10'b0011101010: data <= 11'h7f7; 
        10'b0011101011: data <= 11'h7fb; 
        10'b0011101100: data <= 11'h7fe; 
        10'b0011101101: data <= 11'h7fd; 
        10'b0011101110: data <= 11'h7fe; 
        10'b0011101111: data <= 11'h001; 
        10'b0011110000: data <= 11'h7fc; 
        10'b0011110001: data <= 11'h7ff; 
        10'b0011110010: data <= 11'h000; 
        10'b0011110011: data <= 11'h001; 
        10'b0011110100: data <= 11'h7fd; 
        10'b0011110101: data <= 11'h7fd; 
        10'b0011110110: data <= 11'h7fb; 
        10'b0011110111: data <= 11'h7fa; 
        10'b0011111000: data <= 11'h7fb; 
        10'b0011111001: data <= 11'h7ff; 
        10'b0011111010: data <= 11'h002; 
        10'b0011111011: data <= 11'h002; 
        10'b0011111100: data <= 11'h002; 
        10'b0011111101: data <= 11'h001; 
        10'b0011111110: data <= 11'h001; 
        10'b0011111111: data <= 11'h001; 
        10'b0100000000: data <= 11'h000; 
        10'b0100000001: data <= 11'h000; 
        10'b0100000010: data <= 11'h7fc; 
        10'b0100000011: data <= 11'h7fd; 
        10'b0100000100: data <= 11'h7fa; 
        10'b0100000101: data <= 11'h7f7; 
        10'b0100000110: data <= 11'h7f8; 
        10'b0100000111: data <= 11'h7fd; 
        10'b0100001000: data <= 11'h7fe; 
        10'b0100001001: data <= 11'h002; 
        10'b0100001010: data <= 11'h006; 
        10'b0100001011: data <= 11'h009; 
        10'b0100001100: data <= 11'h003; 
        10'b0100001101: data <= 11'h000; 
        10'b0100001110: data <= 11'h7ff; 
        10'b0100001111: data <= 11'h7fa; 
        10'b0100010000: data <= 11'h7f9; 
        10'b0100010001: data <= 11'h7f9; 
        10'b0100010010: data <= 11'h7f7; 
        10'b0100010011: data <= 11'h7f8; 
        10'b0100010100: data <= 11'h7fc; 
        10'b0100010101: data <= 11'h000; 
        10'b0100010110: data <= 11'h002; 
        10'b0100010111: data <= 11'h001; 
        10'b0100011000: data <= 11'h002; 
        10'b0100011001: data <= 11'h002; 
        10'b0100011010: data <= 11'h002; 
        10'b0100011011: data <= 11'h000; 
        10'b0100011100: data <= 11'h002; 
        10'b0100011101: data <= 11'h7fe; 
        10'b0100011110: data <= 11'h7fd; 
        10'b0100011111: data <= 11'h7fe; 
        10'b0100100000: data <= 11'h7fb; 
        10'b0100100001: data <= 11'h7fb; 
        10'b0100100010: data <= 11'h7fd; 
        10'b0100100011: data <= 11'h7fe; 
        10'b0100100100: data <= 11'h7fe; 
        10'b0100100101: data <= 11'h005; 
        10'b0100100110: data <= 11'h00f; 
        10'b0100100111: data <= 11'h010; 
        10'b0100101000: data <= 11'h008; 
        10'b0100101001: data <= 11'h000; 
        10'b0100101010: data <= 11'h7fb; 
        10'b0100101011: data <= 11'h7fa; 
        10'b0100101100: data <= 11'h7f9; 
        10'b0100101101: data <= 11'h7fa; 
        10'b0100101110: data <= 11'h7fa; 
        10'b0100101111: data <= 11'h7fc; 
        10'b0100110000: data <= 11'h7ff; 
        10'b0100110001: data <= 11'h000; 
        10'b0100110010: data <= 11'h002; 
        10'b0100110011: data <= 11'h001; 
        10'b0100110100: data <= 11'h000; 
        10'b0100110101: data <= 11'h000; 
        10'b0100110110: data <= 11'h002; 
        10'b0100110111: data <= 11'h002; 
        10'b0100111000: data <= 11'h000; 
        10'b0100111001: data <= 11'h7ff; 
        10'b0100111010: data <= 11'h000; 
        10'b0100111011: data <= 11'h7fd; 
        10'b0100111100: data <= 11'h7fe; 
        10'b0100111101: data <= 11'h7fd; 
        10'b0100111110: data <= 11'h7fc; 
        10'b0100111111: data <= 11'h7fa; 
        10'b0101000000: data <= 11'h7ff; 
        10'b0101000001: data <= 11'h008; 
        10'b0101000010: data <= 11'h013; 
        10'b0101000011: data <= 11'h014; 
        10'b0101000100: data <= 11'h007; 
        10'b0101000101: data <= 11'h7fe; 
        10'b0101000110: data <= 11'h7ff; 
        10'b0101000111: data <= 11'h7fc; 
        10'b0101001000: data <= 11'h7fc; 
        10'b0101001001: data <= 11'h7fc; 
        10'b0101001010: data <= 11'h7fc; 
        10'b0101001011: data <= 11'h7fe; 
        10'b0101001100: data <= 11'h7ff; 
        10'b0101001101: data <= 11'h002; 
        10'b0101001110: data <= 11'h002; 
        10'b0101001111: data <= 11'h002; 
        10'b0101010000: data <= 11'h000; 
        10'b0101010001: data <= 11'h002; 
        10'b0101010010: data <= 11'h001; 
        10'b0101010011: data <= 11'h001; 
        10'b0101010100: data <= 11'h002; 
        10'b0101010101: data <= 11'h000; 
        10'b0101010110: data <= 11'h7ff; 
        10'b0101010111: data <= 11'h7ff; 
        10'b0101011000: data <= 11'h7fd; 
        10'b0101011001: data <= 11'h7fc; 
        10'b0101011010: data <= 11'h7f8; 
        10'b0101011011: data <= 11'h7f5; 
        10'b0101011100: data <= 11'h000; 
        10'b0101011101: data <= 11'h008; 
        10'b0101011110: data <= 11'h016; 
        10'b0101011111: data <= 11'h00f; 
        10'b0101100000: data <= 11'h003; 
        10'b0101100001: data <= 11'h002; 
        10'b0101100010: data <= 11'h7ff; 
        10'b0101100011: data <= 11'h7fc; 
        10'b0101100100: data <= 11'h7fd; 
        10'b0101100101: data <= 11'h7ff; 
        10'b0101100110: data <= 11'h7ff; 
        10'b0101100111: data <= 11'h7ff; 
        10'b0101101000: data <= 11'h000; 
        10'b0101101001: data <= 11'h002; 
        10'b0101101010: data <= 11'h000; 
        10'b0101101011: data <= 11'h002; 
        10'b0101101100: data <= 11'h000; 
        10'b0101101101: data <= 11'h001; 
        10'b0101101110: data <= 11'h001; 
        10'b0101101111: data <= 11'h001; 
        10'b0101110000: data <= 11'h002; 
        10'b0101110001: data <= 11'h000; 
        10'b0101110010: data <= 11'h000; 
        10'b0101110011: data <= 11'h7ff; 
        10'b0101110100: data <= 11'h7ff; 
        10'b0101110101: data <= 11'h7fa; 
        10'b0101110110: data <= 11'h7f3; 
        10'b0101110111: data <= 11'h7f3; 
        10'b0101111000: data <= 11'h000; 
        10'b0101111001: data <= 11'h007; 
        10'b0101111010: data <= 11'h012; 
        10'b0101111011: data <= 11'h00a; 
        10'b0101111100: data <= 11'h003; 
        10'b0101111101: data <= 11'h001; 
        10'b0101111110: data <= 11'h7fc; 
        10'b0101111111: data <= 11'h7fa; 
        10'b0110000000: data <= 11'h7fe; 
        10'b0110000001: data <= 11'h7ff; 
        10'b0110000010: data <= 11'h7ff; 
        10'b0110000011: data <= 11'h000; 
        10'b0110000100: data <= 11'h001; 
        10'b0110000101: data <= 11'h002; 
        10'b0110000110: data <= 11'h002; 
        10'b0110000111: data <= 11'h001; 
        10'b0110001000: data <= 11'h001; 
        10'b0110001001: data <= 11'h002; 
        10'b0110001010: data <= 11'h001; 
        10'b0110001011: data <= 11'h002; 
        10'b0110001100: data <= 11'h002; 
        10'b0110001101: data <= 11'h000; 
        10'b0110001110: data <= 11'h000; 
        10'b0110001111: data <= 11'h7ff; 
        10'b0110010000: data <= 11'h7fc; 
        10'b0110010001: data <= 11'h7f9; 
        10'b0110010010: data <= 11'h7f3; 
        10'b0110010011: data <= 11'h7f6; 
        10'b0110010100: data <= 11'h000; 
        10'b0110010101: data <= 11'h007; 
        10'b0110010110: data <= 11'h00f; 
        10'b0110010111: data <= 11'h00a; 
        10'b0110011000: data <= 11'h003; 
        10'b0110011001: data <= 11'h7fb; 
        10'b0110011010: data <= 11'h7f9; 
        10'b0110011011: data <= 11'h7fa; 
        10'b0110011100: data <= 11'h7fd; 
        10'b0110011101: data <= 11'h7ff; 
        10'b0110011110: data <= 11'h7ff; 
        10'b0110011111: data <= 11'h7ff; 
        10'b0110100000: data <= 11'h002; 
        10'b0110100001: data <= 11'h000; 
        10'b0110100010: data <= 11'h000; 
        10'b0110100011: data <= 11'h001; 
        10'b0110100100: data <= 11'h002; 
        10'b0110100101: data <= 11'h000; 
        10'b0110100110: data <= 11'h002; 
        10'b0110100111: data <= 11'h001; 
        10'b0110101000: data <= 11'h001; 
        10'b0110101001: data <= 11'h001; 
        10'b0110101010: data <= 11'h7ff; 
        10'b0110101011: data <= 11'h7fe; 
        10'b0110101100: data <= 11'h7fd; 
        10'b0110101101: data <= 11'h7f8; 
        10'b0110101110: data <= 11'h7f8; 
        10'b0110101111: data <= 11'h7fe; 
        10'b0110110000: data <= 11'h003; 
        10'b0110110001: data <= 11'h00a; 
        10'b0110110010: data <= 11'h010; 
        10'b0110110011: data <= 11'h006; 
        10'b0110110100: data <= 11'h001; 
        10'b0110110101: data <= 11'h7f6; 
        10'b0110110110: data <= 11'h7f7; 
        10'b0110110111: data <= 11'h7fa; 
        10'b0110111000: data <= 11'h7fd; 
        10'b0110111001: data <= 11'h7fe; 
        10'b0110111010: data <= 11'h7ff; 
        10'b0110111011: data <= 11'h000; 
        10'b0110111100: data <= 11'h001; 
        10'b0110111101: data <= 11'h001; 
        10'b0110111110: data <= 11'h002; 
        10'b0110111111: data <= 11'h000; 
        10'b0111000000: data <= 11'h002; 
        10'b0111000001: data <= 11'h001; 
        10'b0111000010: data <= 11'h002; 
        10'b0111000011: data <= 11'h001; 
        10'b0111000100: data <= 11'h001; 
        10'b0111000101: data <= 11'h7ff; 
        10'b0111000110: data <= 11'h7fe; 
        10'b0111000111: data <= 11'h7fe; 
        10'b0111001000: data <= 11'h7fa; 
        10'b0111001001: data <= 11'h7fc; 
        10'b0111001010: data <= 11'h7fd; 
        10'b0111001011: data <= 11'h7fe; 
        10'b0111001100: data <= 11'h000; 
        10'b0111001101: data <= 11'h00d; 
        10'b0111001110: data <= 11'h00f; 
        10'b0111001111: data <= 11'h001; 
        10'b0111010000: data <= 11'h7fb; 
        10'b0111010001: data <= 11'h7f5; 
        10'b0111010010: data <= 11'h7f7; 
        10'b0111010011: data <= 11'h7fa; 
        10'b0111010100: data <= 11'h7fb; 
        10'b0111010101: data <= 11'h7fe; 
        10'b0111010110: data <= 11'h7fe; 
        10'b0111010111: data <= 11'h000; 
        10'b0111011000: data <= 11'h7ff; 
        10'b0111011001: data <= 11'h000; 
        10'b0111011010: data <= 11'h001; 
        10'b0111011011: data <= 11'h001; 
        10'b0111011100: data <= 11'h001; 
        10'b0111011101: data <= 11'h002; 
        10'b0111011110: data <= 11'h001; 
        10'b0111011111: data <= 11'h002; 
        10'b0111100000: data <= 11'h002; 
        10'b0111100001: data <= 11'h7ff; 
        10'b0111100010: data <= 11'h7fb; 
        10'b0111100011: data <= 11'h7fb; 
        10'b0111100100: data <= 11'h7fc; 
        10'b0111100101: data <= 11'h7fe; 
        10'b0111100110: data <= 11'h002; 
        10'b0111100111: data <= 11'h000; 
        10'b0111101000: data <= 11'h004; 
        10'b0111101001: data <= 11'h00f; 
        10'b0111101010: data <= 11'h00d; 
        10'b0111101011: data <= 11'h7fd; 
        10'b0111101100: data <= 11'h7f7; 
        10'b0111101101: data <= 11'h7f5; 
        10'b0111101110: data <= 11'h7f7; 
        10'b0111101111: data <= 11'h7fa; 
        10'b0111110000: data <= 11'h7fe; 
        10'b0111110001: data <= 11'h7ff; 
        10'b0111110010: data <= 11'h7ff; 
        10'b0111110011: data <= 11'h7ff; 
        10'b0111110100: data <= 11'h7fe; 
        10'b0111110101: data <= 11'h001; 
        10'b0111110110: data <= 11'h001; 
        10'b0111110111: data <= 11'h002; 
        10'b0111111000: data <= 11'h001; 
        10'b0111111001: data <= 11'h001; 
        10'b0111111010: data <= 11'h001; 
        10'b0111111011: data <= 11'h002; 
        10'b0111111100: data <= 11'h001; 
        10'b0111111101: data <= 11'h7fe; 
        10'b0111111110: data <= 11'h7fb; 
        10'b0111111111: data <= 11'h7fb; 
        10'b1000000000: data <= 11'h7fe; 
        10'b1000000001: data <= 11'h002; 
        10'b1000000010: data <= 11'h002; 
        10'b1000000011: data <= 11'h003; 
        10'b1000000100: data <= 11'h007; 
        10'b1000000101: data <= 11'h00b; 
        10'b1000000110: data <= 11'h008; 
        10'b1000000111: data <= 11'h7fb; 
        10'b1000001000: data <= 11'h7f8; 
        10'b1000001001: data <= 11'h7f9; 
        10'b1000001010: data <= 11'h7fa; 
        10'b1000001011: data <= 11'h7fc; 
        10'b1000001100: data <= 11'h7fe; 
        10'b1000001101: data <= 11'h7fd; 
        10'b1000001110: data <= 11'h7ff; 
        10'b1000001111: data <= 11'h7fe; 
        10'b1000010000: data <= 11'h7ff; 
        10'b1000010001: data <= 11'h001; 
        10'b1000010010: data <= 11'h002; 
        10'b1000010011: data <= 11'h002; 
        10'b1000010100: data <= 11'h002; 
        10'b1000010101: data <= 11'h002; 
        10'b1000010110: data <= 11'h002; 
        10'b1000010111: data <= 11'h002; 
        10'b1000011000: data <= 11'h000; 
        10'b1000011001: data <= 11'h7fd; 
        10'b1000011010: data <= 11'h7fa; 
        10'b1000011011: data <= 11'h7fc; 
        10'b1000011100: data <= 11'h7fe; 
        10'b1000011101: data <= 11'h001; 
        10'b1000011110: data <= 11'h001; 
        10'b1000011111: data <= 11'h000; 
        10'b1000100000: data <= 11'h001; 
        10'b1000100001: data <= 11'h005; 
        10'b1000100010: data <= 11'h001; 
        10'b1000100011: data <= 11'h7fc; 
        10'b1000100100: data <= 11'h7fd; 
        10'b1000100101: data <= 11'h7fd; 
        10'b1000100110: data <= 11'h7fc; 
        10'b1000100111: data <= 11'h7fd; 
        10'b1000101000: data <= 11'h7fc; 
        10'b1000101001: data <= 11'h7fc; 
        10'b1000101010: data <= 11'h7fe; 
        10'b1000101011: data <= 11'h7fe; 
        10'b1000101100: data <= 11'h000; 
        10'b1000101101: data <= 11'h001; 
        10'b1000101110: data <= 11'h001; 
        10'b1000101111: data <= 11'h000; 
        10'b1000110000: data <= 11'h000; 
        10'b1000110001: data <= 11'h002; 
        10'b1000110010: data <= 11'h001; 
        10'b1000110011: data <= 11'h001; 
        10'b1000110100: data <= 11'h7ff; 
        10'b1000110101: data <= 11'h7fe; 
        10'b1000110110: data <= 11'h000; 
        10'b1000110111: data <= 11'h7ff; 
        10'b1000111000: data <= 11'h000; 
        10'b1000111001: data <= 11'h001; 
        10'b1000111010: data <= 11'h7fe; 
        10'b1000111011: data <= 11'h7ff; 
        10'b1000111100: data <= 11'h7fd; 
        10'b1000111101: data <= 11'h7ff; 
        10'b1000111110: data <= 11'h7ff; 
        10'b1000111111: data <= 11'h000; 
        10'b1001000000: data <= 11'h002; 
        10'b1001000001: data <= 11'h001; 
        10'b1001000010: data <= 11'h7ff; 
        10'b1001000011: data <= 11'h7fd; 
        10'b1001000100: data <= 11'h7fc; 
        10'b1001000101: data <= 11'h7fc; 
        10'b1001000110: data <= 11'h7fd; 
        10'b1001000111: data <= 11'h7ff; 
        10'b1001001000: data <= 11'h000; 
        10'b1001001001: data <= 11'h002; 
        10'b1001001010: data <= 11'h001; 
        10'b1001001011: data <= 11'h002; 
        10'b1001001100: data <= 11'h002; 
        10'b1001001101: data <= 11'h001; 
        10'b1001001110: data <= 11'h001; 
        10'b1001001111: data <= 11'h002; 
        10'b1001010000: data <= 11'h001; 
        10'b1001010001: data <= 11'h004; 
        10'b1001010010: data <= 11'h003; 
        10'b1001010011: data <= 11'h001; 
        10'b1001010100: data <= 11'h000; 
        10'b1001010101: data <= 11'h7ff; 
        10'b1001010110: data <= 11'h000; 
        10'b1001010111: data <= 11'h7fe; 
        10'b1001011000: data <= 11'h7fb; 
        10'b1001011001: data <= 11'h7fb; 
        10'b1001011010: data <= 11'h000; 
        10'b1001011011: data <= 11'h002; 
        10'b1001011100: data <= 11'h003; 
        10'b1001011101: data <= 11'h003; 
        10'b1001011110: data <= 11'h002; 
        10'b1001011111: data <= 11'h7fd; 
        10'b1001100000: data <= 11'h7fd; 
        10'b1001100001: data <= 11'h7fc; 
        10'b1001100010: data <= 11'h7fd; 
        10'b1001100011: data <= 11'h7fe; 
        10'b1001100100: data <= 11'h000; 
        10'b1001100101: data <= 11'h001; 
        10'b1001100110: data <= 11'h000; 
        10'b1001100111: data <= 11'h000; 
        10'b1001101000: data <= 11'h001; 
        10'b1001101001: data <= 11'h001; 
        10'b1001101010: data <= 11'h002; 
        10'b1001101011: data <= 11'h000; 
        10'b1001101100: data <= 11'h003; 
        10'b1001101101: data <= 11'h007; 
        10'b1001101110: data <= 11'h007; 
        10'b1001101111: data <= 11'h004; 
        10'b1001110000: data <= 11'h001; 
        10'b1001110001: data <= 11'h000; 
        10'b1001110010: data <= 11'h7fe; 
        10'b1001110011: data <= 11'h7f9; 
        10'b1001110100: data <= 11'h7f5; 
        10'b1001110101: data <= 11'h7f7; 
        10'b1001110110: data <= 11'h000; 
        10'b1001110111: data <= 11'h002; 
        10'b1001111000: data <= 11'h006; 
        10'b1001111001: data <= 11'h00b; 
        10'b1001111010: data <= 11'h005; 
        10'b1001111011: data <= 11'h001; 
        10'b1001111100: data <= 11'h7fe; 
        10'b1001111101: data <= 11'h7fe; 
        10'b1001111110: data <= 11'h000; 
        10'b1001111111: data <= 11'h000; 
        10'b1010000000: data <= 11'h000; 
        10'b1010000001: data <= 11'h001; 
        10'b1010000010: data <= 11'h002; 
        10'b1010000011: data <= 11'h001; 
        10'b1010000100: data <= 11'h002; 
        10'b1010000101: data <= 11'h001; 
        10'b1010000110: data <= 11'h002; 
        10'b1010000111: data <= 11'h001; 
        10'b1010001000: data <= 11'h003; 
        10'b1010001001: data <= 11'h006; 
        10'b1010001010: data <= 11'h006; 
        10'b1010001011: data <= 11'h003; 
        10'b1010001100: data <= 11'h001; 
        10'b1010001101: data <= 11'h7fe; 
        10'b1010001110: data <= 11'h7ff; 
        10'b1010001111: data <= 11'h7fc; 
        10'b1010010000: data <= 11'h7fd; 
        10'b1010010001: data <= 11'h7fe; 
        10'b1010010010: data <= 11'h7fd; 
        10'b1010010011: data <= 11'h001; 
        10'b1010010100: data <= 11'h008; 
        10'b1010010101: data <= 11'h009; 
        10'b1010010110: data <= 11'h004; 
        10'b1010010111: data <= 11'h7ff; 
        10'b1010011000: data <= 11'h7fe; 
        10'b1010011001: data <= 11'h7fd; 
        10'b1010011010: data <= 11'h7ff; 
        10'b1010011011: data <= 11'h7ff; 
        10'b1010011100: data <= 11'h001; 
        10'b1010011101: data <= 11'h000; 
        10'b1010011110: data <= 11'h001; 
        10'b1010011111: data <= 11'h000; 
        10'b1010100000: data <= 11'h001; 
        10'b1010100001: data <= 11'h000; 
        10'b1010100010: data <= 11'h001; 
        10'b1010100011: data <= 11'h000; 
        10'b1010100100: data <= 11'h001; 
        10'b1010100101: data <= 11'h003; 
        10'b1010100110: data <= 11'h003; 
        10'b1010100111: data <= 11'h7ff; 
        10'b1010101000: data <= 11'h7fc; 
        10'b1010101001: data <= 11'h7fc; 
        10'b1010101010: data <= 11'h7f9; 
        10'b1010101011: data <= 11'h7f9; 
        10'b1010101100: data <= 11'h7fa; 
        10'b1010101101: data <= 11'h7fb; 
        10'b1010101110: data <= 11'h7fb; 
        10'b1010101111: data <= 11'h7fb; 
        10'b1010110000: data <= 11'h7fe; 
        10'b1010110001: data <= 11'h001; 
        10'b1010110010: data <= 11'h001; 
        10'b1010110011: data <= 11'h002; 
        10'b1010110100: data <= 11'h001; 
        10'b1010110101: data <= 11'h000; 
        10'b1010110110: data <= 11'h001; 
        10'b1010110111: data <= 11'h002; 
        10'b1010111000: data <= 11'h001; 
        10'b1010111001: data <= 11'h001; 
        10'b1010111010: data <= 11'h002; 
        10'b1010111011: data <= 11'h001; 
        10'b1010111100: data <= 11'h002; 
        10'b1010111101: data <= 11'h001; 
        10'b1010111110: data <= 11'h001; 
        10'b1010111111: data <= 11'h001; 
        10'b1011000000: data <= 11'h002; 
        10'b1011000001: data <= 11'h002; 
        10'b1011000010: data <= 11'h000; 
        10'b1011000011: data <= 11'h7ff; 
        10'b1011000100: data <= 11'h000; 
        10'b1011000101: data <= 11'h7ff; 
        10'b1011000110: data <= 11'h7fc; 
        10'b1011000111: data <= 11'h7fb; 
        10'b1011001000: data <= 11'h7fc; 
        10'b1011001001: data <= 11'h7fb; 
        10'b1011001010: data <= 11'h7fd; 
        10'b1011001011: data <= 11'h7fc; 
        10'b1011001100: data <= 11'h7fe; 
        10'b1011001101: data <= 11'h000; 
        10'b1011001110: data <= 11'h001; 
        10'b1011001111: data <= 11'h002; 
        10'b1011010000: data <= 11'h000; 
        10'b1011010001: data <= 11'h001; 
        10'b1011010010: data <= 11'h001; 
        10'b1011010011: data <= 11'h002; 
        10'b1011010100: data <= 11'h001; 
        10'b1011010101: data <= 11'h001; 
        10'b1011010110: data <= 11'h001; 
        10'b1011010111: data <= 11'h001; 
        10'b1011011000: data <= 11'h001; 
        10'b1011011001: data <= 11'h002; 
        10'b1011011010: data <= 11'h001; 
        10'b1011011011: data <= 11'h000; 
        10'b1011011100: data <= 11'h002; 
        10'b1011011101: data <= 11'h002; 
        10'b1011011110: data <= 11'h001; 
        10'b1011011111: data <= 11'h001; 
        10'b1011100000: data <= 11'h002; 
        10'b1011100001: data <= 11'h002; 
        10'b1011100010: data <= 11'h000; 
        10'b1011100011: data <= 11'h001; 
        10'b1011100100: data <= 11'h001; 
        10'b1011100101: data <= 11'h001; 
        10'b1011100110: data <= 11'h000; 
        10'b1011100111: data <= 11'h001; 
        10'b1011101000: data <= 11'h001; 
        10'b1011101001: data <= 11'h002; 
        10'b1011101010: data <= 11'h002; 
        10'b1011101011: data <= 11'h000; 
        10'b1011101100: data <= 11'h001; 
        10'b1011101101: data <= 11'h001; 
        10'b1011101110: data <= 11'h001; 
        10'b1011101111: data <= 11'h001; 
        10'b1011110000: data <= 11'h001; 
        10'b1011110001: data <= 11'h002; 
        10'b1011110010: data <= 11'h002; 
        10'b1011110011: data <= 11'h002; 
        10'b1011110100: data <= 11'h002; 
        10'b1011110101: data <= 11'h002; 
        10'b1011110110: data <= 11'h000; 
        10'b1011110111: data <= 11'h001; 
        10'b1011111000: data <= 11'h002; 
        10'b1011111001: data <= 11'h002; 
        10'b1011111010: data <= 11'h002; 
        10'b1011111011: data <= 11'h002; 
        10'b1011111100: data <= 11'h002; 
        10'b1011111101: data <= 11'h001; 
        10'b1011111110: data <= 11'h002; 
        10'b1011111111: data <= 11'h002; 
        10'b1100000000: data <= 11'h000; 
        10'b1100000001: data <= 11'h000; 
        10'b1100000010: data <= 11'h002; 
        10'b1100000011: data <= 11'h002; 
        10'b1100000100: data <= 11'h001; 
        10'b1100000101: data <= 11'h000; 
        10'b1100000110: data <= 11'h001; 
        10'b1100000111: data <= 11'h000; 
        10'b1100001000: data <= 11'h000; 
        10'b1100001001: data <= 11'h001; 
        10'b1100001010: data <= 11'h001; 
        10'b1100001011: data <= 11'h002; 
        10'b1100001100: data <= 11'h002; 
        10'b1100001101: data <= 11'h002; 
        10'b1100001110: data <= 11'h002; 
        10'b1100001111: data <= 11'h001; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 6) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 12'h004; 
        10'b0000000001: data <= 12'h002; 
        10'b0000000010: data <= 12'h002; 
        10'b0000000011: data <= 12'h001; 
        10'b0000000100: data <= 12'h003; 
        10'b0000000101: data <= 12'h003; 
        10'b0000000110: data <= 12'h004; 
        10'b0000000111: data <= 12'h001; 
        10'b0000001000: data <= 12'h003; 
        10'b0000001001: data <= 12'h001; 
        10'b0000001010: data <= 12'h003; 
        10'b0000001011: data <= 12'h002; 
        10'b0000001100: data <= 12'h003; 
        10'b0000001101: data <= 12'h005; 
        10'b0000001110: data <= 12'h004; 
        10'b0000001111: data <= 12'h003; 
        10'b0000010000: data <= 12'h003; 
        10'b0000010001: data <= 12'h001; 
        10'b0000010010: data <= 12'h005; 
        10'b0000010011: data <= 12'h005; 
        10'b0000010100: data <= 12'h003; 
        10'b0000010101: data <= 12'h003; 
        10'b0000010110: data <= 12'h003; 
        10'b0000010111: data <= 12'h004; 
        10'b0000011000: data <= 12'h002; 
        10'b0000011001: data <= 12'h004; 
        10'b0000011010: data <= 12'h003; 
        10'b0000011011: data <= 12'h004; 
        10'b0000011100: data <= 12'h000; 
        10'b0000011101: data <= 12'h004; 
        10'b0000011110: data <= 12'h001; 
        10'b0000011111: data <= 12'h003; 
        10'b0000100000: data <= 12'h003; 
        10'b0000100001: data <= 12'h001; 
        10'b0000100010: data <= 12'h001; 
        10'b0000100011: data <= 12'h004; 
        10'b0000100100: data <= 12'h004; 
        10'b0000100101: data <= 12'h003; 
        10'b0000100110: data <= 12'h003; 
        10'b0000100111: data <= 12'h002; 
        10'b0000101000: data <= 12'h003; 
        10'b0000101001: data <= 12'h004; 
        10'b0000101010: data <= 12'h005; 
        10'b0000101011: data <= 12'h003; 
        10'b0000101100: data <= 12'h002; 
        10'b0000101101: data <= 12'h004; 
        10'b0000101110: data <= 12'h003; 
        10'b0000101111: data <= 12'h002; 
        10'b0000110000: data <= 12'h004; 
        10'b0000110001: data <= 12'h004; 
        10'b0000110010: data <= 12'h002; 
        10'b0000110011: data <= 12'h005; 
        10'b0000110100: data <= 12'h005; 
        10'b0000110101: data <= 12'h003; 
        10'b0000110110: data <= 12'h004; 
        10'b0000110111: data <= 12'h003; 
        10'b0000111000: data <= 12'h004; 
        10'b0000111001: data <= 12'h003; 
        10'b0000111010: data <= 12'h005; 
        10'b0000111011: data <= 12'h001; 
        10'b0000111100: data <= 12'h001; 
        10'b0000111101: data <= 12'h003; 
        10'b0000111110: data <= 12'h002; 
        10'b0000111111: data <= 12'h002; 
        10'b0001000000: data <= 12'h002; 
        10'b0001000001: data <= 12'h003; 
        10'b0001000010: data <= 12'h000; 
        10'b0001000011: data <= 12'h001; 
        10'b0001000100: data <= 12'h000; 
        10'b0001000101: data <= 12'h001; 
        10'b0001000110: data <= 12'h002; 
        10'b0001000111: data <= 12'h004; 
        10'b0001001000: data <= 12'h003; 
        10'b0001001001: data <= 12'h000; 
        10'b0001001010: data <= 12'h003; 
        10'b0001001011: data <= 12'h002; 
        10'b0001001100: data <= 12'h004; 
        10'b0001001101: data <= 12'h002; 
        10'b0001001110: data <= 12'h004; 
        10'b0001001111: data <= 12'h003; 
        10'b0001010000: data <= 12'h003; 
        10'b0001010001: data <= 12'h001; 
        10'b0001010010: data <= 12'h004; 
        10'b0001010011: data <= 12'h004; 
        10'b0001010100: data <= 12'h001; 
        10'b0001010101: data <= 12'h002; 
        10'b0001010110: data <= 12'h003; 
        10'b0001010111: data <= 12'h002; 
        10'b0001011000: data <= 12'h005; 
        10'b0001011001: data <= 12'h002; 
        10'b0001011010: data <= 12'h001; 
        10'b0001011011: data <= 12'h004; 
        10'b0001011100: data <= 12'h000; 
        10'b0001011101: data <= 12'hfff; 
        10'b0001011110: data <= 12'hfff; 
        10'b0001011111: data <= 12'hffd; 
        10'b0001100000: data <= 12'hfff; 
        10'b0001100001: data <= 12'h000; 
        10'b0001100010: data <= 12'h002; 
        10'b0001100011: data <= 12'h004; 
        10'b0001100100: data <= 12'hffe; 
        10'b0001100101: data <= 12'hfff; 
        10'b0001100110: data <= 12'h000; 
        10'b0001100111: data <= 12'hffd; 
        10'b0001101000: data <= 12'h000; 
        10'b0001101001: data <= 12'h001; 
        10'b0001101010: data <= 12'h003; 
        10'b0001101011: data <= 12'h003; 
        10'b0001101100: data <= 12'hfff; 
        10'b0001101101: data <= 12'h004; 
        10'b0001101110: data <= 12'h002; 
        10'b0001101111: data <= 12'h004; 
        10'b0001110000: data <= 12'h003; 
        10'b0001110001: data <= 12'h002; 
        10'b0001110010: data <= 12'h005; 
        10'b0001110011: data <= 12'h005; 
        10'b0001110100: data <= 12'h001; 
        10'b0001110101: data <= 12'h001; 
        10'b0001110110: data <= 12'h004; 
        10'b0001110111: data <= 12'h003; 
        10'b0001111000: data <= 12'h001; 
        10'b0001111001: data <= 12'hffc; 
        10'b0001111010: data <= 12'h000; 
        10'b0001111011: data <= 12'h001; 
        10'b0001111100: data <= 12'h002; 
        10'b0001111101: data <= 12'h004; 
        10'b0001111110: data <= 12'h005; 
        10'b0001111111: data <= 12'h00a; 
        10'b0010000000: data <= 12'h003; 
        10'b0010000001: data <= 12'hffe; 
        10'b0010000010: data <= 12'hffe; 
        10'b0010000011: data <= 12'h002; 
        10'b0010000100: data <= 12'h005; 
        10'b0010000101: data <= 12'h006; 
        10'b0010000110: data <= 12'h006; 
        10'b0010000111: data <= 12'h007; 
        10'b0010001000: data <= 12'h004; 
        10'b0010001001: data <= 12'h002; 
        10'b0010001010: data <= 12'h002; 
        10'b0010001011: data <= 12'h002; 
        10'b0010001100: data <= 12'h001; 
        10'b0010001101: data <= 12'h004; 
        10'b0010001110: data <= 12'h001; 
        10'b0010001111: data <= 12'h003; 
        10'b0010010000: data <= 12'h001; 
        10'b0010010001: data <= 12'h003; 
        10'b0010010010: data <= 12'h001; 
        10'b0010010011: data <= 12'hfff; 
        10'b0010010100: data <= 12'hff7; 
        10'b0010010101: data <= 12'hff7; 
        10'b0010010110: data <= 12'hffc; 
        10'b0010010111: data <= 12'h000; 
        10'b0010011000: data <= 12'h003; 
        10'b0010011001: data <= 12'h004; 
        10'b0010011010: data <= 12'h007; 
        10'b0010011011: data <= 12'h005; 
        10'b0010011100: data <= 12'h003; 
        10'b0010011101: data <= 12'hffb; 
        10'b0010011110: data <= 12'hfff; 
        10'b0010011111: data <= 12'h001; 
        10'b0010100000: data <= 12'h005; 
        10'b0010100001: data <= 12'h008; 
        10'b0010100010: data <= 12'h00d; 
        10'b0010100011: data <= 12'h008; 
        10'b0010100100: data <= 12'h007; 
        10'b0010100101: data <= 12'hffe; 
        10'b0010100110: data <= 12'h002; 
        10'b0010100111: data <= 12'h001; 
        10'b0010101000: data <= 12'h001; 
        10'b0010101001: data <= 12'h003; 
        10'b0010101010: data <= 12'h001; 
        10'b0010101011: data <= 12'h002; 
        10'b0010101100: data <= 12'h001; 
        10'b0010101101: data <= 12'hfff; 
        10'b0010101110: data <= 12'hffb; 
        10'b0010101111: data <= 12'hffb; 
        10'b0010110000: data <= 12'hff5; 
        10'b0010110001: data <= 12'hff3; 
        10'b0010110010: data <= 12'hff8; 
        10'b0010110011: data <= 12'hffe; 
        10'b0010110100: data <= 12'hffe; 
        10'b0010110101: data <= 12'hffc; 
        10'b0010110110: data <= 12'hffe; 
        10'b0010110111: data <= 12'hff6; 
        10'b0010111000: data <= 12'hff6; 
        10'b0010111001: data <= 12'hff6; 
        10'b0010111010: data <= 12'hffc; 
        10'b0010111011: data <= 12'hffd; 
        10'b0010111100: data <= 12'h005; 
        10'b0010111101: data <= 12'h008; 
        10'b0010111110: data <= 12'h007; 
        10'b0010111111: data <= 12'h006; 
        10'b0011000000: data <= 12'h002; 
        10'b0011000001: data <= 12'hfff; 
        10'b0011000010: data <= 12'h000; 
        10'b0011000011: data <= 12'h002; 
        10'b0011000100: data <= 12'h002; 
        10'b0011000101: data <= 12'h001; 
        10'b0011000110: data <= 12'h001; 
        10'b0011000111: data <= 12'h000; 
        10'b0011001000: data <= 12'h003; 
        10'b0011001001: data <= 12'hfff; 
        10'b0011001010: data <= 12'hffb; 
        10'b0011001011: data <= 12'hff6; 
        10'b0011001100: data <= 12'hff1; 
        10'b0011001101: data <= 12'hfed; 
        10'b0011001110: data <= 12'hff3; 
        10'b0011001111: data <= 12'hffa; 
        10'b0011010000: data <= 12'hffb; 
        10'b0011010001: data <= 12'hff9; 
        10'b0011010010: data <= 12'hff7; 
        10'b0011010011: data <= 12'hff2; 
        10'b0011010100: data <= 12'hff3; 
        10'b0011010101: data <= 12'hff4; 
        10'b0011010110: data <= 12'hff5; 
        10'b0011010111: data <= 12'h000; 
        10'b0011011000: data <= 12'h002; 
        10'b0011011001: data <= 12'h001; 
        10'b0011011010: data <= 12'h001; 
        10'b0011011011: data <= 12'hffc; 
        10'b0011011100: data <= 12'hffa; 
        10'b0011011101: data <= 12'hffe; 
        10'b0011011110: data <= 12'h002; 
        10'b0011011111: data <= 12'h002; 
        10'b0011100000: data <= 12'h002; 
        10'b0011100001: data <= 12'h002; 
        10'b0011100010: data <= 12'h002; 
        10'b0011100011: data <= 12'h004; 
        10'b0011100100: data <= 12'h001; 
        10'b0011100101: data <= 12'h000; 
        10'b0011100110: data <= 12'hffa; 
        10'b0011100111: data <= 12'hff8; 
        10'b0011101000: data <= 12'hfee; 
        10'b0011101001: data <= 12'hfed; 
        10'b0011101010: data <= 12'hfee; 
        10'b0011101011: data <= 12'hff6; 
        10'b0011101100: data <= 12'hffc; 
        10'b0011101101: data <= 12'hffa; 
        10'b0011101110: data <= 12'hffc; 
        10'b0011101111: data <= 12'h002; 
        10'b0011110000: data <= 12'hff8; 
        10'b0011110001: data <= 12'hffd; 
        10'b0011110010: data <= 12'h000; 
        10'b0011110011: data <= 12'h001; 
        10'b0011110100: data <= 12'hffa; 
        10'b0011110101: data <= 12'hffa; 
        10'b0011110110: data <= 12'hff7; 
        10'b0011110111: data <= 12'hff4; 
        10'b0011111000: data <= 12'hff6; 
        10'b0011111001: data <= 12'hffe; 
        10'b0011111010: data <= 12'h004; 
        10'b0011111011: data <= 12'h005; 
        10'b0011111100: data <= 12'h005; 
        10'b0011111101: data <= 12'h001; 
        10'b0011111110: data <= 12'h002; 
        10'b0011111111: data <= 12'h002; 
        10'b0100000000: data <= 12'h000; 
        10'b0100000001: data <= 12'hfff; 
        10'b0100000010: data <= 12'hff9; 
        10'b0100000011: data <= 12'hff9; 
        10'b0100000100: data <= 12'hff4; 
        10'b0100000101: data <= 12'hfee; 
        10'b0100000110: data <= 12'hfef; 
        10'b0100000111: data <= 12'hff9; 
        10'b0100001000: data <= 12'hffb; 
        10'b0100001001: data <= 12'h004; 
        10'b0100001010: data <= 12'h00c; 
        10'b0100001011: data <= 12'h011; 
        10'b0100001100: data <= 12'h006; 
        10'b0100001101: data <= 12'h000; 
        10'b0100001110: data <= 12'hffd; 
        10'b0100001111: data <= 12'hff4; 
        10'b0100010000: data <= 12'hff2; 
        10'b0100010001: data <= 12'hff2; 
        10'b0100010010: data <= 12'hfee; 
        10'b0100010011: data <= 12'hff1; 
        10'b0100010100: data <= 12'hff8; 
        10'b0100010101: data <= 12'h001; 
        10'b0100010110: data <= 12'h004; 
        10'b0100010111: data <= 12'h003; 
        10'b0100011000: data <= 12'h004; 
        10'b0100011001: data <= 12'h005; 
        10'b0100011010: data <= 12'h004; 
        10'b0100011011: data <= 12'h001; 
        10'b0100011100: data <= 12'h003; 
        10'b0100011101: data <= 12'hffc; 
        10'b0100011110: data <= 12'hff9; 
        10'b0100011111: data <= 12'hffd; 
        10'b0100100000: data <= 12'hff7; 
        10'b0100100001: data <= 12'hff7; 
        10'b0100100010: data <= 12'hff9; 
        10'b0100100011: data <= 12'hffb; 
        10'b0100100100: data <= 12'hffd; 
        10'b0100100101: data <= 12'h009; 
        10'b0100100110: data <= 12'h01f; 
        10'b0100100111: data <= 12'h020; 
        10'b0100101000: data <= 12'h00f; 
        10'b0100101001: data <= 12'h000; 
        10'b0100101010: data <= 12'hff7; 
        10'b0100101011: data <= 12'hff5; 
        10'b0100101100: data <= 12'hff3; 
        10'b0100101101: data <= 12'hff4; 
        10'b0100101110: data <= 12'hff5; 
        10'b0100101111: data <= 12'hff9; 
        10'b0100110000: data <= 12'hffe; 
        10'b0100110001: data <= 12'h000; 
        10'b0100110010: data <= 12'h004; 
        10'b0100110011: data <= 12'h002; 
        10'b0100110100: data <= 12'h001; 
        10'b0100110101: data <= 12'h001; 
        10'b0100110110: data <= 12'h003; 
        10'b0100110111: data <= 12'h004; 
        10'b0100111000: data <= 12'h000; 
        10'b0100111001: data <= 12'hfff; 
        10'b0100111010: data <= 12'hfff; 
        10'b0100111011: data <= 12'hffa; 
        10'b0100111100: data <= 12'hffc; 
        10'b0100111101: data <= 12'hffa; 
        10'b0100111110: data <= 12'hff7; 
        10'b0100111111: data <= 12'hff3; 
        10'b0101000000: data <= 12'hfff; 
        10'b0101000001: data <= 12'h010; 
        10'b0101000010: data <= 12'h025; 
        10'b0101000011: data <= 12'h027; 
        10'b0101000100: data <= 12'h00f; 
        10'b0101000101: data <= 12'hffd; 
        10'b0101000110: data <= 12'hffd; 
        10'b0101000111: data <= 12'hff8; 
        10'b0101001000: data <= 12'hff8; 
        10'b0101001001: data <= 12'hff8; 
        10'b0101001010: data <= 12'hff9; 
        10'b0101001011: data <= 12'hffd; 
        10'b0101001100: data <= 12'hfff; 
        10'b0101001101: data <= 12'h003; 
        10'b0101001110: data <= 12'h005; 
        10'b0101001111: data <= 12'h003; 
        10'b0101010000: data <= 12'h001; 
        10'b0101010001: data <= 12'h004; 
        10'b0101010010: data <= 12'h002; 
        10'b0101010011: data <= 12'h001; 
        10'b0101010100: data <= 12'h004; 
        10'b0101010101: data <= 12'hfff; 
        10'b0101010110: data <= 12'hfff; 
        10'b0101010111: data <= 12'hffe; 
        10'b0101011000: data <= 12'hffa; 
        10'b0101011001: data <= 12'hff9; 
        10'b0101011010: data <= 12'hff1; 
        10'b0101011011: data <= 12'hfea; 
        10'b0101011100: data <= 12'hfff; 
        10'b0101011101: data <= 12'h010; 
        10'b0101011110: data <= 12'h02c; 
        10'b0101011111: data <= 12'h01e; 
        10'b0101100000: data <= 12'h006; 
        10'b0101100001: data <= 12'h003; 
        10'b0101100010: data <= 12'hffe; 
        10'b0101100011: data <= 12'hff7; 
        10'b0101100100: data <= 12'hffa; 
        10'b0101100101: data <= 12'hffd; 
        10'b0101100110: data <= 12'hffe; 
        10'b0101100111: data <= 12'hffe; 
        10'b0101101000: data <= 12'h000; 
        10'b0101101001: data <= 12'h004; 
        10'b0101101010: data <= 12'h001; 
        10'b0101101011: data <= 12'h003; 
        10'b0101101100: data <= 12'h000; 
        10'b0101101101: data <= 12'h003; 
        10'b0101101110: data <= 12'h003; 
        10'b0101101111: data <= 12'h003; 
        10'b0101110000: data <= 12'h005; 
        10'b0101110001: data <= 12'h000; 
        10'b0101110010: data <= 12'h000; 
        10'b0101110011: data <= 12'hffe; 
        10'b0101110100: data <= 12'hffd; 
        10'b0101110101: data <= 12'hff4; 
        10'b0101110110: data <= 12'hfe6; 
        10'b0101110111: data <= 12'hfe6; 
        10'b0101111000: data <= 12'h000; 
        10'b0101111001: data <= 12'h00e; 
        10'b0101111010: data <= 12'h024; 
        10'b0101111011: data <= 12'h014; 
        10'b0101111100: data <= 12'h005; 
        10'b0101111101: data <= 12'h003; 
        10'b0101111110: data <= 12'hff8; 
        10'b0101111111: data <= 12'hff4; 
        10'b0110000000: data <= 12'hffc; 
        10'b0110000001: data <= 12'hffe; 
        10'b0110000010: data <= 12'hffe; 
        10'b0110000011: data <= 12'hfff; 
        10'b0110000100: data <= 12'h002; 
        10'b0110000101: data <= 12'h003; 
        10'b0110000110: data <= 12'h004; 
        10'b0110000111: data <= 12'h003; 
        10'b0110001000: data <= 12'h002; 
        10'b0110001001: data <= 12'h005; 
        10'b0110001010: data <= 12'h003; 
        10'b0110001011: data <= 12'h004; 
        10'b0110001100: data <= 12'h004; 
        10'b0110001101: data <= 12'h000; 
        10'b0110001110: data <= 12'h001; 
        10'b0110001111: data <= 12'hfff; 
        10'b0110010000: data <= 12'hff8; 
        10'b0110010001: data <= 12'hff2; 
        10'b0110010010: data <= 12'hfe6; 
        10'b0110010011: data <= 12'hfec; 
        10'b0110010100: data <= 12'h000; 
        10'b0110010101: data <= 12'h00e; 
        10'b0110010110: data <= 12'h01f; 
        10'b0110010111: data <= 12'h014; 
        10'b0110011000: data <= 12'h006; 
        10'b0110011001: data <= 12'hff5; 
        10'b0110011010: data <= 12'hff1; 
        10'b0110011011: data <= 12'hff5; 
        10'b0110011100: data <= 12'hff9; 
        10'b0110011101: data <= 12'hffe; 
        10'b0110011110: data <= 12'hffe; 
        10'b0110011111: data <= 12'hfff; 
        10'b0110100000: data <= 12'h003; 
        10'b0110100001: data <= 12'h001; 
        10'b0110100010: data <= 12'h001; 
        10'b0110100011: data <= 12'h003; 
        10'b0110100100: data <= 12'h005; 
        10'b0110100101: data <= 12'h001; 
        10'b0110100110: data <= 12'h003; 
        10'b0110100111: data <= 12'h002; 
        10'b0110101000: data <= 12'h001; 
        10'b0110101001: data <= 12'h003; 
        10'b0110101010: data <= 12'hffd; 
        10'b0110101011: data <= 12'hffd; 
        10'b0110101100: data <= 12'hffb; 
        10'b0110101101: data <= 12'hff1; 
        10'b0110101110: data <= 12'hfef; 
        10'b0110101111: data <= 12'hffc; 
        10'b0110110000: data <= 12'h006; 
        10'b0110110001: data <= 12'h014; 
        10'b0110110010: data <= 12'h021; 
        10'b0110110011: data <= 12'h00c; 
        10'b0110110100: data <= 12'h002; 
        10'b0110110101: data <= 12'hfeb; 
        10'b0110110110: data <= 12'hfee; 
        10'b0110110111: data <= 12'hff5; 
        10'b0110111000: data <= 12'hff9; 
        10'b0110111001: data <= 12'hffb; 
        10'b0110111010: data <= 12'hfff; 
        10'b0110111011: data <= 12'h000; 
        10'b0110111100: data <= 12'h002; 
        10'b0110111101: data <= 12'h002; 
        10'b0110111110: data <= 12'h005; 
        10'b0110111111: data <= 12'h001; 
        10'b0111000000: data <= 12'h005; 
        10'b0111000001: data <= 12'h002; 
        10'b0111000010: data <= 12'h004; 
        10'b0111000011: data <= 12'h003; 
        10'b0111000100: data <= 12'h001; 
        10'b0111000101: data <= 12'hffe; 
        10'b0111000110: data <= 12'hffc; 
        10'b0111000111: data <= 12'hffb; 
        10'b0111001000: data <= 12'hff4; 
        10'b0111001001: data <= 12'hff9; 
        10'b0111001010: data <= 12'hffa; 
        10'b0111001011: data <= 12'hffd; 
        10'b0111001100: data <= 12'hfff; 
        10'b0111001101: data <= 12'h01a; 
        10'b0111001110: data <= 12'h01f; 
        10'b0111001111: data <= 12'h002; 
        10'b0111010000: data <= 12'hff6; 
        10'b0111010001: data <= 12'hfea; 
        10'b0111010010: data <= 12'hfee; 
        10'b0111010011: data <= 12'hff4; 
        10'b0111010100: data <= 12'hff7; 
        10'b0111010101: data <= 12'hffc; 
        10'b0111010110: data <= 12'hffc; 
        10'b0111010111: data <= 12'h000; 
        10'b0111011000: data <= 12'hffe; 
        10'b0111011001: data <= 12'h000; 
        10'b0111011010: data <= 12'h001; 
        10'b0111011011: data <= 12'h002; 
        10'b0111011100: data <= 12'h002; 
        10'b0111011101: data <= 12'h005; 
        10'b0111011110: data <= 12'h001; 
        10'b0111011111: data <= 12'h005; 
        10'b0111100000: data <= 12'h003; 
        10'b0111100001: data <= 12'hffd; 
        10'b0111100010: data <= 12'hff6; 
        10'b0111100011: data <= 12'hff5; 
        10'b0111100100: data <= 12'hff8; 
        10'b0111100101: data <= 12'hffb; 
        10'b0111100110: data <= 12'h003; 
        10'b0111100111: data <= 12'h000; 
        10'b0111101000: data <= 12'h008; 
        10'b0111101001: data <= 12'h01e; 
        10'b0111101010: data <= 12'h019; 
        10'b0111101011: data <= 12'hffb; 
        10'b0111101100: data <= 12'hfee; 
        10'b0111101101: data <= 12'hfea; 
        10'b0111101110: data <= 12'hfee; 
        10'b0111101111: data <= 12'hff4; 
        10'b0111110000: data <= 12'hffc; 
        10'b0111110001: data <= 12'hffe; 
        10'b0111110010: data <= 12'hffe; 
        10'b0111110011: data <= 12'hffe; 
        10'b0111110100: data <= 12'hffc; 
        10'b0111110101: data <= 12'h001; 
        10'b0111110110: data <= 12'h003; 
        10'b0111110111: data <= 12'h003; 
        10'b0111111000: data <= 12'h003; 
        10'b0111111001: data <= 12'h003; 
        10'b0111111010: data <= 12'h002; 
        10'b0111111011: data <= 12'h004; 
        10'b0111111100: data <= 12'h002; 
        10'b0111111101: data <= 12'hffc; 
        10'b0111111110: data <= 12'hff6; 
        10'b0111111111: data <= 12'hff6; 
        10'b1000000000: data <= 12'hffc; 
        10'b1000000001: data <= 12'h004; 
        10'b1000000010: data <= 12'h003; 
        10'b1000000011: data <= 12'h005; 
        10'b1000000100: data <= 12'h00e; 
        10'b1000000101: data <= 12'h016; 
        10'b1000000110: data <= 12'h00f; 
        10'b1000000111: data <= 12'hff6; 
        10'b1000001000: data <= 12'hff0; 
        10'b1000001001: data <= 12'hff2; 
        10'b1000001010: data <= 12'hff4; 
        10'b1000001011: data <= 12'hff8; 
        10'b1000001100: data <= 12'hffc; 
        10'b1000001101: data <= 12'hff9; 
        10'b1000001110: data <= 12'hffd; 
        10'b1000001111: data <= 12'hffb; 
        10'b1000010000: data <= 12'hffd; 
        10'b1000010001: data <= 12'h003; 
        10'b1000010010: data <= 12'h004; 
        10'b1000010011: data <= 12'h004; 
        10'b1000010100: data <= 12'h005; 
        10'b1000010101: data <= 12'h003; 
        10'b1000010110: data <= 12'h003; 
        10'b1000010111: data <= 12'h004; 
        10'b1000011000: data <= 12'h000; 
        10'b1000011001: data <= 12'hffa; 
        10'b1000011010: data <= 12'hff3; 
        10'b1000011011: data <= 12'hff7; 
        10'b1000011100: data <= 12'hffc; 
        10'b1000011101: data <= 12'h002; 
        10'b1000011110: data <= 12'h001; 
        10'b1000011111: data <= 12'h001; 
        10'b1000100000: data <= 12'h002; 
        10'b1000100001: data <= 12'h00a; 
        10'b1000100010: data <= 12'h002; 
        10'b1000100011: data <= 12'hff8; 
        10'b1000100100: data <= 12'hff9; 
        10'b1000100101: data <= 12'hffa; 
        10'b1000100110: data <= 12'hff8; 
        10'b1000100111: data <= 12'hffa; 
        10'b1000101000: data <= 12'hff7; 
        10'b1000101001: data <= 12'hff9; 
        10'b1000101010: data <= 12'hffc; 
        10'b1000101011: data <= 12'hffc; 
        10'b1000101100: data <= 12'h000; 
        10'b1000101101: data <= 12'h001; 
        10'b1000101110: data <= 12'h002; 
        10'b1000101111: data <= 12'h001; 
        10'b1000110000: data <= 12'h001; 
        10'b1000110001: data <= 12'h005; 
        10'b1000110010: data <= 12'h003; 
        10'b1000110011: data <= 12'h002; 
        10'b1000110100: data <= 12'hfff; 
        10'b1000110101: data <= 12'hffc; 
        10'b1000110110: data <= 12'hfff; 
        10'b1000110111: data <= 12'hffd; 
        10'b1000111000: data <= 12'h000; 
        10'b1000111001: data <= 12'h001; 
        10'b1000111010: data <= 12'hffd; 
        10'b1000111011: data <= 12'hfff; 
        10'b1000111100: data <= 12'hffb; 
        10'b1000111101: data <= 12'hffe; 
        10'b1000111110: data <= 12'hfff; 
        10'b1000111111: data <= 12'h000; 
        10'b1001000000: data <= 12'h005; 
        10'b1001000001: data <= 12'h002; 
        10'b1001000010: data <= 12'hffe; 
        10'b1001000011: data <= 12'hff9; 
        10'b1001000100: data <= 12'hff7; 
        10'b1001000101: data <= 12'hff8; 
        10'b1001000110: data <= 12'hffa; 
        10'b1001000111: data <= 12'hfff; 
        10'b1001001000: data <= 12'h001; 
        10'b1001001001: data <= 12'h004; 
        10'b1001001010: data <= 12'h002; 
        10'b1001001011: data <= 12'h005; 
        10'b1001001100: data <= 12'h003; 
        10'b1001001101: data <= 12'h002; 
        10'b1001001110: data <= 12'h003; 
        10'b1001001111: data <= 12'h003; 
        10'b1001010000: data <= 12'h003; 
        10'b1001010001: data <= 12'h007; 
        10'b1001010010: data <= 12'h006; 
        10'b1001010011: data <= 12'h003; 
        10'b1001010100: data <= 12'h000; 
        10'b1001010101: data <= 12'hffe; 
        10'b1001010110: data <= 12'h000; 
        10'b1001010111: data <= 12'hffc; 
        10'b1001011000: data <= 12'hff6; 
        10'b1001011001: data <= 12'hff5; 
        10'b1001011010: data <= 12'hfff; 
        10'b1001011011: data <= 12'h003; 
        10'b1001011100: data <= 12'h005; 
        10'b1001011101: data <= 12'h006; 
        10'b1001011110: data <= 12'h004; 
        10'b1001011111: data <= 12'hff9; 
        10'b1001100000: data <= 12'hff9; 
        10'b1001100001: data <= 12'hff8; 
        10'b1001100010: data <= 12'hffb; 
        10'b1001100011: data <= 12'hffd; 
        10'b1001100100: data <= 12'h001; 
        10'b1001100101: data <= 12'h002; 
        10'b1001100110: data <= 12'h000; 
        10'b1001100111: data <= 12'h001; 
        10'b1001101000: data <= 12'h003; 
        10'b1001101001: data <= 12'h003; 
        10'b1001101010: data <= 12'h003; 
        10'b1001101011: data <= 12'h001; 
        10'b1001101100: data <= 12'h006; 
        10'b1001101101: data <= 12'h00e; 
        10'b1001101110: data <= 12'h00f; 
        10'b1001101111: data <= 12'h009; 
        10'b1001110000: data <= 12'h001; 
        10'b1001110001: data <= 12'hfff; 
        10'b1001110010: data <= 12'hffd; 
        10'b1001110011: data <= 12'hff2; 
        10'b1001110100: data <= 12'hfe9; 
        10'b1001110101: data <= 12'hfef; 
        10'b1001110110: data <= 12'h000; 
        10'b1001110111: data <= 12'h003; 
        10'b1001111000: data <= 12'h00d; 
        10'b1001111001: data <= 12'h015; 
        10'b1001111010: data <= 12'h009; 
        10'b1001111011: data <= 12'h002; 
        10'b1001111100: data <= 12'hffb; 
        10'b1001111101: data <= 12'hffc; 
        10'b1001111110: data <= 12'h000; 
        10'b1001111111: data <= 12'h001; 
        10'b1010000000: data <= 12'h000; 
        10'b1010000001: data <= 12'h002; 
        10'b1010000010: data <= 12'h005; 
        10'b1010000011: data <= 12'h002; 
        10'b1010000100: data <= 12'h004; 
        10'b1010000101: data <= 12'h003; 
        10'b1010000110: data <= 12'h003; 
        10'b1010000111: data <= 12'h002; 
        10'b1010001000: data <= 12'h006; 
        10'b1010001001: data <= 12'h00c; 
        10'b1010001010: data <= 12'h00d; 
        10'b1010001011: data <= 12'h006; 
        10'b1010001100: data <= 12'h002; 
        10'b1010001101: data <= 12'hffd; 
        10'b1010001110: data <= 12'hffe; 
        10'b1010001111: data <= 12'hff8; 
        10'b1010010000: data <= 12'hffb; 
        10'b1010010001: data <= 12'hffb; 
        10'b1010010010: data <= 12'hff9; 
        10'b1010010011: data <= 12'h003; 
        10'b1010010100: data <= 12'h00f; 
        10'b1010010101: data <= 12'h012; 
        10'b1010010110: data <= 12'h008; 
        10'b1010010111: data <= 12'hfff; 
        10'b1010011000: data <= 12'hffd; 
        10'b1010011001: data <= 12'hffb; 
        10'b1010011010: data <= 12'hffe; 
        10'b1010011011: data <= 12'hffe; 
        10'b1010011100: data <= 12'h001; 
        10'b1010011101: data <= 12'h001; 
        10'b1010011110: data <= 12'h001; 
        10'b1010011111: data <= 12'h000; 
        10'b1010100000: data <= 12'h001; 
        10'b1010100001: data <= 12'h001; 
        10'b1010100010: data <= 12'h002; 
        10'b1010100011: data <= 12'h001; 
        10'b1010100100: data <= 12'h003; 
        10'b1010100101: data <= 12'h005; 
        10'b1010100110: data <= 12'h006; 
        10'b1010100111: data <= 12'hffe; 
        10'b1010101000: data <= 12'hff8; 
        10'b1010101001: data <= 12'hff8; 
        10'b1010101010: data <= 12'hff2; 
        10'b1010101011: data <= 12'hff2; 
        10'b1010101100: data <= 12'hff4; 
        10'b1010101101: data <= 12'hff6; 
        10'b1010101110: data <= 12'hff6; 
        10'b1010101111: data <= 12'hff6; 
        10'b1010110000: data <= 12'hffd; 
        10'b1010110001: data <= 12'h001; 
        10'b1010110010: data <= 12'h002; 
        10'b1010110011: data <= 12'h003; 
        10'b1010110100: data <= 12'h003; 
        10'b1010110101: data <= 12'h001; 
        10'b1010110110: data <= 12'h001; 
        10'b1010110111: data <= 12'h004; 
        10'b1010111000: data <= 12'h001; 
        10'b1010111001: data <= 12'h002; 
        10'b1010111010: data <= 12'h004; 
        10'b1010111011: data <= 12'h001; 
        10'b1010111100: data <= 12'h005; 
        10'b1010111101: data <= 12'h002; 
        10'b1010111110: data <= 12'h002; 
        10'b1010111111: data <= 12'h003; 
        10'b1011000000: data <= 12'h004; 
        10'b1011000001: data <= 12'h003; 
        10'b1011000010: data <= 12'h000; 
        10'b1011000011: data <= 12'hffe; 
        10'b1011000100: data <= 12'hfff; 
        10'b1011000101: data <= 12'hffe; 
        10'b1011000110: data <= 12'hff8; 
        10'b1011000111: data <= 12'hff6; 
        10'b1011001000: data <= 12'hff9; 
        10'b1011001001: data <= 12'hff6; 
        10'b1011001010: data <= 12'hffa; 
        10'b1011001011: data <= 12'hff8; 
        10'b1011001100: data <= 12'hffc; 
        10'b1011001101: data <= 12'hfff; 
        10'b1011001110: data <= 12'h002; 
        10'b1011001111: data <= 12'h003; 
        10'b1011010000: data <= 12'h000; 
        10'b1011010001: data <= 12'h003; 
        10'b1011010010: data <= 12'h002; 
        10'b1011010011: data <= 12'h004; 
        10'b1011010100: data <= 12'h001; 
        10'b1011010101: data <= 12'h001; 
        10'b1011010110: data <= 12'h002; 
        10'b1011010111: data <= 12'h002; 
        10'b1011011000: data <= 12'h002; 
        10'b1011011001: data <= 12'h003; 
        10'b1011011010: data <= 12'h003; 
        10'b1011011011: data <= 12'h001; 
        10'b1011011100: data <= 12'h003; 
        10'b1011011101: data <= 12'h004; 
        10'b1011011110: data <= 12'h003; 
        10'b1011011111: data <= 12'h003; 
        10'b1011100000: data <= 12'h004; 
        10'b1011100001: data <= 12'h003; 
        10'b1011100010: data <= 12'h000; 
        10'b1011100011: data <= 12'h003; 
        10'b1011100100: data <= 12'h002; 
        10'b1011100101: data <= 12'h001; 
        10'b1011100110: data <= 12'h000; 
        10'b1011100111: data <= 12'h001; 
        10'b1011101000: data <= 12'h003; 
        10'b1011101001: data <= 12'h004; 
        10'b1011101010: data <= 12'h003; 
        10'b1011101011: data <= 12'h001; 
        10'b1011101100: data <= 12'h003; 
        10'b1011101101: data <= 12'h003; 
        10'b1011101110: data <= 12'h003; 
        10'b1011101111: data <= 12'h001; 
        10'b1011110000: data <= 12'h001; 
        10'b1011110001: data <= 12'h003; 
        10'b1011110010: data <= 12'h004; 
        10'b1011110011: data <= 12'h004; 
        10'b1011110100: data <= 12'h004; 
        10'b1011110101: data <= 12'h005; 
        10'b1011110110: data <= 12'h001; 
        10'b1011110111: data <= 12'h003; 
        10'b1011111000: data <= 12'h005; 
        10'b1011111001: data <= 12'h004; 
        10'b1011111010: data <= 12'h004; 
        10'b1011111011: data <= 12'h004; 
        10'b1011111100: data <= 12'h004; 
        10'b1011111101: data <= 12'h002; 
        10'b1011111110: data <= 12'h004; 
        10'b1011111111: data <= 12'h004; 
        10'b1100000000: data <= 12'h000; 
        10'b1100000001: data <= 12'h001; 
        10'b1100000010: data <= 12'h005; 
        10'b1100000011: data <= 12'h003; 
        10'b1100000100: data <= 12'h003; 
        10'b1100000101: data <= 12'h000; 
        10'b1100000110: data <= 12'h002; 
        10'b1100000111: data <= 12'h001; 
        10'b1100001000: data <= 12'h001; 
        10'b1100001001: data <= 12'h002; 
        10'b1100001010: data <= 12'h003; 
        10'b1100001011: data <= 12'h004; 
        10'b1100001100: data <= 12'h004; 
        10'b1100001101: data <= 12'h004; 
        10'b1100001110: data <= 12'h004; 
        10'b1100001111: data <= 12'h001; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 7) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 13'h0008; 
        10'b0000000001: data <= 13'h0004; 
        10'b0000000010: data <= 13'h0004; 
        10'b0000000011: data <= 13'h0002; 
        10'b0000000100: data <= 13'h0007; 
        10'b0000000101: data <= 13'h0007; 
        10'b0000000110: data <= 13'h0007; 
        10'b0000000111: data <= 13'h0002; 
        10'b0000001000: data <= 13'h0006; 
        10'b0000001001: data <= 13'h0002; 
        10'b0000001010: data <= 13'h0006; 
        10'b0000001011: data <= 13'h0005; 
        10'b0000001100: data <= 13'h0007; 
        10'b0000001101: data <= 13'h0009; 
        10'b0000001110: data <= 13'h0008; 
        10'b0000001111: data <= 13'h0005; 
        10'b0000010000: data <= 13'h0006; 
        10'b0000010001: data <= 13'h0002; 
        10'b0000010010: data <= 13'h0009; 
        10'b0000010011: data <= 13'h0009; 
        10'b0000010100: data <= 13'h0005; 
        10'b0000010101: data <= 13'h0007; 
        10'b0000010110: data <= 13'h0005; 
        10'b0000010111: data <= 13'h0008; 
        10'b0000011000: data <= 13'h0003; 
        10'b0000011001: data <= 13'h0009; 
        10'b0000011010: data <= 13'h0005; 
        10'b0000011011: data <= 13'h0008; 
        10'b0000011100: data <= 13'h0001; 
        10'b0000011101: data <= 13'h0008; 
        10'b0000011110: data <= 13'h0002; 
        10'b0000011111: data <= 13'h0006; 
        10'b0000100000: data <= 13'h0005; 
        10'b0000100001: data <= 13'h0002; 
        10'b0000100010: data <= 13'h0003; 
        10'b0000100011: data <= 13'h0008; 
        10'b0000100100: data <= 13'h0007; 
        10'b0000100101: data <= 13'h0006; 
        10'b0000100110: data <= 13'h0006; 
        10'b0000100111: data <= 13'h0004; 
        10'b0000101000: data <= 13'h0007; 
        10'b0000101001: data <= 13'h0008; 
        10'b0000101010: data <= 13'h000a; 
        10'b0000101011: data <= 13'h0005; 
        10'b0000101100: data <= 13'h0004; 
        10'b0000101101: data <= 13'h0008; 
        10'b0000101110: data <= 13'h0005; 
        10'b0000101111: data <= 13'h0004; 
        10'b0000110000: data <= 13'h0009; 
        10'b0000110001: data <= 13'h0008; 
        10'b0000110010: data <= 13'h0003; 
        10'b0000110011: data <= 13'h0009; 
        10'b0000110100: data <= 13'h000a; 
        10'b0000110101: data <= 13'h0005; 
        10'b0000110110: data <= 13'h0008; 
        10'b0000110111: data <= 13'h0007; 
        10'b0000111000: data <= 13'h0008; 
        10'b0000111001: data <= 13'h0006; 
        10'b0000111010: data <= 13'h000a; 
        10'b0000111011: data <= 13'h0002; 
        10'b0000111100: data <= 13'h0002; 
        10'b0000111101: data <= 13'h0006; 
        10'b0000111110: data <= 13'h0005; 
        10'b0000111111: data <= 13'h0005; 
        10'b0001000000: data <= 13'h0003; 
        10'b0001000001: data <= 13'h0005; 
        10'b0001000010: data <= 13'h0000; 
        10'b0001000011: data <= 13'h0003; 
        10'b0001000100: data <= 13'h0000; 
        10'b0001000101: data <= 13'h0002; 
        10'b0001000110: data <= 13'h0005; 
        10'b0001000111: data <= 13'h0008; 
        10'b0001001000: data <= 13'h0006; 
        10'b0001001001: data <= 13'h0000; 
        10'b0001001010: data <= 13'h0006; 
        10'b0001001011: data <= 13'h0004; 
        10'b0001001100: data <= 13'h0008; 
        10'b0001001101: data <= 13'h0003; 
        10'b0001001110: data <= 13'h0009; 
        10'b0001001111: data <= 13'h0006; 
        10'b0001010000: data <= 13'h0007; 
        10'b0001010001: data <= 13'h0001; 
        10'b0001010010: data <= 13'h0007; 
        10'b0001010011: data <= 13'h0008; 
        10'b0001010100: data <= 13'h0003; 
        10'b0001010101: data <= 13'h0003; 
        10'b0001010110: data <= 13'h0006; 
        10'b0001010111: data <= 13'h0005; 
        10'b0001011000: data <= 13'h0009; 
        10'b0001011001: data <= 13'h0005; 
        10'b0001011010: data <= 13'h0001; 
        10'b0001011011: data <= 13'h0009; 
        10'b0001011100: data <= 13'h1fff; 
        10'b0001011101: data <= 13'h1ffe; 
        10'b0001011110: data <= 13'h1ffe; 
        10'b0001011111: data <= 13'h1ffb; 
        10'b0001100000: data <= 13'h1ffe; 
        10'b0001100001: data <= 13'h0001; 
        10'b0001100010: data <= 13'h0004; 
        10'b0001100011: data <= 13'h0007; 
        10'b0001100100: data <= 13'h1ffc; 
        10'b0001100101: data <= 13'h1fff; 
        10'b0001100110: data <= 13'h0000; 
        10'b0001100111: data <= 13'h1ffa; 
        10'b0001101000: data <= 13'h1fff; 
        10'b0001101001: data <= 13'h0002; 
        10'b0001101010: data <= 13'h0006; 
        10'b0001101011: data <= 13'h0006; 
        10'b0001101100: data <= 13'h1fff; 
        10'b0001101101: data <= 13'h0008; 
        10'b0001101110: data <= 13'h0003; 
        10'b0001101111: data <= 13'h0009; 
        10'b0001110000: data <= 13'h0007; 
        10'b0001110001: data <= 13'h0004; 
        10'b0001110010: data <= 13'h0009; 
        10'b0001110011: data <= 13'h0009; 
        10'b0001110100: data <= 13'h0001; 
        10'b0001110101: data <= 13'h0002; 
        10'b0001110110: data <= 13'h0008; 
        10'b0001110111: data <= 13'h0005; 
        10'b0001111000: data <= 13'h0002; 
        10'b0001111001: data <= 13'h1ff8; 
        10'b0001111010: data <= 13'h0001; 
        10'b0001111011: data <= 13'h0003; 
        10'b0001111100: data <= 13'h0005; 
        10'b0001111101: data <= 13'h0008; 
        10'b0001111110: data <= 13'h000a; 
        10'b0001111111: data <= 13'h0014; 
        10'b0010000000: data <= 13'h0005; 
        10'b0010000001: data <= 13'h1ffc; 
        10'b0010000010: data <= 13'h1ffb; 
        10'b0010000011: data <= 13'h0003; 
        10'b0010000100: data <= 13'h000b; 
        10'b0010000101: data <= 13'h000c; 
        10'b0010000110: data <= 13'h000c; 
        10'b0010000111: data <= 13'h000e; 
        10'b0010001000: data <= 13'h0007; 
        10'b0010001001: data <= 13'h0004; 
        10'b0010001010: data <= 13'h0003; 
        10'b0010001011: data <= 13'h0003; 
        10'b0010001100: data <= 13'h0001; 
        10'b0010001101: data <= 13'h0008; 
        10'b0010001110: data <= 13'h0002; 
        10'b0010001111: data <= 13'h0006; 
        10'b0010010000: data <= 13'h0001; 
        10'b0010010001: data <= 13'h0005; 
        10'b0010010010: data <= 13'h0002; 
        10'b0010010011: data <= 13'h1ffe; 
        10'b0010010100: data <= 13'h1fee; 
        10'b0010010101: data <= 13'h1fee; 
        10'b0010010110: data <= 13'h1ff8; 
        10'b0010010111: data <= 13'h0000; 
        10'b0010011000: data <= 13'h0007; 
        10'b0010011001: data <= 13'h0008; 
        10'b0010011010: data <= 13'h000d; 
        10'b0010011011: data <= 13'h000a; 
        10'b0010011100: data <= 13'h0006; 
        10'b0010011101: data <= 13'h1ff6; 
        10'b0010011110: data <= 13'h1fff; 
        10'b0010011111: data <= 13'h0002; 
        10'b0010100000: data <= 13'h000a; 
        10'b0010100001: data <= 13'h0010; 
        10'b0010100010: data <= 13'h001a; 
        10'b0010100011: data <= 13'h0010; 
        10'b0010100100: data <= 13'h000d; 
        10'b0010100101: data <= 13'h1ffd; 
        10'b0010100110: data <= 13'h0004; 
        10'b0010100111: data <= 13'h0002; 
        10'b0010101000: data <= 13'h0002; 
        10'b0010101001: data <= 13'h0006; 
        10'b0010101010: data <= 13'h0001; 
        10'b0010101011: data <= 13'h0005; 
        10'b0010101100: data <= 13'h0001; 
        10'b0010101101: data <= 13'h1ffd; 
        10'b0010101110: data <= 13'h1ff6; 
        10'b0010101111: data <= 13'h1ff6; 
        10'b0010110000: data <= 13'h1fea; 
        10'b0010110001: data <= 13'h1fe5; 
        10'b0010110010: data <= 13'h1fef; 
        10'b0010110011: data <= 13'h1ffc; 
        10'b0010110100: data <= 13'h1ffc; 
        10'b0010110101: data <= 13'h1ff8; 
        10'b0010110110: data <= 13'h1ffc; 
        10'b0010110111: data <= 13'h1fed; 
        10'b0010111000: data <= 13'h1feb; 
        10'b0010111001: data <= 13'h1feb; 
        10'b0010111010: data <= 13'h1ff7; 
        10'b0010111011: data <= 13'h1ffa; 
        10'b0010111100: data <= 13'h000a; 
        10'b0010111101: data <= 13'h0010; 
        10'b0010111110: data <= 13'h000f; 
        10'b0010111111: data <= 13'h000d; 
        10'b0011000000: data <= 13'h0003; 
        10'b0011000001: data <= 13'h1ffd; 
        10'b0011000010: data <= 13'h0000; 
        10'b0011000011: data <= 13'h0005; 
        10'b0011000100: data <= 13'h0004; 
        10'b0011000101: data <= 13'h0002; 
        10'b0011000110: data <= 13'h0003; 
        10'b0011000111: data <= 13'h0001; 
        10'b0011001000: data <= 13'h0006; 
        10'b0011001001: data <= 13'h1fff; 
        10'b0011001010: data <= 13'h1ff7; 
        10'b0011001011: data <= 13'h1fed; 
        10'b0011001100: data <= 13'h1fe2; 
        10'b0011001101: data <= 13'h1fda; 
        10'b0011001110: data <= 13'h1fe6; 
        10'b0011001111: data <= 13'h1ff5; 
        10'b0011010000: data <= 13'h1ff6; 
        10'b0011010001: data <= 13'h1ff1; 
        10'b0011010010: data <= 13'h1fee; 
        10'b0011010011: data <= 13'h1fe3; 
        10'b0011010100: data <= 13'h1fe7; 
        10'b0011010101: data <= 13'h1fe8; 
        10'b0011010110: data <= 13'h1feb; 
        10'b0011010111: data <= 13'h1fff; 
        10'b0011011000: data <= 13'h0004; 
        10'b0011011001: data <= 13'h0003; 
        10'b0011011010: data <= 13'h0003; 
        10'b0011011011: data <= 13'h1ff8; 
        10'b0011011100: data <= 13'h1ff5; 
        10'b0011011101: data <= 13'h1ffc; 
        10'b0011011110: data <= 13'h0004; 
        10'b0011011111: data <= 13'h0004; 
        10'b0011100000: data <= 13'h0005; 
        10'b0011100001: data <= 13'h0004; 
        10'b0011100010: data <= 13'h0004; 
        10'b0011100011: data <= 13'h0008; 
        10'b0011100100: data <= 13'h0003; 
        10'b0011100101: data <= 13'h0000; 
        10'b0011100110: data <= 13'h1ff5; 
        10'b0011100111: data <= 13'h1fef; 
        10'b0011101000: data <= 13'h1fdd; 
        10'b0011101001: data <= 13'h1fda; 
        10'b0011101010: data <= 13'h1fdc; 
        10'b0011101011: data <= 13'h1fed; 
        10'b0011101100: data <= 13'h1ff7; 
        10'b0011101101: data <= 13'h1ff5; 
        10'b0011101110: data <= 13'h1ff7; 
        10'b0011101111: data <= 13'h0004; 
        10'b0011110000: data <= 13'h1ff0; 
        10'b0011110001: data <= 13'h1ffb; 
        10'b0011110010: data <= 13'h1fff; 
        10'b0011110011: data <= 13'h0002; 
        10'b0011110100: data <= 13'h1ff4; 
        10'b0011110101: data <= 13'h1ff4; 
        10'b0011110110: data <= 13'h1fed; 
        10'b0011110111: data <= 13'h1fe8; 
        10'b0011111000: data <= 13'h1fed; 
        10'b0011111001: data <= 13'h1ffb; 
        10'b0011111010: data <= 13'h0007; 
        10'b0011111011: data <= 13'h0009; 
        10'b0011111100: data <= 13'h000a; 
        10'b0011111101: data <= 13'h0002; 
        10'b0011111110: data <= 13'h0004; 
        10'b0011111111: data <= 13'h0003; 
        10'b0100000000: data <= 13'h1fff; 
        10'b0100000001: data <= 13'h1fff; 
        10'b0100000010: data <= 13'h1ff2; 
        10'b0100000011: data <= 13'h1ff3; 
        10'b0100000100: data <= 13'h1fe8; 
        10'b0100000101: data <= 13'h1fdb; 
        10'b0100000110: data <= 13'h1fde; 
        10'b0100000111: data <= 13'h1ff3; 
        10'b0100001000: data <= 13'h1ff6; 
        10'b0100001001: data <= 13'h0008; 
        10'b0100001010: data <= 13'h0018; 
        10'b0100001011: data <= 13'h0022; 
        10'b0100001100: data <= 13'h000d; 
        10'b0100001101: data <= 13'h1fff; 
        10'b0100001110: data <= 13'h1ffa; 
        10'b0100001111: data <= 13'h1fe9; 
        10'b0100010000: data <= 13'h1fe4; 
        10'b0100010001: data <= 13'h1fe4; 
        10'b0100010010: data <= 13'h1fdd; 
        10'b0100010011: data <= 13'h1fe1; 
        10'b0100010100: data <= 13'h1ff0; 
        10'b0100010101: data <= 13'h0002; 
        10'b0100010110: data <= 13'h0008; 
        10'b0100010111: data <= 13'h0006; 
        10'b0100011000: data <= 13'h0009; 
        10'b0100011001: data <= 13'h000a; 
        10'b0100011010: data <= 13'h0008; 
        10'b0100011011: data <= 13'h0001; 
        10'b0100011100: data <= 13'h0007; 
        10'b0100011101: data <= 13'h1ff8; 
        10'b0100011110: data <= 13'h1ff3; 
        10'b0100011111: data <= 13'h1ffa; 
        10'b0100100000: data <= 13'h1fed; 
        10'b0100100001: data <= 13'h1fed; 
        10'b0100100010: data <= 13'h1ff2; 
        10'b0100100011: data <= 13'h1ff7; 
        10'b0100100100: data <= 13'h1ffa; 
        10'b0100100101: data <= 13'h0013; 
        10'b0100100110: data <= 13'h003d; 
        10'b0100100111: data <= 13'h0041; 
        10'b0100101000: data <= 13'h001f; 
        10'b0100101001: data <= 13'h1fff; 
        10'b0100101010: data <= 13'h1fee; 
        10'b0100101011: data <= 13'h1fea; 
        10'b0100101100: data <= 13'h1fe5; 
        10'b0100101101: data <= 13'h1fe8; 
        10'b0100101110: data <= 13'h1fe9; 
        10'b0100101111: data <= 13'h1ff2; 
        10'b0100110000: data <= 13'h1ffb; 
        10'b0100110001: data <= 13'h1fff; 
        10'b0100110010: data <= 13'h0008; 
        10'b0100110011: data <= 13'h0003; 
        10'b0100110100: data <= 13'h0002; 
        10'b0100110101: data <= 13'h0001; 
        10'b0100110110: data <= 13'h0007; 
        10'b0100110111: data <= 13'h0007; 
        10'b0100111000: data <= 13'h0000; 
        10'b0100111001: data <= 13'h1ffe; 
        10'b0100111010: data <= 13'h1fff; 
        10'b0100111011: data <= 13'h1ff4; 
        10'b0100111100: data <= 13'h1ff8; 
        10'b0100111101: data <= 13'h1ff4; 
        10'b0100111110: data <= 13'h1fef; 
        10'b0100111111: data <= 13'h1fe6; 
        10'b0101000000: data <= 13'h1ffd; 
        10'b0101000001: data <= 13'h0020; 
        10'b0101000010: data <= 13'h004a; 
        10'b0101000011: data <= 13'h004f; 
        10'b0101000100: data <= 13'h001d; 
        10'b0101000101: data <= 13'h1ffa; 
        10'b0101000110: data <= 13'h1ffa; 
        10'b0101000111: data <= 13'h1ff1; 
        10'b0101001000: data <= 13'h1ff0; 
        10'b0101001001: data <= 13'h1ff1; 
        10'b0101001010: data <= 13'h1ff2; 
        10'b0101001011: data <= 13'h1ff9; 
        10'b0101001100: data <= 13'h1ffd; 
        10'b0101001101: data <= 13'h0007; 
        10'b0101001110: data <= 13'h0009; 
        10'b0101001111: data <= 13'h0006; 
        10'b0101010000: data <= 13'h0001; 
        10'b0101010001: data <= 13'h0009; 
        10'b0101010010: data <= 13'h0004; 
        10'b0101010011: data <= 13'h0003; 
        10'b0101010100: data <= 13'h0009; 
        10'b0101010101: data <= 13'h1ffe; 
        10'b0101010110: data <= 13'h1ffd; 
        10'b0101010111: data <= 13'h1ffc; 
        10'b0101011000: data <= 13'h1ff5; 
        10'b0101011001: data <= 13'h1ff1; 
        10'b0101011010: data <= 13'h1fe1; 
        10'b0101011011: data <= 13'h1fd5; 
        10'b0101011100: data <= 13'h1fff; 
        10'b0101011101: data <= 13'h0021; 
        10'b0101011110: data <= 13'h0057; 
        10'b0101011111: data <= 13'h003d; 
        10'b0101100000: data <= 13'h000c; 
        10'b0101100001: data <= 13'h0006; 
        10'b0101100010: data <= 13'h1ffc; 
        10'b0101100011: data <= 13'h1fee; 
        10'b0101100100: data <= 13'h1ff5; 
        10'b0101100101: data <= 13'h1ffb; 
        10'b0101100110: data <= 13'h1ffd; 
        10'b0101100111: data <= 13'h1ffc; 
        10'b0101101000: data <= 13'h0001; 
        10'b0101101001: data <= 13'h0009; 
        10'b0101101010: data <= 13'h0001; 
        10'b0101101011: data <= 13'h0006; 
        10'b0101101100: data <= 13'h0001; 
        10'b0101101101: data <= 13'h0006; 
        10'b0101101110: data <= 13'h0006; 
        10'b0101101111: data <= 13'h0006; 
        10'b0101110000: data <= 13'h000a; 
        10'b0101110001: data <= 13'h0000; 
        10'b0101110010: data <= 13'h0001; 
        10'b0101110011: data <= 13'h1ffc; 
        10'b0101110100: data <= 13'h1ffa; 
        10'b0101110101: data <= 13'h1fe8; 
        10'b0101110110: data <= 13'h1fcc; 
        10'b0101110111: data <= 13'h1fcc; 
        10'b0101111000: data <= 13'h0000; 
        10'b0101111001: data <= 13'h001c; 
        10'b0101111010: data <= 13'h0048; 
        10'b0101111011: data <= 13'h0029; 
        10'b0101111100: data <= 13'h000b; 
        10'b0101111101: data <= 13'h0005; 
        10'b0101111110: data <= 13'h1ff0; 
        10'b0101111111: data <= 13'h1fe8; 
        10'b0110000000: data <= 13'h1ff7; 
        10'b0110000001: data <= 13'h1ffd; 
        10'b0110000010: data <= 13'h1ffd; 
        10'b0110000011: data <= 13'h1fff; 
        10'b0110000100: data <= 13'h0004; 
        10'b0110000101: data <= 13'h0006; 
        10'b0110000110: data <= 13'h0009; 
        10'b0110000111: data <= 13'h0006; 
        10'b0110001000: data <= 13'h0004; 
        10'b0110001001: data <= 13'h0009; 
        10'b0110001010: data <= 13'h0005; 
        10'b0110001011: data <= 13'h0007; 
        10'b0110001100: data <= 13'h0008; 
        10'b0110001101: data <= 13'h0000; 
        10'b0110001110: data <= 13'h0001; 
        10'b0110001111: data <= 13'h1ffd; 
        10'b0110010000: data <= 13'h1ff0; 
        10'b0110010001: data <= 13'h1fe4; 
        10'b0110010010: data <= 13'h1fcd; 
        10'b0110010011: data <= 13'h1fd9; 
        10'b0110010100: data <= 13'h1fff; 
        10'b0110010101: data <= 13'h001c; 
        10'b0110010110: data <= 13'h003d; 
        10'b0110010111: data <= 13'h0027; 
        10'b0110011000: data <= 13'h000c; 
        10'b0110011001: data <= 13'h1fea; 
        10'b0110011010: data <= 13'h1fe2; 
        10'b0110011011: data <= 13'h1fe9; 
        10'b0110011100: data <= 13'h1ff3; 
        10'b0110011101: data <= 13'h1ffc; 
        10'b0110011110: data <= 13'h1ffc; 
        10'b0110011111: data <= 13'h1ffd; 
        10'b0110100000: data <= 13'h0007; 
        10'b0110100001: data <= 13'h0001; 
        10'b0110100010: data <= 13'h0002; 
        10'b0110100011: data <= 13'h0005; 
        10'b0110100100: data <= 13'h000a; 
        10'b0110100101: data <= 13'h0002; 
        10'b0110100110: data <= 13'h0006; 
        10'b0110100111: data <= 13'h0004; 
        10'b0110101000: data <= 13'h0002; 
        10'b0110101001: data <= 13'h0006; 
        10'b0110101010: data <= 13'h1ffa; 
        10'b0110101011: data <= 13'h1ffa; 
        10'b0110101100: data <= 13'h1ff6; 
        10'b0110101101: data <= 13'h1fe2; 
        10'b0110101110: data <= 13'h1fde; 
        10'b0110101111: data <= 13'h1ff7; 
        10'b0110110000: data <= 13'h000c; 
        10'b0110110001: data <= 13'h0027; 
        10'b0110110010: data <= 13'h0042; 
        10'b0110110011: data <= 13'h0017; 
        10'b0110110100: data <= 13'h0004; 
        10'b0110110101: data <= 13'h1fd7; 
        10'b0110110110: data <= 13'h1fdb; 
        10'b0110110111: data <= 13'h1fea; 
        10'b0110111000: data <= 13'h1ff3; 
        10'b0110111001: data <= 13'h1ff6; 
        10'b0110111010: data <= 13'h1ffe; 
        10'b0110111011: data <= 13'h0001; 
        10'b0110111100: data <= 13'h0003; 
        10'b0110111101: data <= 13'h0004; 
        10'b0110111110: data <= 13'h0009; 
        10'b0110111111: data <= 13'h0002; 
        10'b0111000000: data <= 13'h000a; 
        10'b0111000001: data <= 13'h0005; 
        10'b0111000010: data <= 13'h0009; 
        10'b0111000011: data <= 13'h0005; 
        10'b0111000100: data <= 13'h0003; 
        10'b0111000101: data <= 13'h1ffc; 
        10'b0111000110: data <= 13'h1ff7; 
        10'b0111000111: data <= 13'h1ff6; 
        10'b0111001000: data <= 13'h1fe9; 
        10'b0111001001: data <= 13'h1ff2; 
        10'b0111001010: data <= 13'h1ff5; 
        10'b0111001011: data <= 13'h1ffa; 
        10'b0111001100: data <= 13'h1ffe; 
        10'b0111001101: data <= 13'h0034; 
        10'b0111001110: data <= 13'h003e; 
        10'b0111001111: data <= 13'h0004; 
        10'b0111010000: data <= 13'h1fed; 
        10'b0111010001: data <= 13'h1fd3; 
        10'b0111010010: data <= 13'h1fdb; 
        10'b0111010011: data <= 13'h1fe8; 
        10'b0111010100: data <= 13'h1fee; 
        10'b0111010101: data <= 13'h1ff8; 
        10'b0111010110: data <= 13'h1ff8; 
        10'b0111010111: data <= 13'h0000; 
        10'b0111011000: data <= 13'h1ffd; 
        10'b0111011001: data <= 13'h0001; 
        10'b0111011010: data <= 13'h0002; 
        10'b0111011011: data <= 13'h0005; 
        10'b0111011100: data <= 13'h0004; 
        10'b0111011101: data <= 13'h0009; 
        10'b0111011110: data <= 13'h0002; 
        10'b0111011111: data <= 13'h0009; 
        10'b0111100000: data <= 13'h0007; 
        10'b0111100001: data <= 13'h1ffb; 
        10'b0111100010: data <= 13'h1fec; 
        10'b0111100011: data <= 13'h1feb; 
        10'b0111100100: data <= 13'h1ff1; 
        10'b0111100101: data <= 13'h1ff6; 
        10'b0111100110: data <= 13'h0007; 
        10'b0111100111: data <= 13'h0000; 
        10'b0111101000: data <= 13'h0011; 
        10'b0111101001: data <= 13'h003b; 
        10'b0111101010: data <= 13'h0033; 
        10'b0111101011: data <= 13'h1ff6; 
        10'b0111101100: data <= 13'h1fdd; 
        10'b0111101101: data <= 13'h1fd3; 
        10'b0111101110: data <= 13'h1fdb; 
        10'b0111101111: data <= 13'h1fe9; 
        10'b0111110000: data <= 13'h1ff7; 
        10'b0111110001: data <= 13'h1ffc; 
        10'b0111110010: data <= 13'h1ffd; 
        10'b0111110011: data <= 13'h1ffc; 
        10'b0111110100: data <= 13'h1ff9; 
        10'b0111110101: data <= 13'h0002; 
        10'b0111110110: data <= 13'h0006; 
        10'b0111110111: data <= 13'h0006; 
        10'b0111111000: data <= 13'h0006; 
        10'b0111111001: data <= 13'h0005; 
        10'b0111111010: data <= 13'h0003; 
        10'b0111111011: data <= 13'h0008; 
        10'b0111111100: data <= 13'h0004; 
        10'b0111111101: data <= 13'h1ff8; 
        10'b0111111110: data <= 13'h1feb; 
        10'b0111111111: data <= 13'h1feb; 
        10'b1000000000: data <= 13'h1ff8; 
        10'b1000000001: data <= 13'h0008; 
        10'b1000000010: data <= 13'h0007; 
        10'b1000000011: data <= 13'h000b; 
        10'b1000000100: data <= 13'h001b; 
        10'b1000000101: data <= 13'h002c; 
        10'b1000000110: data <= 13'h001f; 
        10'b1000000111: data <= 13'h1fec; 
        10'b1000001000: data <= 13'h1fdf; 
        10'b1000001001: data <= 13'h1fe4; 
        10'b1000001010: data <= 13'h1fe8; 
        10'b1000001011: data <= 13'h1ff0; 
        10'b1000001100: data <= 13'h1ff8; 
        10'b1000001101: data <= 13'h1ff3; 
        10'b1000001110: data <= 13'h1ffa; 
        10'b1000001111: data <= 13'h1ff7; 
        10'b1000010000: data <= 13'h1ffa; 
        10'b1000010001: data <= 13'h0005; 
        10'b1000010010: data <= 13'h0009; 
        10'b1000010011: data <= 13'h0009; 
        10'b1000010100: data <= 13'h0009; 
        10'b1000010101: data <= 13'h0007; 
        10'b1000010110: data <= 13'h0007; 
        10'b1000010111: data <= 13'h0008; 
        10'b1000011000: data <= 13'h0001; 
        10'b1000011001: data <= 13'h1ff4; 
        10'b1000011010: data <= 13'h1fe6; 
        10'b1000011011: data <= 13'h1fee; 
        10'b1000011100: data <= 13'h1ff9; 
        10'b1000011101: data <= 13'h0004; 
        10'b1000011110: data <= 13'h0002; 
        10'b1000011111: data <= 13'h0001; 
        10'b1000100000: data <= 13'h0004; 
        10'b1000100001: data <= 13'h0014; 
        10'b1000100010: data <= 13'h0004; 
        10'b1000100011: data <= 13'h1fef; 
        10'b1000100100: data <= 13'h1ff2; 
        10'b1000100101: data <= 13'h1ff4; 
        10'b1000100110: data <= 13'h1ff1; 
        10'b1000100111: data <= 13'h1ff4; 
        10'b1000101000: data <= 13'h1fef; 
        10'b1000101001: data <= 13'h1ff2; 
        10'b1000101010: data <= 13'h1ff7; 
        10'b1000101011: data <= 13'h1ff8; 
        10'b1000101100: data <= 13'h0000; 
        10'b1000101101: data <= 13'h0003; 
        10'b1000101110: data <= 13'h0003; 
        10'b1000101111: data <= 13'h0001; 
        10'b1000110000: data <= 13'h0001; 
        10'b1000110001: data <= 13'h000a; 
        10'b1000110010: data <= 13'h0005; 
        10'b1000110011: data <= 13'h0003; 
        10'b1000110100: data <= 13'h1ffd; 
        10'b1000110101: data <= 13'h1ff8; 
        10'b1000110110: data <= 13'h1ffe; 
        10'b1000110111: data <= 13'h1ffa; 
        10'b1000111000: data <= 13'h0000; 
        10'b1000111001: data <= 13'h0002; 
        10'b1000111010: data <= 13'h1ffa; 
        10'b1000111011: data <= 13'h1ffe; 
        10'b1000111100: data <= 13'h1ff6; 
        10'b1000111101: data <= 13'h1ffc; 
        10'b1000111110: data <= 13'h1ffd; 
        10'b1000111111: data <= 13'h0001; 
        10'b1001000000: data <= 13'h000a; 
        10'b1001000001: data <= 13'h0004; 
        10'b1001000010: data <= 13'h1ffc; 
        10'b1001000011: data <= 13'h1ff2; 
        10'b1001000100: data <= 13'h1fef; 
        10'b1001000101: data <= 13'h1ff0; 
        10'b1001000110: data <= 13'h1ff4; 
        10'b1001000111: data <= 13'h1ffd; 
        10'b1001001000: data <= 13'h0001; 
        10'b1001001001: data <= 13'h0008; 
        10'b1001001010: data <= 13'h0003; 
        10'b1001001011: data <= 13'h000a; 
        10'b1001001100: data <= 13'h0007; 
        10'b1001001101: data <= 13'h0004; 
        10'b1001001110: data <= 13'h0006; 
        10'b1001001111: data <= 13'h0007; 
        10'b1001010000: data <= 13'h0005; 
        10'b1001010001: data <= 13'h000f; 
        10'b1001010010: data <= 13'h000c; 
        10'b1001010011: data <= 13'h0006; 
        10'b1001010100: data <= 13'h0001; 
        10'b1001010101: data <= 13'h1ffc; 
        10'b1001010110: data <= 13'h0000; 
        10'b1001010111: data <= 13'h1ff8; 
        10'b1001011000: data <= 13'h1fed; 
        10'b1001011001: data <= 13'h1fea; 
        10'b1001011010: data <= 13'h1ffe; 
        10'b1001011011: data <= 13'h0007; 
        10'b1001011100: data <= 13'h000a; 
        10'b1001011101: data <= 13'h000c; 
        10'b1001011110: data <= 13'h0008; 
        10'b1001011111: data <= 13'h1ff2; 
        10'b1001100000: data <= 13'h1ff2; 
        10'b1001100001: data <= 13'h1ff0; 
        10'b1001100010: data <= 13'h1ff5; 
        10'b1001100011: data <= 13'h1ffa; 
        10'b1001100100: data <= 13'h0001; 
        10'b1001100101: data <= 13'h0004; 
        10'b1001100110: data <= 13'h0001; 
        10'b1001100111: data <= 13'h0001; 
        10'b1001101000: data <= 13'h0005; 
        10'b1001101001: data <= 13'h0005; 
        10'b1001101010: data <= 13'h0006; 
        10'b1001101011: data <= 13'h0001; 
        10'b1001101100: data <= 13'h000d; 
        10'b1001101101: data <= 13'h001c; 
        10'b1001101110: data <= 13'h001d; 
        10'b1001101111: data <= 13'h0012; 
        10'b1001110000: data <= 13'h0002; 
        10'b1001110001: data <= 13'h1ffe; 
        10'b1001110010: data <= 13'h1ff9; 
        10'b1001110011: data <= 13'h1fe4; 
        10'b1001110100: data <= 13'h1fd3; 
        10'b1001110101: data <= 13'h1fde; 
        10'b1001110110: data <= 13'h0000; 
        10'b1001110111: data <= 13'h0007; 
        10'b1001111000: data <= 13'h001a; 
        10'b1001111001: data <= 13'h002a; 
        10'b1001111010: data <= 13'h0013; 
        10'b1001111011: data <= 13'h0004; 
        10'b1001111100: data <= 13'h1ff6; 
        10'b1001111101: data <= 13'h1ff9; 
        10'b1001111110: data <= 13'h1fff; 
        10'b1001111111: data <= 13'h0001; 
        10'b1010000000: data <= 13'h0001; 
        10'b1010000001: data <= 13'h0004; 
        10'b1010000010: data <= 13'h0009; 
        10'b1010000011: data <= 13'h0005; 
        10'b1010000100: data <= 13'h0009; 
        10'b1010000101: data <= 13'h0005; 
        10'b1010000110: data <= 13'h0007; 
        10'b1010000111: data <= 13'h0004; 
        10'b1010001000: data <= 13'h000b; 
        10'b1010001001: data <= 13'h0018; 
        10'b1010001010: data <= 13'h001a; 
        10'b1010001011: data <= 13'h000c; 
        10'b1010001100: data <= 13'h0003; 
        10'b1010001101: data <= 13'h1ffa; 
        10'b1010001110: data <= 13'h1ffc; 
        10'b1010001111: data <= 13'h1ff0; 
        10'b1010010000: data <= 13'h1ff5; 
        10'b1010010001: data <= 13'h1ff6; 
        10'b1010010010: data <= 13'h1ff3; 
        10'b1010010011: data <= 13'h0005; 
        10'b1010010100: data <= 13'h001e; 
        10'b1010010101: data <= 13'h0024; 
        10'b1010010110: data <= 13'h0010; 
        10'b1010010111: data <= 13'h1ffd; 
        10'b1010011000: data <= 13'h1ff9; 
        10'b1010011001: data <= 13'h1ff5; 
        10'b1010011010: data <= 13'h1ffc; 
        10'b1010011011: data <= 13'h1ffd; 
        10'b1010011100: data <= 13'h0002; 
        10'b1010011101: data <= 13'h0001; 
        10'b1010011110: data <= 13'h0002; 
        10'b1010011111: data <= 13'h0001; 
        10'b1010100000: data <= 13'h0002; 
        10'b1010100001: data <= 13'h0001; 
        10'b1010100010: data <= 13'h0004; 
        10'b1010100011: data <= 13'h0001; 
        10'b1010100100: data <= 13'h0005; 
        10'b1010100101: data <= 13'h000b; 
        10'b1010100110: data <= 13'h000b; 
        10'b1010100111: data <= 13'h1ffc; 
        10'b1010101000: data <= 13'h1ff0; 
        10'b1010101001: data <= 13'h1ff0; 
        10'b1010101010: data <= 13'h1fe4; 
        10'b1010101011: data <= 13'h1fe5; 
        10'b1010101100: data <= 13'h1fe8; 
        10'b1010101101: data <= 13'h1feb; 
        10'b1010101110: data <= 13'h1feb; 
        10'b1010101111: data <= 13'h1feb; 
        10'b1010110000: data <= 13'h1ffa; 
        10'b1010110001: data <= 13'h0003; 
        10'b1010110010: data <= 13'h0005; 
        10'b1010110011: data <= 13'h0007; 
        10'b1010110100: data <= 13'h0006; 
        10'b1010110101: data <= 13'h0001; 
        10'b1010110110: data <= 13'h0003; 
        10'b1010110111: data <= 13'h0008; 
        10'b1010111000: data <= 13'h0002; 
        10'b1010111001: data <= 13'h0004; 
        10'b1010111010: data <= 13'h0007; 
        10'b1010111011: data <= 13'h0002; 
        10'b1010111100: data <= 13'h0009; 
        10'b1010111101: data <= 13'h0003; 
        10'b1010111110: data <= 13'h0004; 
        10'b1010111111: data <= 13'h0005; 
        10'b1011000000: data <= 13'h0007; 
        10'b1011000001: data <= 13'h0007; 
        10'b1011000010: data <= 13'h0000; 
        10'b1011000011: data <= 13'h1ffc; 
        10'b1011000100: data <= 13'h1ffe; 
        10'b1011000101: data <= 13'h1ffc; 
        10'b1011000110: data <= 13'h1ff0; 
        10'b1011000111: data <= 13'h1fed; 
        10'b1011001000: data <= 13'h1ff2; 
        10'b1011001001: data <= 13'h1fec; 
        10'b1011001010: data <= 13'h1ff4; 
        10'b1011001011: data <= 13'h1ff1; 
        10'b1011001100: data <= 13'h1ff7; 
        10'b1011001101: data <= 13'h1ffe; 
        10'b1011001110: data <= 13'h0003; 
        10'b1011001111: data <= 13'h0006; 
        10'b1011010000: data <= 13'h0001; 
        10'b1011010001: data <= 13'h0006; 
        10'b1011010010: data <= 13'h0003; 
        10'b1011010011: data <= 13'h0008; 
        10'b1011010100: data <= 13'h0002; 
        10'b1011010101: data <= 13'h0002; 
        10'b1011010110: data <= 13'h0004; 
        10'b1011010111: data <= 13'h0003; 
        10'b1011011000: data <= 13'h0003; 
        10'b1011011001: data <= 13'h0007; 
        10'b1011011010: data <= 13'h0006; 
        10'b1011011011: data <= 13'h0002; 
        10'b1011011100: data <= 13'h0006; 
        10'b1011011101: data <= 13'h0009; 
        10'b1011011110: data <= 13'h0006; 
        10'b1011011111: data <= 13'h0005; 
        10'b1011100000: data <= 13'h0008; 
        10'b1011100001: data <= 13'h0006; 
        10'b1011100010: data <= 13'h0001; 
        10'b1011100011: data <= 13'h0005; 
        10'b1011100100: data <= 13'h0005; 
        10'b1011100101: data <= 13'h0003; 
        10'b1011100110: data <= 13'h0000; 
        10'b1011100111: data <= 13'h0003; 
        10'b1011101000: data <= 13'h0006; 
        10'b1011101001: data <= 13'h0009; 
        10'b1011101010: data <= 13'h0006; 
        10'b1011101011: data <= 13'h0001; 
        10'b1011101100: data <= 13'h0006; 
        10'b1011101101: data <= 13'h0006; 
        10'b1011101110: data <= 13'h0005; 
        10'b1011101111: data <= 13'h0003; 
        10'b1011110000: data <= 13'h0002; 
        10'b1011110001: data <= 13'h0006; 
        10'b1011110010: data <= 13'h0009; 
        10'b1011110011: data <= 13'h0007; 
        10'b1011110100: data <= 13'h0007; 
        10'b1011110101: data <= 13'h0009; 
        10'b1011110110: data <= 13'h0001; 
        10'b1011110111: data <= 13'h0005; 
        10'b1011111000: data <= 13'h000a; 
        10'b1011111001: data <= 13'h0008; 
        10'b1011111010: data <= 13'h0009; 
        10'b1011111011: data <= 13'h0008; 
        10'b1011111100: data <= 13'h0009; 
        10'b1011111101: data <= 13'h0004; 
        10'b1011111110: data <= 13'h0008; 
        10'b1011111111: data <= 13'h0008; 
        10'b1100000000: data <= 13'h0001; 
        10'b1100000001: data <= 13'h0002; 
        10'b1100000010: data <= 13'h0009; 
        10'b1100000011: data <= 13'h0006; 
        10'b1100000100: data <= 13'h0006; 
        10'b1100000101: data <= 13'h0001; 
        10'b1100000110: data <= 13'h0004; 
        10'b1100000111: data <= 13'h0002; 
        10'b1100001000: data <= 13'h0002; 
        10'b1100001001: data <= 13'h0003; 
        10'b1100001010: data <= 13'h0006; 
        10'b1100001011: data <= 13'h0008; 
        10'b1100001100: data <= 13'h0009; 
        10'b1100001101: data <= 13'h0009; 
        10'b1100001110: data <= 13'h0009; 
        10'b1100001111: data <= 13'h0003; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 8) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 14'h0010; 
        10'b0000000001: data <= 14'h0008; 
        10'b0000000010: data <= 14'h0008; 
        10'b0000000011: data <= 14'h0003; 
        10'b0000000100: data <= 14'h000e; 
        10'b0000000101: data <= 14'h000d; 
        10'b0000000110: data <= 14'h000f; 
        10'b0000000111: data <= 14'h0004; 
        10'b0000001000: data <= 14'h000d; 
        10'b0000001001: data <= 14'h0004; 
        10'b0000001010: data <= 14'h000c; 
        10'b0000001011: data <= 14'h000a; 
        10'b0000001100: data <= 14'h000e; 
        10'b0000001101: data <= 14'h0012; 
        10'b0000001110: data <= 14'h0010; 
        10'b0000001111: data <= 14'h000b; 
        10'b0000010000: data <= 14'h000b; 
        10'b0000010001: data <= 14'h0004; 
        10'b0000010010: data <= 14'h0013; 
        10'b0000010011: data <= 14'h0012; 
        10'b0000010100: data <= 14'h000b; 
        10'b0000010101: data <= 14'h000e; 
        10'b0000010110: data <= 14'h000a; 
        10'b0000010111: data <= 14'h0010; 
        10'b0000011000: data <= 14'h0006; 
        10'b0000011001: data <= 14'h0011; 
        10'b0000011010: data <= 14'h000a; 
        10'b0000011011: data <= 14'h000f; 
        10'b0000011100: data <= 14'h0002; 
        10'b0000011101: data <= 14'h0010; 
        10'b0000011110: data <= 14'h0005; 
        10'b0000011111: data <= 14'h000b; 
        10'b0000100000: data <= 14'h000a; 
        10'b0000100001: data <= 14'h0004; 
        10'b0000100010: data <= 14'h0006; 
        10'b0000100011: data <= 14'h000f; 
        10'b0000100100: data <= 14'h000e; 
        10'b0000100101: data <= 14'h000c; 
        10'b0000100110: data <= 14'h000c; 
        10'b0000100111: data <= 14'h0009; 
        10'b0000101000: data <= 14'h000e; 
        10'b0000101001: data <= 14'h0010; 
        10'b0000101010: data <= 14'h0014; 
        10'b0000101011: data <= 14'h000a; 
        10'b0000101100: data <= 14'h0008; 
        10'b0000101101: data <= 14'h0010; 
        10'b0000101110: data <= 14'h000b; 
        10'b0000101111: data <= 14'h0007; 
        10'b0000110000: data <= 14'h0012; 
        10'b0000110001: data <= 14'h0011; 
        10'b0000110010: data <= 14'h0007; 
        10'b0000110011: data <= 14'h0012; 
        10'b0000110100: data <= 14'h0013; 
        10'b0000110101: data <= 14'h000a; 
        10'b0000110110: data <= 14'h0011; 
        10'b0000110111: data <= 14'h000d; 
        10'b0000111000: data <= 14'h0010; 
        10'b0000111001: data <= 14'h000c; 
        10'b0000111010: data <= 14'h0014; 
        10'b0000111011: data <= 14'h0004; 
        10'b0000111100: data <= 14'h0004; 
        10'b0000111101: data <= 14'h000d; 
        10'b0000111110: data <= 14'h000a; 
        10'b0000111111: data <= 14'h0009; 
        10'b0001000000: data <= 14'h0006; 
        10'b0001000001: data <= 14'h000b; 
        10'b0001000010: data <= 14'h0000; 
        10'b0001000011: data <= 14'h0005; 
        10'b0001000100: data <= 14'h0001; 
        10'b0001000101: data <= 14'h0005; 
        10'b0001000110: data <= 14'h000a; 
        10'b0001000111: data <= 14'h0010; 
        10'b0001001000: data <= 14'h000c; 
        10'b0001001001: data <= 14'h0000; 
        10'b0001001010: data <= 14'h000c; 
        10'b0001001011: data <= 14'h0007; 
        10'b0001001100: data <= 14'h0010; 
        10'b0001001101: data <= 14'h0007; 
        10'b0001001110: data <= 14'h0011; 
        10'b0001001111: data <= 14'h000d; 
        10'b0001010000: data <= 14'h000e; 
        10'b0001010001: data <= 14'h0002; 
        10'b0001010010: data <= 14'h000f; 
        10'b0001010011: data <= 14'h000f; 
        10'b0001010100: data <= 14'h0006; 
        10'b0001010101: data <= 14'h0007; 
        10'b0001010110: data <= 14'h000b; 
        10'b0001010111: data <= 14'h0009; 
        10'b0001011000: data <= 14'h0012; 
        10'b0001011001: data <= 14'h000a; 
        10'b0001011010: data <= 14'h0002; 
        10'b0001011011: data <= 14'h0012; 
        10'b0001011100: data <= 14'h3ffe; 
        10'b0001011101: data <= 14'h3ffc; 
        10'b0001011110: data <= 14'h3ffd; 
        10'b0001011111: data <= 14'h3ff6; 
        10'b0001100000: data <= 14'h3ffc; 
        10'b0001100001: data <= 14'h0001; 
        10'b0001100010: data <= 14'h0007; 
        10'b0001100011: data <= 14'h000f; 
        10'b0001100100: data <= 14'h3ff9; 
        10'b0001100101: data <= 14'h3ffd; 
        10'b0001100110: data <= 14'h0000; 
        10'b0001100111: data <= 14'h3ff4; 
        10'b0001101000: data <= 14'h3fff; 
        10'b0001101001: data <= 14'h0005; 
        10'b0001101010: data <= 14'h000c; 
        10'b0001101011: data <= 14'h000c; 
        10'b0001101100: data <= 14'h3ffe; 
        10'b0001101101: data <= 14'h0011; 
        10'b0001101110: data <= 14'h0006; 
        10'b0001101111: data <= 14'h0012; 
        10'b0001110000: data <= 14'h000d; 
        10'b0001110001: data <= 14'h0008; 
        10'b0001110010: data <= 14'h0013; 
        10'b0001110011: data <= 14'h0012; 
        10'b0001110100: data <= 14'h0002; 
        10'b0001110101: data <= 14'h0004; 
        10'b0001110110: data <= 14'h0010; 
        10'b0001110111: data <= 14'h000a; 
        10'b0001111000: data <= 14'h0004; 
        10'b0001111001: data <= 14'h3fef; 
        10'b0001111010: data <= 14'h0002; 
        10'b0001111011: data <= 14'h0006; 
        10'b0001111100: data <= 14'h0009; 
        10'b0001111101: data <= 14'h0011; 
        10'b0001111110: data <= 14'h0013; 
        10'b0001111111: data <= 14'h0028; 
        10'b0010000000: data <= 14'h000b; 
        10'b0010000001: data <= 14'h3ff8; 
        10'b0010000010: data <= 14'h3ff7; 
        10'b0010000011: data <= 14'h0006; 
        10'b0010000100: data <= 14'h0016; 
        10'b0010000101: data <= 14'h0019; 
        10'b0010000110: data <= 14'h0018; 
        10'b0010000111: data <= 14'h001d; 
        10'b0010001000: data <= 14'h000f; 
        10'b0010001001: data <= 14'h0007; 
        10'b0010001010: data <= 14'h0006; 
        10'b0010001011: data <= 14'h0007; 
        10'b0010001100: data <= 14'h0002; 
        10'b0010001101: data <= 14'h0010; 
        10'b0010001110: data <= 14'h0003; 
        10'b0010001111: data <= 14'h000b; 
        10'b0010010000: data <= 14'h0003; 
        10'b0010010001: data <= 14'h000b; 
        10'b0010010010: data <= 14'h0003; 
        10'b0010010011: data <= 14'h3ffc; 
        10'b0010010100: data <= 14'h3fdc; 
        10'b0010010101: data <= 14'h3fdc; 
        10'b0010010110: data <= 14'h3ff0; 
        10'b0010010111: data <= 14'h0000; 
        10'b0010011000: data <= 14'h000d; 
        10'b0010011001: data <= 14'h000f; 
        10'b0010011010: data <= 14'h001a; 
        10'b0010011011: data <= 14'h0015; 
        10'b0010011100: data <= 14'h000c; 
        10'b0010011101: data <= 14'h3fec; 
        10'b0010011110: data <= 14'h3ffe; 
        10'b0010011111: data <= 14'h0004; 
        10'b0010100000: data <= 14'h0014; 
        10'b0010100001: data <= 14'h001f; 
        10'b0010100010: data <= 14'h0034; 
        10'b0010100011: data <= 14'h0021; 
        10'b0010100100: data <= 14'h001b; 
        10'b0010100101: data <= 14'h3ff9; 
        10'b0010100110: data <= 14'h0007; 
        10'b0010100111: data <= 14'h0004; 
        10'b0010101000: data <= 14'h0003; 
        10'b0010101001: data <= 14'h000c; 
        10'b0010101010: data <= 14'h0002; 
        10'b0010101011: data <= 14'h0009; 
        10'b0010101100: data <= 14'h0002; 
        10'b0010101101: data <= 14'h3ffb; 
        10'b0010101110: data <= 14'h3fec; 
        10'b0010101111: data <= 14'h3fed; 
        10'b0010110000: data <= 14'h3fd3; 
        10'b0010110001: data <= 14'h3fca; 
        10'b0010110010: data <= 14'h3fde; 
        10'b0010110011: data <= 14'h3ff8; 
        10'b0010110100: data <= 14'h3ff8; 
        10'b0010110101: data <= 14'h3fef; 
        10'b0010110110: data <= 14'h3ff8; 
        10'b0010110111: data <= 14'h3fd9; 
        10'b0010111000: data <= 14'h3fd6; 
        10'b0010111001: data <= 14'h3fd6; 
        10'b0010111010: data <= 14'h3fee; 
        10'b0010111011: data <= 14'h3ff3; 
        10'b0010111100: data <= 14'h0014; 
        10'b0010111101: data <= 14'h0020; 
        10'b0010111110: data <= 14'h001e; 
        10'b0010111111: data <= 14'h0019; 
        10'b0011000000: data <= 14'h0007; 
        10'b0011000001: data <= 14'h3ffb; 
        10'b0011000010: data <= 14'h0000; 
        10'b0011000011: data <= 14'h0009; 
        10'b0011000100: data <= 14'h0008; 
        10'b0011000101: data <= 14'h0004; 
        10'b0011000110: data <= 14'h0005; 
        10'b0011000111: data <= 14'h0001; 
        10'b0011001000: data <= 14'h000d; 
        10'b0011001001: data <= 14'h3ffd; 
        10'b0011001010: data <= 14'h3fed; 
        10'b0011001011: data <= 14'h3fda; 
        10'b0011001100: data <= 14'h3fc4; 
        10'b0011001101: data <= 14'h3fb3; 
        10'b0011001110: data <= 14'h3fcc; 
        10'b0011001111: data <= 14'h3fe9; 
        10'b0011010000: data <= 14'h3feb; 
        10'b0011010001: data <= 14'h3fe2; 
        10'b0011010010: data <= 14'h3fdb; 
        10'b0011010011: data <= 14'h3fc6; 
        10'b0011010100: data <= 14'h3fce; 
        10'b0011010101: data <= 14'h3fd1; 
        10'b0011010110: data <= 14'h3fd6; 
        10'b0011010111: data <= 14'h3fff; 
        10'b0011011000: data <= 14'h0009; 
        10'b0011011001: data <= 14'h0006; 
        10'b0011011010: data <= 14'h0005; 
        10'b0011011011: data <= 14'h3ff0; 
        10'b0011011100: data <= 14'h3fea; 
        10'b0011011101: data <= 14'h3ff7; 
        10'b0011011110: data <= 14'h0007; 
        10'b0011011111: data <= 14'h0008; 
        10'b0011100000: data <= 14'h0009; 
        10'b0011100001: data <= 14'h0008; 
        10'b0011100010: data <= 14'h0008; 
        10'b0011100011: data <= 14'h0010; 
        10'b0011100100: data <= 14'h0005; 
        10'b0011100101: data <= 14'h3fff; 
        10'b0011100110: data <= 14'h3fea; 
        10'b0011100111: data <= 14'h3fde; 
        10'b0011101000: data <= 14'h3fba; 
        10'b0011101001: data <= 14'h3fb4; 
        10'b0011101010: data <= 14'h3fb8; 
        10'b0011101011: data <= 14'h3fd9; 
        10'b0011101100: data <= 14'h3fee; 
        10'b0011101101: data <= 14'h3fea; 
        10'b0011101110: data <= 14'h3fee; 
        10'b0011101111: data <= 14'h0008; 
        10'b0011110000: data <= 14'h3fe0; 
        10'b0011110001: data <= 14'h3ff5; 
        10'b0011110010: data <= 14'h3ffe; 
        10'b0011110011: data <= 14'h0004; 
        10'b0011110100: data <= 14'h3fe8; 
        10'b0011110101: data <= 14'h3fe9; 
        10'b0011110110: data <= 14'h3fdb; 
        10'b0011110111: data <= 14'h3fcf; 
        10'b0011111000: data <= 14'h3fd9; 
        10'b0011111001: data <= 14'h3ff6; 
        10'b0011111010: data <= 14'h000e; 
        10'b0011111011: data <= 14'h0013; 
        10'b0011111100: data <= 14'h0013; 
        10'b0011111101: data <= 14'h0004; 
        10'b0011111110: data <= 14'h0008; 
        10'b0011111111: data <= 14'h0007; 
        10'b0100000000: data <= 14'h3fff; 
        10'b0100000001: data <= 14'h3ffe; 
        10'b0100000010: data <= 14'h3fe4; 
        10'b0100000011: data <= 14'h3fe5; 
        10'b0100000100: data <= 14'h3fd0; 
        10'b0100000101: data <= 14'h3fb6; 
        10'b0100000110: data <= 14'h3fbd; 
        10'b0100000111: data <= 14'h3fe5; 
        10'b0100001000: data <= 14'h3fec; 
        10'b0100001001: data <= 14'h000f; 
        10'b0100001010: data <= 14'h0030; 
        10'b0100001011: data <= 14'h0044; 
        10'b0100001100: data <= 14'h0019; 
        10'b0100001101: data <= 14'h3ffe; 
        10'b0100001110: data <= 14'h3ff5; 
        10'b0100001111: data <= 14'h3fd2; 
        10'b0100010000: data <= 14'h3fc7; 
        10'b0100010001: data <= 14'h3fc8; 
        10'b0100010010: data <= 14'h3fb9; 
        10'b0100010011: data <= 14'h3fc3; 
        10'b0100010100: data <= 14'h3fdf; 
        10'b0100010101: data <= 14'h0004; 
        10'b0100010110: data <= 14'h0010; 
        10'b0100010111: data <= 14'h000b; 
        10'b0100011000: data <= 14'h0011; 
        10'b0100011001: data <= 14'h0013; 
        10'b0100011010: data <= 14'h0010; 
        10'b0100011011: data <= 14'h0002; 
        10'b0100011100: data <= 14'h000d; 
        10'b0100011101: data <= 14'h3ff1; 
        10'b0100011110: data <= 14'h3fe5; 
        10'b0100011111: data <= 14'h3ff4; 
        10'b0100100000: data <= 14'h3fdb; 
        10'b0100100001: data <= 14'h3fda; 
        10'b0100100010: data <= 14'h3fe4; 
        10'b0100100011: data <= 14'h3fed; 
        10'b0100100100: data <= 14'h3ff4; 
        10'b0100100101: data <= 14'h0026; 
        10'b0100100110: data <= 14'h007b; 
        10'b0100100111: data <= 14'h0082; 
        10'b0100101000: data <= 14'h003e; 
        10'b0100101001: data <= 14'h3fff; 
        10'b0100101010: data <= 14'h3fdb; 
        10'b0100101011: data <= 14'h3fd4; 
        10'b0100101100: data <= 14'h3fca; 
        10'b0100101101: data <= 14'h3fcf; 
        10'b0100101110: data <= 14'h3fd2; 
        10'b0100101111: data <= 14'h3fe4; 
        10'b0100110000: data <= 14'h3ff6; 
        10'b0100110001: data <= 14'h3ffe; 
        10'b0100110010: data <= 14'h0010; 
        10'b0100110011: data <= 14'h0007; 
        10'b0100110100: data <= 14'h0003; 
        10'b0100110101: data <= 14'h0003; 
        10'b0100110110: data <= 14'h000d; 
        10'b0100110111: data <= 14'h000e; 
        10'b0100111000: data <= 14'h0000; 
        10'b0100111001: data <= 14'h3ffc; 
        10'b0100111010: data <= 14'h3ffe; 
        10'b0100111011: data <= 14'h3fe9; 
        10'b0100111100: data <= 14'h3ff1; 
        10'b0100111101: data <= 14'h3fe9; 
        10'b0100111110: data <= 14'h3fde; 
        10'b0100111111: data <= 14'h3fcc; 
        10'b0101000000: data <= 14'h3ffa; 
        10'b0101000001: data <= 14'h0041; 
        10'b0101000010: data <= 14'h0094; 
        10'b0101000011: data <= 14'h009d; 
        10'b0101000100: data <= 14'h003a; 
        10'b0101000101: data <= 14'h3ff3; 
        10'b0101000110: data <= 14'h3ff4; 
        10'b0101000111: data <= 14'h3fe1; 
        10'b0101001000: data <= 14'h3fdf; 
        10'b0101001001: data <= 14'h3fe2; 
        10'b0101001010: data <= 14'h3fe4; 
        10'b0101001011: data <= 14'h3ff3; 
        10'b0101001100: data <= 14'h3ffa; 
        10'b0101001101: data <= 14'h000d; 
        10'b0101001110: data <= 14'h0012; 
        10'b0101001111: data <= 14'h000d; 
        10'b0101010000: data <= 14'h0002; 
        10'b0101010001: data <= 14'h0012; 
        10'b0101010010: data <= 14'h0008; 
        10'b0101010011: data <= 14'h0006; 
        10'b0101010100: data <= 14'h0012; 
        10'b0101010101: data <= 14'h3ffd; 
        10'b0101010110: data <= 14'h3ffb; 
        10'b0101010111: data <= 14'h3ff8; 
        10'b0101011000: data <= 14'h3fea; 
        10'b0101011001: data <= 14'h3fe3; 
        10'b0101011010: data <= 14'h3fc2; 
        10'b0101011011: data <= 14'h3fa9; 
        10'b0101011100: data <= 14'h3ffd; 
        10'b0101011101: data <= 14'h0042; 
        10'b0101011110: data <= 14'h00af; 
        10'b0101011111: data <= 14'h0079; 
        10'b0101100000: data <= 14'h0018; 
        10'b0101100001: data <= 14'h000d; 
        10'b0101100010: data <= 14'h3ff9; 
        10'b0101100011: data <= 14'h3fdd; 
        10'b0101100100: data <= 14'h3fea; 
        10'b0101100101: data <= 14'h3ff5; 
        10'b0101100110: data <= 14'h3ffa; 
        10'b0101100111: data <= 14'h3ff8; 
        10'b0101101000: data <= 14'h0001; 
        10'b0101101001: data <= 14'h0012; 
        10'b0101101010: data <= 14'h0003; 
        10'b0101101011: data <= 14'h000d; 
        10'b0101101100: data <= 14'h0002; 
        10'b0101101101: data <= 14'h000c; 
        10'b0101101110: data <= 14'h000b; 
        10'b0101101111: data <= 14'h000c; 
        10'b0101110000: data <= 14'h0014; 
        10'b0101110001: data <= 14'h0000; 
        10'b0101110010: data <= 14'h0002; 
        10'b0101110011: data <= 14'h3ff7; 
        10'b0101110100: data <= 14'h3ff4; 
        10'b0101110101: data <= 14'h3fcf; 
        10'b0101110110: data <= 14'h3f99; 
        10'b0101110111: data <= 14'h3f97; 
        10'b0101111000: data <= 14'h0000; 
        10'b0101111001: data <= 14'h0037; 
        10'b0101111010: data <= 14'h0090; 
        10'b0101111011: data <= 14'h0051; 
        10'b0101111100: data <= 14'h0015; 
        10'b0101111101: data <= 14'h000a; 
        10'b0101111110: data <= 14'h3fdf; 
        10'b0101111111: data <= 14'h3fd0; 
        10'b0110000000: data <= 14'h3fef; 
        10'b0110000001: data <= 14'h3ffa; 
        10'b0110000010: data <= 14'h3ffa; 
        10'b0110000011: data <= 14'h3ffe; 
        10'b0110000100: data <= 14'h0008; 
        10'b0110000101: data <= 14'h000c; 
        10'b0110000110: data <= 14'h0011; 
        10'b0110000111: data <= 14'h000b; 
        10'b0110001000: data <= 14'h0009; 
        10'b0110001001: data <= 14'h0013; 
        10'b0110001010: data <= 14'h000b; 
        10'b0110001011: data <= 14'h000f; 
        10'b0110001100: data <= 14'h000f; 
        10'b0110001101: data <= 14'h0000; 
        10'b0110001110: data <= 14'h0003; 
        10'b0110001111: data <= 14'h3ffa; 
        10'b0110010000: data <= 14'h3fe0; 
        10'b0110010001: data <= 14'h3fc9; 
        10'b0110010010: data <= 14'h3f99; 
        10'b0110010011: data <= 14'h3fb2; 
        10'b0110010100: data <= 14'h3ffe; 
        10'b0110010101: data <= 14'h0038; 
        10'b0110010110: data <= 14'h007b; 
        10'b0110010111: data <= 14'h004f; 
        10'b0110011000: data <= 14'h0018; 
        10'b0110011001: data <= 14'h3fd4; 
        10'b0110011010: data <= 14'h3fc5; 
        10'b0110011011: data <= 14'h3fd3; 
        10'b0110011100: data <= 14'h3fe5; 
        10'b0110011101: data <= 14'h3ff8; 
        10'b0110011110: data <= 14'h3ff8; 
        10'b0110011111: data <= 14'h3ffa; 
        10'b0110100000: data <= 14'h000d; 
        10'b0110100001: data <= 14'h0002; 
        10'b0110100010: data <= 14'h0004; 
        10'b0110100011: data <= 14'h000b; 
        10'b0110100100: data <= 14'h0014; 
        10'b0110100101: data <= 14'h0003; 
        10'b0110100110: data <= 14'h000d; 
        10'b0110100111: data <= 14'h0008; 
        10'b0110101000: data <= 14'h0005; 
        10'b0110101001: data <= 14'h000c; 
        10'b0110101010: data <= 14'h3ff5; 
        10'b0110101011: data <= 14'h3ff3; 
        10'b0110101100: data <= 14'h3fec; 
        10'b0110101101: data <= 14'h3fc3; 
        10'b0110101110: data <= 14'h3fbc; 
        10'b0110101111: data <= 14'h3fef; 
        10'b0110110000: data <= 14'h0019; 
        10'b0110110001: data <= 14'h004f; 
        10'b0110110010: data <= 14'h0083; 
        10'b0110110011: data <= 14'h002e; 
        10'b0110110100: data <= 14'h0008; 
        10'b0110110101: data <= 14'h3fad; 
        10'b0110110110: data <= 14'h3fb7; 
        10'b0110110111: data <= 14'h3fd3; 
        10'b0110111000: data <= 14'h3fe5; 
        10'b0110111001: data <= 14'h3fed; 
        10'b0110111010: data <= 14'h3ffb; 
        10'b0110111011: data <= 14'h0001; 
        10'b0110111100: data <= 14'h0007; 
        10'b0110111101: data <= 14'h0009; 
        10'b0110111110: data <= 14'h0012; 
        10'b0110111111: data <= 14'h0003; 
        10'b0111000000: data <= 14'h0013; 
        10'b0111000001: data <= 14'h0009; 
        10'b0111000010: data <= 14'h0012; 
        10'b0111000011: data <= 14'h000b; 
        10'b0111000100: data <= 14'h0006; 
        10'b0111000101: data <= 14'h3ff8; 
        10'b0111000110: data <= 14'h3fee; 
        10'b0111000111: data <= 14'h3fed; 
        10'b0111001000: data <= 14'h3fd1; 
        10'b0111001001: data <= 14'h3fe4; 
        10'b0111001010: data <= 14'h3fea; 
        10'b0111001011: data <= 14'h3ff4; 
        10'b0111001100: data <= 14'h3ffd; 
        10'b0111001101: data <= 14'h0067; 
        10'b0111001110: data <= 14'h007c; 
        10'b0111001111: data <= 14'h0007; 
        10'b0111010000: data <= 14'h3fda; 
        10'b0111010001: data <= 14'h3fa7; 
        10'b0111010010: data <= 14'h3fb6; 
        10'b0111010011: data <= 14'h3fd0; 
        10'b0111010100: data <= 14'h3fdc; 
        10'b0111010101: data <= 14'h3ff1; 
        10'b0111010110: data <= 14'h3ff0; 
        10'b0111010111: data <= 14'h0000; 
        10'b0111011000: data <= 14'h3ff9; 
        10'b0111011001: data <= 14'h0001; 
        10'b0111011010: data <= 14'h0005; 
        10'b0111011011: data <= 14'h000a; 
        10'b0111011100: data <= 14'h0008; 
        10'b0111011101: data <= 14'h0013; 
        10'b0111011110: data <= 14'h0004; 
        10'b0111011111: data <= 14'h0013; 
        10'b0111100000: data <= 14'h000e; 
        10'b0111100001: data <= 14'h3ff5; 
        10'b0111100010: data <= 14'h3fd9; 
        10'b0111100011: data <= 14'h3fd5; 
        10'b0111100100: data <= 14'h3fe2; 
        10'b0111100101: data <= 14'h3fed; 
        10'b0111100110: data <= 14'h000e; 
        10'b0111100111: data <= 14'h0000; 
        10'b0111101000: data <= 14'h0022; 
        10'b0111101001: data <= 14'h0076; 
        10'b0111101010: data <= 14'h0065; 
        10'b0111101011: data <= 14'h3feb; 
        10'b0111101100: data <= 14'h3fba; 
        10'b0111101101: data <= 14'h3fa6; 
        10'b0111101110: data <= 14'h3fb7; 
        10'b0111101111: data <= 14'h3fd2; 
        10'b0111110000: data <= 14'h3fef; 
        10'b0111110001: data <= 14'h3ff7; 
        10'b0111110010: data <= 14'h3ffa; 
        10'b0111110011: data <= 14'h3ff8; 
        10'b0111110100: data <= 14'h3ff2; 
        10'b0111110101: data <= 14'h0004; 
        10'b0111110110: data <= 14'h000b; 
        10'b0111110111: data <= 14'h000d; 
        10'b0111111000: data <= 14'h000c; 
        10'b0111111001: data <= 14'h000b; 
        10'b0111111010: data <= 14'h0007; 
        10'b0111111011: data <= 14'h0010; 
        10'b0111111100: data <= 14'h0009; 
        10'b0111111101: data <= 14'h3ff1; 
        10'b0111111110: data <= 14'h3fd6; 
        10'b0111111111: data <= 14'h3fd6; 
        10'b1000000000: data <= 14'h3ff0; 
        10'b1000000001: data <= 14'h0010; 
        10'b1000000010: data <= 14'h000d; 
        10'b1000000011: data <= 14'h0015; 
        10'b1000000100: data <= 14'h0037; 
        10'b1000000101: data <= 14'h0058; 
        10'b1000000110: data <= 14'h003d; 
        10'b1000000111: data <= 14'h3fd8; 
        10'b1000001000: data <= 14'h3fbe; 
        10'b1000001001: data <= 14'h3fc7; 
        10'b1000001010: data <= 14'h3fd0; 
        10'b1000001011: data <= 14'h3fe0; 
        10'b1000001100: data <= 14'h3ff0; 
        10'b1000001101: data <= 14'h3fe5; 
        10'b1000001110: data <= 14'h3ff4; 
        10'b1000001111: data <= 14'h3fee; 
        10'b1000010000: data <= 14'h3ff5; 
        10'b1000010001: data <= 14'h000a; 
        10'b1000010010: data <= 14'h0012; 
        10'b1000010011: data <= 14'h0012; 
        10'b1000010100: data <= 14'h0012; 
        10'b1000010101: data <= 14'h000d; 
        10'b1000010110: data <= 14'h000e; 
        10'b1000010111: data <= 14'h000f; 
        10'b1000011000: data <= 14'h0002; 
        10'b1000011001: data <= 14'h3fe9; 
        10'b1000011010: data <= 14'h3fcc; 
        10'b1000011011: data <= 14'h3fdd; 
        10'b1000011100: data <= 14'h3ff2; 
        10'b1000011101: data <= 14'h0008; 
        10'b1000011110: data <= 14'h0004; 
        10'b1000011111: data <= 14'h0003; 
        10'b1000100000: data <= 14'h0007; 
        10'b1000100001: data <= 14'h0029; 
        10'b1000100010: data <= 14'h0009; 
        10'b1000100011: data <= 14'h3fdf; 
        10'b1000100100: data <= 14'h3fe4; 
        10'b1000100101: data <= 14'h3fe8; 
        10'b1000100110: data <= 14'h3fe2; 
        10'b1000100111: data <= 14'h3fe9; 
        10'b1000101000: data <= 14'h3fde; 
        10'b1000101001: data <= 14'h3fe3; 
        10'b1000101010: data <= 14'h3fef; 
        10'b1000101011: data <= 14'h3ff1; 
        10'b1000101100: data <= 14'h0001; 
        10'b1000101101: data <= 14'h0006; 
        10'b1000101110: data <= 14'h0006; 
        10'b1000101111: data <= 14'h0003; 
        10'b1000110000: data <= 14'h0003; 
        10'b1000110001: data <= 14'h0013; 
        10'b1000110010: data <= 14'h000a; 
        10'b1000110011: data <= 14'h0007; 
        10'b1000110100: data <= 14'h3ffb; 
        10'b1000110101: data <= 14'h3fef; 
        10'b1000110110: data <= 14'h3ffd; 
        10'b1000110111: data <= 14'h3ff5; 
        10'b1000111000: data <= 14'h0000; 
        10'b1000111001: data <= 14'h0005; 
        10'b1000111010: data <= 14'h3ff3; 
        10'b1000111011: data <= 14'h3ffb; 
        10'b1000111100: data <= 14'h3feb; 
        10'b1000111101: data <= 14'h3ff9; 
        10'b1000111110: data <= 14'h3ffb; 
        10'b1000111111: data <= 14'h0001; 
        10'b1001000000: data <= 14'h0014; 
        10'b1001000001: data <= 14'h0007; 
        10'b1001000010: data <= 14'h3ff9; 
        10'b1001000011: data <= 14'h3fe4; 
        10'b1001000100: data <= 14'h3fde; 
        10'b1001000101: data <= 14'h3fe0; 
        10'b1001000110: data <= 14'h3fe7; 
        10'b1001000111: data <= 14'h3ffa; 
        10'b1001001000: data <= 14'h0003; 
        10'b1001001001: data <= 14'h0010; 
        10'b1001001010: data <= 14'h0006; 
        10'b1001001011: data <= 14'h0014; 
        10'b1001001100: data <= 14'h000e; 
        10'b1001001101: data <= 14'h0007; 
        10'b1001001110: data <= 14'h000b; 
        10'b1001001111: data <= 14'h000e; 
        10'b1001010000: data <= 14'h000b; 
        10'b1001010001: data <= 14'h001d; 
        10'b1001010010: data <= 14'h0018; 
        10'b1001010011: data <= 14'h000b; 
        10'b1001010100: data <= 14'h0002; 
        10'b1001010101: data <= 14'h3ff8; 
        10'b1001010110: data <= 14'h0000; 
        10'b1001010111: data <= 14'h3fef; 
        10'b1001011000: data <= 14'h3fda; 
        10'b1001011001: data <= 14'h3fd4; 
        10'b1001011010: data <= 14'h3ffc; 
        10'b1001011011: data <= 14'h000d; 
        10'b1001011100: data <= 14'h0015; 
        10'b1001011101: data <= 14'h0018; 
        10'b1001011110: data <= 14'h0010; 
        10'b1001011111: data <= 14'h3fe4; 
        10'b1001100000: data <= 14'h3fe5; 
        10'b1001100001: data <= 14'h3fe1; 
        10'b1001100010: data <= 14'h3feb; 
        10'b1001100011: data <= 14'h3ff4; 
        10'b1001100100: data <= 14'h0003; 
        10'b1001100101: data <= 14'h0008; 
        10'b1001100110: data <= 14'h0002; 
        10'b1001100111: data <= 14'h0002; 
        10'b1001101000: data <= 14'h000b; 
        10'b1001101001: data <= 14'h000b; 
        10'b1001101010: data <= 14'h000c; 
        10'b1001101011: data <= 14'h0003; 
        10'b1001101100: data <= 14'h0019; 
        10'b1001101101: data <= 14'h0038; 
        10'b1001101110: data <= 14'h003a; 
        10'b1001101111: data <= 14'h0023; 
        10'b1001110000: data <= 14'h0005; 
        10'b1001110001: data <= 14'h3ffc; 
        10'b1001110010: data <= 14'h3ff3; 
        10'b1001110011: data <= 14'h3fc8; 
        10'b1001110100: data <= 14'h3fa6; 
        10'b1001110101: data <= 14'h3fbb; 
        10'b1001110110: data <= 14'h0000; 
        10'b1001110111: data <= 14'h000e; 
        10'b1001111000: data <= 14'h0034; 
        10'b1001111001: data <= 14'h0055; 
        10'b1001111010: data <= 14'h0025; 
        10'b1001111011: data <= 14'h0008; 
        10'b1001111100: data <= 14'h3fed; 
        10'b1001111101: data <= 14'h3ff1; 
        10'b1001111110: data <= 14'h3fff; 
        10'b1001111111: data <= 14'h0003; 
        10'b1010000000: data <= 14'h0001; 
        10'b1010000001: data <= 14'h0008; 
        10'b1010000010: data <= 14'h0013; 
        10'b1010000011: data <= 14'h0009; 
        10'b1010000100: data <= 14'h0011; 
        10'b1010000101: data <= 14'h000b; 
        10'b1010000110: data <= 14'h000e; 
        10'b1010000111: data <= 14'h0008; 
        10'b1010001000: data <= 14'h0017; 
        10'b1010001001: data <= 14'h0030; 
        10'b1010001010: data <= 14'h0034; 
        10'b1010001011: data <= 14'h0018; 
        10'b1010001100: data <= 14'h0007; 
        10'b1010001101: data <= 14'h3ff4; 
        10'b1010001110: data <= 14'h3ff8; 
        10'b1010001111: data <= 14'h3fe1; 
        10'b1010010000: data <= 14'h3fea; 
        10'b1010010001: data <= 14'h3fec; 
        10'b1010010010: data <= 14'h3fe6; 
        10'b1010010011: data <= 14'h000a; 
        10'b1010010100: data <= 14'h003c; 
        10'b1010010101: data <= 14'h0049; 
        10'b1010010110: data <= 14'h0021; 
        10'b1010010111: data <= 14'h3ffa; 
        10'b1010011000: data <= 14'h3ff2; 
        10'b1010011001: data <= 14'h3feb; 
        10'b1010011010: data <= 14'h3ff9; 
        10'b1010011011: data <= 14'h3ff9; 
        10'b1010011100: data <= 14'h0004; 
        10'b1010011101: data <= 14'h0002; 
        10'b1010011110: data <= 14'h0004; 
        10'b1010011111: data <= 14'h0002; 
        10'b1010100000: data <= 14'h0004; 
        10'b1010100001: data <= 14'h0003; 
        10'b1010100010: data <= 14'h0007; 
        10'b1010100011: data <= 14'h0002; 
        10'b1010100100: data <= 14'h000b; 
        10'b1010100101: data <= 14'h0015; 
        10'b1010100110: data <= 14'h0016; 
        10'b1010100111: data <= 14'h3ff9; 
        10'b1010101000: data <= 14'h3fe0; 
        10'b1010101001: data <= 14'h3fe0; 
        10'b1010101010: data <= 14'h3fc7; 
        10'b1010101011: data <= 14'h3fca; 
        10'b1010101100: data <= 14'h3fcf; 
        10'b1010101101: data <= 14'h3fd6; 
        10'b1010101110: data <= 14'h3fd6; 
        10'b1010101111: data <= 14'h3fd6; 
        10'b1010110000: data <= 14'h3ff4; 
        10'b1010110001: data <= 14'h0005; 
        10'b1010110010: data <= 14'h0009; 
        10'b1010110011: data <= 14'h000d; 
        10'b1010110100: data <= 14'h000b; 
        10'b1010110101: data <= 14'h0003; 
        10'b1010110110: data <= 14'h0006; 
        10'b1010110111: data <= 14'h000f; 
        10'b1010111000: data <= 14'h0005; 
        10'b1010111001: data <= 14'h0008; 
        10'b1010111010: data <= 14'h000f; 
        10'b1010111011: data <= 14'h0005; 
        10'b1010111100: data <= 14'h0013; 
        10'b1010111101: data <= 14'h0006; 
        10'b1010111110: data <= 14'h0007; 
        10'b1010111111: data <= 14'h000a; 
        10'b1011000000: data <= 14'h000f; 
        10'b1011000001: data <= 14'h000d; 
        10'b1011000010: data <= 14'h0000; 
        10'b1011000011: data <= 14'h3ff8; 
        10'b1011000100: data <= 14'h3ffd; 
        10'b1011000101: data <= 14'h3ff8; 
        10'b1011000110: data <= 14'h3fe0; 
        10'b1011000111: data <= 14'h3fd9; 
        10'b1011001000: data <= 14'h3fe3; 
        10'b1011001001: data <= 14'h3fd8; 
        10'b1011001010: data <= 14'h3fe8; 
        10'b1011001011: data <= 14'h3fe1; 
        10'b1011001100: data <= 14'h3fee; 
        10'b1011001101: data <= 14'h3ffd; 
        10'b1011001110: data <= 14'h0006; 
        10'b1011001111: data <= 14'h000d; 
        10'b1011010000: data <= 14'h0001; 
        10'b1011010001: data <= 14'h000c; 
        10'b1011010010: data <= 14'h0007; 
        10'b1011010011: data <= 14'h0011; 
        10'b1011010100: data <= 14'h0004; 
        10'b1011010101: data <= 14'h0005; 
        10'b1011010110: data <= 14'h0007; 
        10'b1011010111: data <= 14'h0006; 
        10'b1011011000: data <= 14'h0007; 
        10'b1011011001: data <= 14'h000d; 
        10'b1011011010: data <= 14'h000c; 
        10'b1011011011: data <= 14'h0004; 
        10'b1011011100: data <= 14'h000d; 
        10'b1011011101: data <= 14'h0011; 
        10'b1011011110: data <= 14'h000c; 
        10'b1011011111: data <= 14'h000b; 
        10'b1011100000: data <= 14'h000f; 
        10'b1011100001: data <= 14'h000d; 
        10'b1011100010: data <= 14'h0002; 
        10'b1011100011: data <= 14'h000b; 
        10'b1011100100: data <= 14'h000a; 
        10'b1011100101: data <= 14'h0006; 
        10'b1011100110: data <= 14'h0000; 
        10'b1011100111: data <= 14'h0005; 
        10'b1011101000: data <= 14'h000b; 
        10'b1011101001: data <= 14'h0011; 
        10'b1011101010: data <= 14'h000d; 
        10'b1011101011: data <= 14'h0002; 
        10'b1011101100: data <= 14'h000c; 
        10'b1011101101: data <= 14'h000b; 
        10'b1011101110: data <= 14'h000b; 
        10'b1011101111: data <= 14'h0005; 
        10'b1011110000: data <= 14'h0004; 
        10'b1011110001: data <= 14'h000d; 
        10'b1011110010: data <= 14'h0012; 
        10'b1011110011: data <= 14'h000e; 
        10'b1011110100: data <= 14'h000e; 
        10'b1011110101: data <= 14'h0012; 
        10'b1011110110: data <= 14'h0003; 
        10'b1011110111: data <= 14'h000a; 
        10'b1011111000: data <= 14'h0013; 
        10'b1011111001: data <= 14'h000f; 
        10'b1011111010: data <= 14'h0011; 
        10'b1011111011: data <= 14'h0010; 
        10'b1011111100: data <= 14'h0011; 
        10'b1011111101: data <= 14'h0008; 
        10'b1011111110: data <= 14'h000f; 
        10'b1011111111: data <= 14'h0010; 
        10'b1100000000: data <= 14'h0002; 
        10'b1100000001: data <= 14'h0003; 
        10'b1100000010: data <= 14'h0013; 
        10'b1100000011: data <= 14'h000c; 
        10'b1100000100: data <= 14'h000b; 
        10'b1100000101: data <= 14'h0002; 
        10'b1100000110: data <= 14'h0008; 
        10'b1100000111: data <= 14'h0004; 
        10'b1100001000: data <= 14'h0003; 
        10'b1100001001: data <= 14'h0006; 
        10'b1100001010: data <= 14'h000b; 
        10'b1100001011: data <= 14'h0010; 
        10'b1100001100: data <= 14'h0012; 
        10'b1100001101: data <= 14'h0011; 
        10'b1100001110: data <= 14'h0011; 
        10'b1100001111: data <= 14'h0006; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 9) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 15'h0020; 
        10'b0000000001: data <= 15'h000f; 
        10'b0000000010: data <= 15'h0011; 
        10'b0000000011: data <= 15'h0007; 
        10'b0000000100: data <= 15'h001b; 
        10'b0000000101: data <= 15'h001a; 
        10'b0000000110: data <= 15'h001d; 
        10'b0000000111: data <= 15'h0007; 
        10'b0000001000: data <= 15'h0019; 
        10'b0000001001: data <= 15'h0008; 
        10'b0000001010: data <= 15'h0018; 
        10'b0000001011: data <= 15'h0013; 
        10'b0000001100: data <= 15'h001b; 
        10'b0000001101: data <= 15'h0024; 
        10'b0000001110: data <= 15'h0020; 
        10'b0000001111: data <= 15'h0016; 
        10'b0000010000: data <= 15'h0016; 
        10'b0000010001: data <= 15'h0008; 
        10'b0000010010: data <= 15'h0025; 
        10'b0000010011: data <= 15'h0025; 
        10'b0000010100: data <= 15'h0015; 
        10'b0000010101: data <= 15'h001b; 
        10'b0000010110: data <= 15'h0015; 
        10'b0000010111: data <= 15'h0020; 
        10'b0000011000: data <= 15'h000c; 
        10'b0000011001: data <= 15'h0022; 
        10'b0000011010: data <= 15'h0015; 
        10'b0000011011: data <= 15'h001e; 
        10'b0000011100: data <= 15'h0004; 
        10'b0000011101: data <= 15'h0020; 
        10'b0000011110: data <= 15'h0009; 
        10'b0000011111: data <= 15'h0017; 
        10'b0000100000: data <= 15'h0014; 
        10'b0000100001: data <= 15'h0008; 
        10'b0000100010: data <= 15'h000b; 
        10'b0000100011: data <= 15'h001e; 
        10'b0000100100: data <= 15'h001d; 
        10'b0000100101: data <= 15'h0018; 
        10'b0000100110: data <= 15'h0017; 
        10'b0000100111: data <= 15'h0011; 
        10'b0000101000: data <= 15'h001c; 
        10'b0000101001: data <= 15'h001f; 
        10'b0000101010: data <= 15'h0028; 
        10'b0000101011: data <= 15'h0014; 
        10'b0000101100: data <= 15'h0010; 
        10'b0000101101: data <= 15'h0020; 
        10'b0000101110: data <= 15'h0016; 
        10'b0000101111: data <= 15'h000f; 
        10'b0000110000: data <= 15'h0023; 
        10'b0000110001: data <= 15'h0022; 
        10'b0000110010: data <= 15'h000e; 
        10'b0000110011: data <= 15'h0024; 
        10'b0000110100: data <= 15'h0027; 
        10'b0000110101: data <= 15'h0015; 
        10'b0000110110: data <= 15'h0021; 
        10'b0000110111: data <= 15'h001b; 
        10'b0000111000: data <= 15'h0021; 
        10'b0000111001: data <= 15'h0019; 
        10'b0000111010: data <= 15'h0027; 
        10'b0000111011: data <= 15'h0008; 
        10'b0000111100: data <= 15'h0007; 
        10'b0000111101: data <= 15'h001a; 
        10'b0000111110: data <= 15'h0013; 
        10'b0000111111: data <= 15'h0012; 
        10'b0001000000: data <= 15'h000c; 
        10'b0001000001: data <= 15'h0016; 
        10'b0001000010: data <= 15'h0001; 
        10'b0001000011: data <= 15'h000b; 
        10'b0001000100: data <= 15'h0001; 
        10'b0001000101: data <= 15'h0009; 
        10'b0001000110: data <= 15'h0014; 
        10'b0001000111: data <= 15'h0020; 
        10'b0001001000: data <= 15'h0018; 
        10'b0001001001: data <= 15'h0000; 
        10'b0001001010: data <= 15'h0018; 
        10'b0001001011: data <= 15'h000e; 
        10'b0001001100: data <= 15'h001f; 
        10'b0001001101: data <= 15'h000e; 
        10'b0001001110: data <= 15'h0022; 
        10'b0001001111: data <= 15'h0019; 
        10'b0001010000: data <= 15'h001b; 
        10'b0001010001: data <= 15'h0005; 
        10'b0001010010: data <= 15'h001d; 
        10'b0001010011: data <= 15'h001e; 
        10'b0001010100: data <= 15'h000c; 
        10'b0001010101: data <= 15'h000d; 
        10'b0001010110: data <= 15'h0016; 
        10'b0001010111: data <= 15'h0012; 
        10'b0001011000: data <= 15'h0025; 
        10'b0001011001: data <= 15'h0013; 
        10'b0001011010: data <= 15'h0004; 
        10'b0001011011: data <= 15'h0024; 
        10'b0001011100: data <= 15'h7ffc; 
        10'b0001011101: data <= 15'h7ff9; 
        10'b0001011110: data <= 15'h7ff9; 
        10'b0001011111: data <= 15'h7fec; 
        10'b0001100000: data <= 15'h7ff9; 
        10'b0001100001: data <= 15'h0003; 
        10'b0001100010: data <= 15'h000f; 
        10'b0001100011: data <= 15'h001e; 
        10'b0001100100: data <= 15'h7ff1; 
        10'b0001100101: data <= 15'h7ffb; 
        10'b0001100110: data <= 15'h7fff; 
        10'b0001100111: data <= 15'h7fe9; 
        10'b0001101000: data <= 15'h7ffe; 
        10'b0001101001: data <= 15'h000a; 
        10'b0001101010: data <= 15'h0018; 
        10'b0001101011: data <= 15'h0017; 
        10'b0001101100: data <= 15'h7ffc; 
        10'b0001101101: data <= 15'h0021; 
        10'b0001101110: data <= 15'h000c; 
        10'b0001101111: data <= 15'h0023; 
        10'b0001110000: data <= 15'h001b; 
        10'b0001110001: data <= 15'h0010; 
        10'b0001110010: data <= 15'h0025; 
        10'b0001110011: data <= 15'h0025; 
        10'b0001110100: data <= 15'h0004; 
        10'b0001110101: data <= 15'h0007; 
        10'b0001110110: data <= 15'h0020; 
        10'b0001110111: data <= 15'h0015; 
        10'b0001111000: data <= 15'h0008; 
        10'b0001111001: data <= 15'h7fde; 
        10'b0001111010: data <= 15'h0003; 
        10'b0001111011: data <= 15'h000c; 
        10'b0001111100: data <= 15'h0012; 
        10'b0001111101: data <= 15'h0021; 
        10'b0001111110: data <= 15'h0027; 
        10'b0001111111: data <= 15'h004f; 
        10'b0010000000: data <= 15'h0016; 
        10'b0010000001: data <= 15'h7fef; 
        10'b0010000010: data <= 15'h7fee; 
        10'b0010000011: data <= 15'h000c; 
        10'b0010000100: data <= 15'h002c; 
        10'b0010000101: data <= 15'h0031; 
        10'b0010000110: data <= 15'h0031; 
        10'b0010000111: data <= 15'h0039; 
        10'b0010001000: data <= 15'h001e; 
        10'b0010001001: data <= 15'h000e; 
        10'b0010001010: data <= 15'h000c; 
        10'b0010001011: data <= 15'h000e; 
        10'b0010001100: data <= 15'h0005; 
        10'b0010001101: data <= 15'h0020; 
        10'b0010001110: data <= 15'h0006; 
        10'b0010001111: data <= 15'h0016; 
        10'b0010010000: data <= 15'h0006; 
        10'b0010010001: data <= 15'h0016; 
        10'b0010010010: data <= 15'h0006; 
        10'b0010010011: data <= 15'h7ff8; 
        10'b0010010100: data <= 15'h7fb9; 
        10'b0010010101: data <= 15'h7fb8; 
        10'b0010010110: data <= 15'h7fdf; 
        10'b0010010111: data <= 15'h0000; 
        10'b0010011000: data <= 15'h001b; 
        10'b0010011001: data <= 15'h001e; 
        10'b0010011010: data <= 15'h0035; 
        10'b0010011011: data <= 15'h0029; 
        10'b0010011100: data <= 15'h0018; 
        10'b0010011101: data <= 15'h7fd8; 
        10'b0010011110: data <= 15'h7ffc; 
        10'b0010011111: data <= 15'h0008; 
        10'b0010100000: data <= 15'h0027; 
        10'b0010100001: data <= 15'h003f; 
        10'b0010100010: data <= 15'h0069; 
        10'b0010100011: data <= 15'h0041; 
        10'b0010100100: data <= 15'h0035; 
        10'b0010100101: data <= 15'h7ff2; 
        10'b0010100110: data <= 15'h000f; 
        10'b0010100111: data <= 15'h0008; 
        10'b0010101000: data <= 15'h0007; 
        10'b0010101001: data <= 15'h0017; 
        10'b0010101010: data <= 15'h0004; 
        10'b0010101011: data <= 15'h0012; 
        10'b0010101100: data <= 15'h0004; 
        10'b0010101101: data <= 15'h7ff5; 
        10'b0010101110: data <= 15'h7fd9; 
        10'b0010101111: data <= 15'h7fd9; 
        10'b0010110000: data <= 15'h7fa7; 
        10'b0010110001: data <= 15'h7f94; 
        10'b0010110010: data <= 15'h7fbd; 
        10'b0010110011: data <= 15'h7ff0; 
        10'b0010110100: data <= 15'h7ff0; 
        10'b0010110101: data <= 15'h7fde; 
        10'b0010110110: data <= 15'h7ff0; 
        10'b0010110111: data <= 15'h7fb3; 
        10'b0010111000: data <= 15'h7fad; 
        10'b0010111001: data <= 15'h7fac; 
        10'b0010111010: data <= 15'h7fdd; 
        10'b0010111011: data <= 15'h7fe6; 
        10'b0010111100: data <= 15'h0027; 
        10'b0010111101: data <= 15'h0041; 
        10'b0010111110: data <= 15'h003c; 
        10'b0010111111: data <= 15'h0032; 
        10'b0011000000: data <= 15'h000d; 
        10'b0011000001: data <= 15'h7ff5; 
        10'b0011000010: data <= 15'h0001; 
        10'b0011000011: data <= 15'h0013; 
        10'b0011000100: data <= 15'h000f; 
        10'b0011000101: data <= 15'h0009; 
        10'b0011000110: data <= 15'h000b; 
        10'b0011000111: data <= 15'h0002; 
        10'b0011001000: data <= 15'h0019; 
        10'b0011001001: data <= 15'h7ffb; 
        10'b0011001010: data <= 15'h7fda; 
        10'b0011001011: data <= 15'h7fb3; 
        10'b0011001100: data <= 15'h7f88; 
        10'b0011001101: data <= 15'h7f67; 
        10'b0011001110: data <= 15'h7f98; 
        10'b0011001111: data <= 15'h7fd3; 
        10'b0011010000: data <= 15'h7fd6; 
        10'b0011010001: data <= 15'h7fc4; 
        10'b0011010010: data <= 15'h7fb6; 
        10'b0011010011: data <= 15'h7f8d; 
        10'b0011010100: data <= 15'h7f9c; 
        10'b0011010101: data <= 15'h7fa2; 
        10'b0011010110: data <= 15'h7fab; 
        10'b0011010111: data <= 15'h7ffd; 
        10'b0011011000: data <= 15'h0012; 
        10'b0011011001: data <= 15'h000b; 
        10'b0011011010: data <= 15'h000b; 
        10'b0011011011: data <= 15'h7fe0; 
        10'b0011011100: data <= 15'h7fd4; 
        10'b0011011101: data <= 15'h7fee; 
        10'b0011011110: data <= 15'h000e; 
        10'b0011011111: data <= 15'h0011; 
        10'b0011100000: data <= 15'h0013; 
        10'b0011100001: data <= 15'h0010; 
        10'b0011100010: data <= 15'h000f; 
        10'b0011100011: data <= 15'h0021; 
        10'b0011100100: data <= 15'h000a; 
        10'b0011100101: data <= 15'h7fff; 
        10'b0011100110: data <= 15'h7fd3; 
        10'b0011100111: data <= 15'h7fbc; 
        10'b0011101000: data <= 15'h7f74; 
        10'b0011101001: data <= 15'h7f68; 
        10'b0011101010: data <= 15'h7f6f; 
        10'b0011101011: data <= 15'h7fb2; 
        10'b0011101100: data <= 15'h7fdc; 
        10'b0011101101: data <= 15'h7fd4; 
        10'b0011101110: data <= 15'h7fdc; 
        10'b0011101111: data <= 15'h0010; 
        10'b0011110000: data <= 15'h7fc0; 
        10'b0011110001: data <= 15'h7fea; 
        10'b0011110010: data <= 15'h7ffc; 
        10'b0011110011: data <= 15'h0008; 
        10'b0011110100: data <= 15'h7fd0; 
        10'b0011110101: data <= 15'h7fd2; 
        10'b0011110110: data <= 15'h7fb6; 
        10'b0011110111: data <= 15'h7f9f; 
        10'b0011111000: data <= 15'h7fb3; 
        10'b0011111001: data <= 15'h7fed; 
        10'b0011111010: data <= 15'h001d; 
        10'b0011111011: data <= 15'h0026; 
        10'b0011111100: data <= 15'h0026; 
        10'b0011111101: data <= 15'h0009; 
        10'b0011111110: data <= 15'h0010; 
        10'b0011111111: data <= 15'h000d; 
        10'b0100000000: data <= 15'h7ffe; 
        10'b0100000001: data <= 15'h7ffc; 
        10'b0100000010: data <= 15'h7fc7; 
        10'b0100000011: data <= 15'h7fca; 
        10'b0100000100: data <= 15'h7fa0; 
        10'b0100000101: data <= 15'h7f6d; 
        10'b0100000110: data <= 15'h7f79; 
        10'b0100000111: data <= 15'h7fcb; 
        10'b0100001000: data <= 15'h7fd8; 
        10'b0100001001: data <= 15'h001e; 
        10'b0100001010: data <= 15'h005f; 
        10'b0100001011: data <= 15'h0088; 
        10'b0100001100: data <= 15'h0033; 
        10'b0100001101: data <= 15'h7ffc; 
        10'b0100001110: data <= 15'h7fe9; 
        10'b0100001111: data <= 15'h7fa4; 
        10'b0100010000: data <= 15'h7f8e; 
        10'b0100010001: data <= 15'h7f90; 
        10'b0100010010: data <= 15'h7f73; 
        10'b0100010011: data <= 15'h7f86; 
        10'b0100010100: data <= 15'h7fbe; 
        10'b0100010101: data <= 15'h0008; 
        10'b0100010110: data <= 15'h0020; 
        10'b0100010111: data <= 15'h0017; 
        10'b0100011000: data <= 15'h0023; 
        10'b0100011001: data <= 15'h0027; 
        10'b0100011010: data <= 15'h0020; 
        10'b0100011011: data <= 15'h0004; 
        10'b0100011100: data <= 15'h001a; 
        10'b0100011101: data <= 15'h7fe2; 
        10'b0100011110: data <= 15'h7fca; 
        10'b0100011111: data <= 15'h7fe7; 
        10'b0100100000: data <= 15'h7fb5; 
        10'b0100100001: data <= 15'h7fb4; 
        10'b0100100010: data <= 15'h7fc9; 
        10'b0100100011: data <= 15'h7fdb; 
        10'b0100100100: data <= 15'h7fe7; 
        10'b0100100101: data <= 15'h004c; 
        10'b0100100110: data <= 15'h00f6; 
        10'b0100100111: data <= 15'h0104; 
        10'b0100101000: data <= 15'h007b; 
        10'b0100101001: data <= 15'h7ffd; 
        10'b0100101010: data <= 15'h7fb6; 
        10'b0100101011: data <= 15'h7fa7; 
        10'b0100101100: data <= 15'h7f94; 
        10'b0100101101: data <= 15'h7f9f; 
        10'b0100101110: data <= 15'h7fa4; 
        10'b0100101111: data <= 15'h7fc7; 
        10'b0100110000: data <= 15'h7fed; 
        10'b0100110001: data <= 15'h7ffd; 
        10'b0100110010: data <= 15'h0021; 
        10'b0100110011: data <= 15'h000e; 
        10'b0100110100: data <= 15'h0007; 
        10'b0100110101: data <= 15'h0006; 
        10'b0100110110: data <= 15'h001b; 
        10'b0100110111: data <= 15'h001c; 
        10'b0100111000: data <= 15'h0000; 
        10'b0100111001: data <= 15'h7ff7; 
        10'b0100111010: data <= 15'h7ffc; 
        10'b0100111011: data <= 15'h7fd1; 
        10'b0100111100: data <= 15'h7fe2; 
        10'b0100111101: data <= 15'h7fd1; 
        10'b0100111110: data <= 15'h7fbb; 
        10'b0100111111: data <= 15'h7f98; 
        10'b0101000000: data <= 15'h7ff4; 
        10'b0101000001: data <= 15'h0082; 
        10'b0101000010: data <= 15'h0129; 
        10'b0101000011: data <= 15'h013a; 
        10'b0101000100: data <= 15'h0074; 
        10'b0101000101: data <= 15'h7fe7; 
        10'b0101000110: data <= 15'h7fe9; 
        10'b0101000111: data <= 15'h7fc2; 
        10'b0101001000: data <= 15'h7fbe; 
        10'b0101001001: data <= 15'h7fc3; 
        10'b0101001010: data <= 15'h7fc8; 
        10'b0101001011: data <= 15'h7fe6; 
        10'b0101001100: data <= 15'h7ff5; 
        10'b0101001101: data <= 15'h001a; 
        10'b0101001110: data <= 15'h0025; 
        10'b0101001111: data <= 15'h001a; 
        10'b0101010000: data <= 15'h0004; 
        10'b0101010001: data <= 15'h0023; 
        10'b0101010010: data <= 15'h0011; 
        10'b0101010011: data <= 15'h000b; 
        10'b0101010100: data <= 15'h0024; 
        10'b0101010101: data <= 15'h7ff9; 
        10'b0101010110: data <= 15'h7ff5; 
        10'b0101010111: data <= 15'h7ff0; 
        10'b0101011000: data <= 15'h7fd3; 
        10'b0101011001: data <= 15'h7fc6; 
        10'b0101011010: data <= 15'h7f84; 
        10'b0101011011: data <= 15'h7f52; 
        10'b0101011100: data <= 15'h7ffa; 
        10'b0101011101: data <= 15'h0084; 
        10'b0101011110: data <= 15'h015d; 
        10'b0101011111: data <= 15'h00f2; 
        10'b0101100000: data <= 15'h0030; 
        10'b0101100001: data <= 15'h0019; 
        10'b0101100010: data <= 15'h7ff1; 
        10'b0101100011: data <= 15'h7fb9; 
        10'b0101100100: data <= 15'h7fd3; 
        10'b0101100101: data <= 15'h7fea; 
        10'b0101100110: data <= 15'h7ff4; 
        10'b0101100111: data <= 15'h7ff1; 
        10'b0101101000: data <= 15'h0002; 
        10'b0101101001: data <= 15'h0024; 
        10'b0101101010: data <= 15'h0005; 
        10'b0101101011: data <= 15'h0019; 
        10'b0101101100: data <= 15'h0004; 
        10'b0101101101: data <= 15'h0018; 
        10'b0101101110: data <= 15'h0016; 
        10'b0101101111: data <= 15'h0018; 
        10'b0101110000: data <= 15'h0027; 
        10'b0101110001: data <= 15'h0000; 
        10'b0101110010: data <= 15'h0003; 
        10'b0101110011: data <= 15'h7fee; 
        10'b0101110100: data <= 15'h7fe8; 
        10'b0101110101: data <= 15'h7f9f; 
        10'b0101110110: data <= 15'h7f31; 
        10'b0101110111: data <= 15'h7f2e; 
        10'b0101111000: data <= 15'h0000; 
        10'b0101111001: data <= 15'h006e; 
        10'b0101111010: data <= 15'h0120; 
        10'b0101111011: data <= 15'h00a3; 
        10'b0101111100: data <= 15'h002b; 
        10'b0101111101: data <= 15'h0015; 
        10'b0101111110: data <= 15'h7fbe; 
        10'b0101111111: data <= 15'h7fa1; 
        10'b0110000000: data <= 15'h7fdd; 
        10'b0110000001: data <= 15'h7ff4; 
        10'b0110000010: data <= 15'h7ff3; 
        10'b0110000011: data <= 15'h7ffb; 
        10'b0110000100: data <= 15'h0010; 
        10'b0110000101: data <= 15'h0018; 
        10'b0110000110: data <= 15'h0023; 
        10'b0110000111: data <= 15'h0016; 
        10'b0110001000: data <= 15'h0012; 
        10'b0110001001: data <= 15'h0025; 
        10'b0110001010: data <= 15'h0015; 
        10'b0110001011: data <= 15'h001e; 
        10'b0110001100: data <= 15'h001e; 
        10'b0110001101: data <= 15'h0000; 
        10'b0110001110: data <= 15'h0005; 
        10'b0110001111: data <= 15'h7ff4; 
        10'b0110010000: data <= 15'h7fc0; 
        10'b0110010001: data <= 15'h7f91; 
        10'b0110010010: data <= 15'h7f32; 
        10'b0110010011: data <= 15'h7f64; 
        10'b0110010100: data <= 15'h7ffd; 
        10'b0110010101: data <= 15'h0070; 
        10'b0110010110: data <= 15'h00f5; 
        10'b0110010111: data <= 15'h009e; 
        10'b0110011000: data <= 15'h002f; 
        10'b0110011001: data <= 15'h7fa8; 
        10'b0110011010: data <= 15'h7f89; 
        10'b0110011011: data <= 15'h7fa6; 
        10'b0110011100: data <= 15'h7fcb; 
        10'b0110011101: data <= 15'h7ff1; 
        10'b0110011110: data <= 15'h7fef; 
        10'b0110011111: data <= 15'h7ff5; 
        10'b0110100000: data <= 15'h001b; 
        10'b0110100001: data <= 15'h0004; 
        10'b0110100010: data <= 15'h0007; 
        10'b0110100011: data <= 15'h0015; 
        10'b0110100100: data <= 15'h0028; 
        10'b0110100101: data <= 15'h0007; 
        10'b0110100110: data <= 15'h0019; 
        10'b0110100111: data <= 15'h0010; 
        10'b0110101000: data <= 15'h0009; 
        10'b0110101001: data <= 15'h0017; 
        10'b0110101010: data <= 15'h7fe9; 
        10'b0110101011: data <= 15'h7fe6; 
        10'b0110101100: data <= 15'h7fd7; 
        10'b0110101101: data <= 15'h7f87; 
        10'b0110101110: data <= 15'h7f78; 
        10'b0110101111: data <= 15'h7fde; 
        10'b0110110000: data <= 15'h0032; 
        10'b0110110001: data <= 15'h009d; 
        10'b0110110010: data <= 15'h0107; 
        10'b0110110011: data <= 15'h005d; 
        10'b0110110100: data <= 15'h0011; 
        10'b0110110101: data <= 15'h7f5b; 
        10'b0110110110: data <= 15'h7f6e; 
        10'b0110110111: data <= 15'h7fa6; 
        10'b0110111000: data <= 15'h7fca; 
        10'b0110111001: data <= 15'h7fd9; 
        10'b0110111010: data <= 15'h7ff6; 
        10'b0110111011: data <= 15'h0003; 
        10'b0110111100: data <= 15'h000e; 
        10'b0110111101: data <= 15'h0012; 
        10'b0110111110: data <= 15'h0025; 
        10'b0110111111: data <= 15'h0006; 
        10'b0111000000: data <= 15'h0026; 
        10'b0111000001: data <= 15'h0013; 
        10'b0111000010: data <= 15'h0023; 
        10'b0111000011: data <= 15'h0015; 
        10'b0111000100: data <= 15'h000b; 
        10'b0111000101: data <= 15'h7ff0; 
        10'b0111000110: data <= 15'h7fdc; 
        10'b0111000111: data <= 15'h7fda; 
        10'b0111001000: data <= 15'h7fa2; 
        10'b0111001001: data <= 15'h7fc8; 
        10'b0111001010: data <= 15'h7fd3; 
        10'b0111001011: data <= 15'h7fe7; 
        10'b0111001100: data <= 15'h7ffa; 
        10'b0111001101: data <= 15'h00cf; 
        10'b0111001110: data <= 15'h00f8; 
        10'b0111001111: data <= 15'h000e; 
        10'b0111010000: data <= 15'h7fb3; 
        10'b0111010001: data <= 15'h7f4d; 
        10'b0111010010: data <= 15'h7f6c; 
        10'b0111010011: data <= 15'h7fa1; 
        10'b0111010100: data <= 15'h7fb8; 
        10'b0111010101: data <= 15'h7fe1; 
        10'b0111010110: data <= 15'h7fe1; 
        10'b0111010111: data <= 15'h0000; 
        10'b0111011000: data <= 15'h7ff2; 
        10'b0111011001: data <= 15'h0002; 
        10'b0111011010: data <= 15'h0009; 
        10'b0111011011: data <= 15'h0014; 
        10'b0111011100: data <= 15'h0010; 
        10'b0111011101: data <= 15'h0026; 
        10'b0111011110: data <= 15'h0008; 
        10'b0111011111: data <= 15'h0025; 
        10'b0111100000: data <= 15'h001c; 
        10'b0111100001: data <= 15'h7fea; 
        10'b0111100010: data <= 15'h7fb2; 
        10'b0111100011: data <= 15'h7fab; 
        10'b0111100100: data <= 15'h7fc3; 
        10'b0111100101: data <= 15'h7fd9; 
        10'b0111100110: data <= 15'h001c; 
        10'b0111100111: data <= 15'h0000; 
        10'b0111101000: data <= 15'h0043; 
        10'b0111101001: data <= 15'h00ed; 
        10'b0111101010: data <= 15'h00cb; 
        10'b0111101011: data <= 15'h7fd7; 
        10'b0111101100: data <= 15'h7f73; 
        10'b0111101101: data <= 15'h7f4d; 
        10'b0111101110: data <= 15'h7f6d; 
        10'b0111101111: data <= 15'h7fa3; 
        10'b0111110000: data <= 15'h7fdd; 
        10'b0111110001: data <= 15'h7fee; 
        10'b0111110010: data <= 15'h7ff3; 
        10'b0111110011: data <= 15'h7fef; 
        10'b0111110100: data <= 15'h7fe3; 
        10'b0111110101: data <= 15'h0008; 
        10'b0111110110: data <= 15'h0016; 
        10'b0111110111: data <= 15'h001a; 
        10'b0111111000: data <= 15'h0017; 
        10'b0111111001: data <= 15'h0016; 
        10'b0111111010: data <= 15'h000d; 
        10'b0111111011: data <= 15'h001f; 
        10'b0111111100: data <= 15'h0011; 
        10'b0111111101: data <= 15'h7fe1; 
        10'b0111111110: data <= 15'h7fac; 
        10'b0111111111: data <= 15'h7fad; 
        10'b1000000000: data <= 15'h7fe1; 
        10'b1000000001: data <= 15'h0020; 
        10'b1000000010: data <= 15'h001a; 
        10'b1000000011: data <= 15'h002a; 
        10'b1000000100: data <= 15'h006e; 
        10'b1000000101: data <= 15'h00b1; 
        10'b1000000110: data <= 15'h007a; 
        10'b1000000111: data <= 15'h7fb0; 
        10'b1000001000: data <= 15'h7f7c; 
        10'b1000001001: data <= 15'h7f8f; 
        10'b1000001010: data <= 15'h7f9f; 
        10'b1000001011: data <= 15'h7fbf; 
        10'b1000001100: data <= 15'h7fe0; 
        10'b1000001101: data <= 15'h7fca; 
        10'b1000001110: data <= 15'h7fe8; 
        10'b1000001111: data <= 15'h7fdb; 
        10'b1000010000: data <= 15'h7fea; 
        10'b1000010001: data <= 15'h0014; 
        10'b1000010010: data <= 15'h0023; 
        10'b1000010011: data <= 15'h0024; 
        10'b1000010100: data <= 15'h0025; 
        10'b1000010101: data <= 15'h001a; 
        10'b1000010110: data <= 15'h001b; 
        10'b1000010111: data <= 15'h001e; 
        10'b1000011000: data <= 15'h0003; 
        10'b1000011001: data <= 15'h7fd1; 
        10'b1000011010: data <= 15'h7f98; 
        10'b1000011011: data <= 15'h7fba; 
        10'b1000011100: data <= 15'h7fe3; 
        10'b1000011101: data <= 15'h0010; 
        10'b1000011110: data <= 15'h0008; 
        10'b1000011111: data <= 15'h0006; 
        10'b1000100000: data <= 15'h000f; 
        10'b1000100001: data <= 15'h0051; 
        10'b1000100010: data <= 15'h0012; 
        10'b1000100011: data <= 15'h7fbe; 
        10'b1000100100: data <= 15'h7fc9; 
        10'b1000100101: data <= 15'h7fd0; 
        10'b1000100110: data <= 15'h7fc4; 
        10'b1000100111: data <= 15'h7fd1; 
        10'b1000101000: data <= 15'h7fbb; 
        10'b1000101001: data <= 15'h7fc7; 
        10'b1000101010: data <= 15'h7fdd; 
        10'b1000101011: data <= 15'h7fe2; 
        10'b1000101100: data <= 15'h0002; 
        10'b1000101101: data <= 15'h000c; 
        10'b1000101110: data <= 15'h000d; 
        10'b1000101111: data <= 15'h0005; 
        10'b1000110000: data <= 15'h0006; 
        10'b1000110001: data <= 15'h0027; 
        10'b1000110010: data <= 15'h0015; 
        10'b1000110011: data <= 15'h000d; 
        10'b1000110100: data <= 15'h7ff6; 
        10'b1000110101: data <= 15'h7fdf; 
        10'b1000110110: data <= 15'h7ffa; 
        10'b1000110111: data <= 15'h7fe9; 
        10'b1000111000: data <= 15'h7fff; 
        10'b1000111001: data <= 15'h000a; 
        10'b1000111010: data <= 15'h7fe6; 
        10'b1000111011: data <= 15'h7ff7; 
        10'b1000111100: data <= 15'h7fd6; 
        10'b1000111101: data <= 15'h7ff2; 
        10'b1000111110: data <= 15'h7ff6; 
        10'b1000111111: data <= 15'h0003; 
        10'b1001000000: data <= 15'h0028; 
        10'b1001000001: data <= 15'h000e; 
        10'b1001000010: data <= 15'h7ff1; 
        10'b1001000011: data <= 15'h7fc8; 
        10'b1001000100: data <= 15'h7fbc; 
        10'b1001000101: data <= 15'h7fc1; 
        10'b1001000110: data <= 15'h7fce; 
        10'b1001000111: data <= 15'h7ff5; 
        10'b1001001000: data <= 15'h0005; 
        10'b1001001001: data <= 15'h0020; 
        10'b1001001010: data <= 15'h000d; 
        10'b1001001011: data <= 15'h0027; 
        10'b1001001100: data <= 15'h001c; 
        10'b1001001101: data <= 15'h000f; 
        10'b1001001110: data <= 15'h0017; 
        10'b1001001111: data <= 15'h001b; 
        10'b1001010000: data <= 15'h0016; 
        10'b1001010001: data <= 15'h003a; 
        10'b1001010010: data <= 15'h0030; 
        10'b1001010011: data <= 15'h0017; 
        10'b1001010100: data <= 15'h0004; 
        10'b1001010101: data <= 15'h7fef; 
        10'b1001010110: data <= 15'h0001; 
        10'b1001010111: data <= 15'h7fde; 
        10'b1001011000: data <= 15'h7fb4; 
        10'b1001011001: data <= 15'h7fa9; 
        10'b1001011010: data <= 15'h7ff8; 
        10'b1001011011: data <= 15'h001a; 
        10'b1001011100: data <= 15'h002a; 
        10'b1001011101: data <= 15'h0030; 
        10'b1001011110: data <= 15'h0021; 
        10'b1001011111: data <= 15'h7fc9; 
        10'b1001100000: data <= 15'h7fca; 
        10'b1001100001: data <= 15'h7fc2; 
        10'b1001100010: data <= 15'h7fd5; 
        10'b1001100011: data <= 15'h7fe7; 
        10'b1001100100: data <= 15'h0006; 
        10'b1001100101: data <= 15'h0011; 
        10'b1001100110: data <= 15'h0003; 
        10'b1001100111: data <= 15'h0005; 
        10'b1001101000: data <= 15'h0016; 
        10'b1001101001: data <= 15'h0016; 
        10'b1001101010: data <= 15'h0019; 
        10'b1001101011: data <= 15'h0005; 
        10'b1001101100: data <= 15'h0032; 
        10'b1001101101: data <= 15'h0071; 
        10'b1001101110: data <= 15'h0075; 
        10'b1001101111: data <= 15'h0046; 
        10'b1001110000: data <= 15'h000a; 
        10'b1001110001: data <= 15'h7ff8; 
        10'b1001110010: data <= 15'h7fe5; 
        10'b1001110011: data <= 15'h7f91; 
        10'b1001110100: data <= 15'h7f4c; 
        10'b1001110101: data <= 15'h7f76; 
        10'b1001110110: data <= 15'h0000; 
        10'b1001110111: data <= 15'h001b; 
        10'b1001111000: data <= 15'h0067; 
        10'b1001111001: data <= 15'h00aa; 
        10'b1001111010: data <= 15'h004a; 
        10'b1001111011: data <= 15'h000f; 
        10'b1001111100: data <= 15'h7fda; 
        10'b1001111101: data <= 15'h7fe2; 
        10'b1001111110: data <= 15'h7ffd; 
        10'b1001111111: data <= 15'h0005; 
        10'b1010000000: data <= 15'h0002; 
        10'b1010000001: data <= 15'h0010; 
        10'b1010000010: data <= 15'h0026; 
        10'b1010000011: data <= 15'h0012; 
        10'b1010000100: data <= 15'h0023; 
        10'b1010000101: data <= 15'h0016; 
        10'b1010000110: data <= 15'h001c; 
        10'b1010000111: data <= 15'h0010; 
        10'b1010001000: data <= 15'h002d; 
        10'b1010001001: data <= 15'h0061; 
        10'b1010001010: data <= 15'h0067; 
        10'b1010001011: data <= 15'h002f; 
        10'b1010001100: data <= 15'h000d; 
        10'b1010001101: data <= 15'h7fe8; 
        10'b1010001110: data <= 15'h7ff0; 
        10'b1010001111: data <= 15'h7fc1; 
        10'b1010010000: data <= 15'h7fd4; 
        10'b1010010001: data <= 15'h7fd9; 
        10'b1010010010: data <= 15'h7fcc; 
        10'b1010010011: data <= 15'h0015; 
        10'b1010010100: data <= 15'h0078; 
        10'b1010010101: data <= 15'h0091; 
        10'b1010010110: data <= 15'h0041; 
        10'b1010010111: data <= 15'h7ff4; 
        10'b1010011000: data <= 15'h7fe4; 
        10'b1010011001: data <= 15'h7fd5; 
        10'b1010011010: data <= 15'h7ff1; 
        10'b1010011011: data <= 15'h7ff2; 
        10'b1010011100: data <= 15'h0009; 
        10'b1010011101: data <= 15'h0004; 
        10'b1010011110: data <= 15'h0008; 
        10'b1010011111: data <= 15'h0004; 
        10'b1010100000: data <= 15'h0008; 
        10'b1010100001: data <= 15'h0005; 
        10'b1010100010: data <= 15'h000e; 
        10'b1010100011: data <= 15'h0004; 
        10'b1010100100: data <= 15'h0016; 
        10'b1010100101: data <= 15'h002b; 
        10'b1010100110: data <= 15'h002c; 
        10'b1010100111: data <= 15'h7ff2; 
        10'b1010101000: data <= 15'h7fc0; 
        10'b1010101001: data <= 15'h7fc0; 
        10'b1010101010: data <= 15'h7f8f; 
        10'b1010101011: data <= 15'h7f93; 
        10'b1010101100: data <= 15'h7f9f; 
        10'b1010101101: data <= 15'h7fad; 
        10'b1010101110: data <= 15'h7fad; 
        10'b1010101111: data <= 15'h7fad; 
        10'b1010110000: data <= 15'h7fe8; 
        10'b1010110001: data <= 15'h000a; 
        10'b1010110010: data <= 15'h0012; 
        10'b1010110011: data <= 15'h001b; 
        10'b1010110100: data <= 15'h0016; 
        10'b1010110101: data <= 15'h0005; 
        10'b1010110110: data <= 15'h000c; 
        10'b1010110111: data <= 15'h001f; 
        10'b1010111000: data <= 15'h0009; 
        10'b1010111001: data <= 15'h000f; 
        10'b1010111010: data <= 15'h001d; 
        10'b1010111011: data <= 15'h000a; 
        10'b1010111100: data <= 15'h0026; 
        10'b1010111101: data <= 15'h000c; 
        10'b1010111110: data <= 15'h000e; 
        10'b1010111111: data <= 15'h0014; 
        10'b1011000000: data <= 15'h001d; 
        10'b1011000001: data <= 15'h001b; 
        10'b1011000010: data <= 15'h0000; 
        10'b1011000011: data <= 15'h7fef; 
        10'b1011000100: data <= 15'h7ff9; 
        10'b1011000101: data <= 15'h7ff1; 
        10'b1011000110: data <= 15'h7fc1; 
        10'b1011000111: data <= 15'h7fb3; 
        10'b1011001000: data <= 15'h7fc7; 
        10'b1011001001: data <= 15'h7fb0; 
        10'b1011001010: data <= 15'h7fcf; 
        10'b1011001011: data <= 15'h7fc2; 
        10'b1011001100: data <= 15'h7fdc; 
        10'b1011001101: data <= 15'h7ffa; 
        10'b1011001110: data <= 15'h000c; 
        10'b1011001111: data <= 15'h001a; 
        10'b1011010000: data <= 15'h0002; 
        10'b1011010001: data <= 15'h0017; 
        10'b1011010010: data <= 15'h000e; 
        10'b1011010011: data <= 15'h0021; 
        10'b1011010100: data <= 15'h0008; 
        10'b1011010101: data <= 15'h000a; 
        10'b1011010110: data <= 15'h000e; 
        10'b1011010111: data <= 15'h000c; 
        10'b1011011000: data <= 15'h000e; 
        10'b1011011001: data <= 15'h001b; 
        10'b1011011010: data <= 15'h0018; 
        10'b1011011011: data <= 15'h0007; 
        10'b1011011100: data <= 15'h001a; 
        10'b1011011101: data <= 15'h0022; 
        10'b1011011110: data <= 15'h0017; 
        10'b1011011111: data <= 15'h0015; 
        10'b1011100000: data <= 15'h001f; 
        10'b1011100001: data <= 15'h001a; 
        10'b1011100010: data <= 15'h0004; 
        10'b1011100011: data <= 15'h0015; 
        10'b1011100100: data <= 15'h0013; 
        10'b1011100101: data <= 15'h000b; 
        10'b1011100110: data <= 15'h7fff; 
        10'b1011100111: data <= 15'h000a; 
        10'b1011101000: data <= 15'h0017; 
        10'b1011101001: data <= 15'h0023; 
        10'b1011101010: data <= 15'h001a; 
        10'b1011101011: data <= 15'h0004; 
        10'b1011101100: data <= 15'h0018; 
        10'b1011101101: data <= 15'h0016; 
        10'b1011101110: data <= 15'h0015; 
        10'b1011101111: data <= 15'h000a; 
        10'b1011110000: data <= 15'h0009; 
        10'b1011110001: data <= 15'h001a; 
        10'b1011110010: data <= 15'h0023; 
        10'b1011110011: data <= 15'h001d; 
        10'b1011110100: data <= 15'h001d; 
        10'b1011110101: data <= 15'h0025; 
        10'b1011110110: data <= 15'h0006; 
        10'b1011110111: data <= 15'h0014; 
        10'b1011111000: data <= 15'h0026; 
        10'b1011111001: data <= 15'h001f; 
        10'b1011111010: data <= 15'h0023; 
        10'b1011111011: data <= 15'h0020; 
        10'b1011111100: data <= 15'h0023; 
        10'b1011111101: data <= 15'h0010; 
        10'b1011111110: data <= 15'h001e; 
        10'b1011111111: data <= 15'h0020; 
        10'b1100000000: data <= 15'h0003; 
        10'b1100000001: data <= 15'h0007; 
        10'b1100000010: data <= 15'h0026; 
        10'b1100000011: data <= 15'h0019; 
        10'b1100000100: data <= 15'h0017; 
        10'b1100000101: data <= 15'h0003; 
        10'b1100000110: data <= 15'h0010; 
        10'b1100000111: data <= 15'h0007; 
        10'b1100001000: data <= 15'h0007; 
        10'b1100001001: data <= 15'h000c; 
        10'b1100001010: data <= 15'h0016; 
        10'b1100001011: data <= 15'h0020; 
        10'b1100001100: data <= 15'h0023; 
        10'b1100001101: data <= 15'h0023; 
        10'b1100001110: data <= 15'h0022; 
        10'b1100001111: data <= 15'h000b; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 10) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 16'h0040; 
        10'b0000000001: data <= 16'h001e; 
        10'b0000000010: data <= 16'h0022; 
        10'b0000000011: data <= 16'h000e; 
        10'b0000000100: data <= 16'h0036; 
        10'b0000000101: data <= 16'h0035; 
        10'b0000000110: data <= 16'h003a; 
        10'b0000000111: data <= 16'h000e; 
        10'b0000001000: data <= 16'h0033; 
        10'b0000001001: data <= 16'h0010; 
        10'b0000001010: data <= 16'h0030; 
        10'b0000001011: data <= 16'h0027; 
        10'b0000001100: data <= 16'h0036; 
        10'b0000001101: data <= 16'h0048; 
        10'b0000001110: data <= 16'h0040; 
        10'b0000001111: data <= 16'h002c; 
        10'b0000010000: data <= 16'h002c; 
        10'b0000010001: data <= 16'h0010; 
        10'b0000010010: data <= 16'h004a; 
        10'b0000010011: data <= 16'h004a; 
        10'b0000010100: data <= 16'h002a; 
        10'b0000010101: data <= 16'h0036; 
        10'b0000010110: data <= 16'h002a; 
        10'b0000010111: data <= 16'h0041; 
        10'b0000011000: data <= 16'h0019; 
        10'b0000011001: data <= 16'h0045; 
        10'b0000011010: data <= 16'h002a; 
        10'b0000011011: data <= 16'h003c; 
        10'b0000011100: data <= 16'h0008; 
        10'b0000011101: data <= 16'h0040; 
        10'b0000011110: data <= 16'h0013; 
        10'b0000011111: data <= 16'h002e; 
        10'b0000100000: data <= 16'h0029; 
        10'b0000100001: data <= 16'h0010; 
        10'b0000100010: data <= 16'h0017; 
        10'b0000100011: data <= 16'h003c; 
        10'b0000100100: data <= 16'h003a; 
        10'b0000100101: data <= 16'h002f; 
        10'b0000100110: data <= 16'h002f; 
        10'b0000100111: data <= 16'h0022; 
        10'b0000101000: data <= 16'h0037; 
        10'b0000101001: data <= 16'h003e; 
        10'b0000101010: data <= 16'h0051; 
        10'b0000101011: data <= 16'h0028; 
        10'b0000101100: data <= 16'h0020; 
        10'b0000101101: data <= 16'h0041; 
        10'b0000101110: data <= 16'h002c; 
        10'b0000101111: data <= 16'h001e; 
        10'b0000110000: data <= 16'h0046; 
        10'b0000110001: data <= 16'h0044; 
        10'b0000110010: data <= 16'h001c; 
        10'b0000110011: data <= 16'h0049; 
        10'b0000110100: data <= 16'h004e; 
        10'b0000110101: data <= 16'h0029; 
        10'b0000110110: data <= 16'h0042; 
        10'b0000110111: data <= 16'h0035; 
        10'b0000111000: data <= 16'h0041; 
        10'b0000111001: data <= 16'h0031; 
        10'b0000111010: data <= 16'h004e; 
        10'b0000111011: data <= 16'h000f; 
        10'b0000111100: data <= 16'h000f; 
        10'b0000111101: data <= 16'h0033; 
        10'b0000111110: data <= 16'h0026; 
        10'b0000111111: data <= 16'h0025; 
        10'b0001000000: data <= 16'h0019; 
        10'b0001000001: data <= 16'h002b; 
        10'b0001000010: data <= 16'h0001; 
        10'b0001000011: data <= 16'h0016; 
        10'b0001000100: data <= 16'h0003; 
        10'b0001000101: data <= 16'h0013; 
        10'b0001000110: data <= 16'h0028; 
        10'b0001000111: data <= 16'h0040; 
        10'b0001001000: data <= 16'h0030; 
        10'b0001001001: data <= 16'h0000; 
        10'b0001001010: data <= 16'h0030; 
        10'b0001001011: data <= 16'h001d; 
        10'b0001001100: data <= 16'h003f; 
        10'b0001001101: data <= 16'h001b; 
        10'b0001001110: data <= 16'h0045; 
        10'b0001001111: data <= 16'h0032; 
        10'b0001010000: data <= 16'h0036; 
        10'b0001010001: data <= 16'h0009; 
        10'b0001010010: data <= 16'h003b; 
        10'b0001010011: data <= 16'h003c; 
        10'b0001010100: data <= 16'h0017; 
        10'b0001010101: data <= 16'h001a; 
        10'b0001010110: data <= 16'h002c; 
        10'b0001010111: data <= 16'h0024; 
        10'b0001011000: data <= 16'h004a; 
        10'b0001011001: data <= 16'h0027; 
        10'b0001011010: data <= 16'h0008; 
        10'b0001011011: data <= 16'h0048; 
        10'b0001011100: data <= 16'hfff8; 
        10'b0001011101: data <= 16'hfff1; 
        10'b0001011110: data <= 16'hfff2; 
        10'b0001011111: data <= 16'hffd8; 
        10'b0001100000: data <= 16'hfff2; 
        10'b0001100001: data <= 16'h0005; 
        10'b0001100010: data <= 16'h001e; 
        10'b0001100011: data <= 16'h003c; 
        10'b0001100100: data <= 16'hffe2; 
        10'b0001100101: data <= 16'hfff5; 
        10'b0001100110: data <= 16'hfffe; 
        10'b0001100111: data <= 16'hffd2; 
        10'b0001101000: data <= 16'hfffb; 
        10'b0001101001: data <= 16'h0013; 
        10'b0001101010: data <= 16'h0030; 
        10'b0001101011: data <= 16'h002f; 
        10'b0001101100: data <= 16'hfff7; 
        10'b0001101101: data <= 16'h0042; 
        10'b0001101110: data <= 16'h0019; 
        10'b0001101111: data <= 16'h0046; 
        10'b0001110000: data <= 16'h0036; 
        10'b0001110001: data <= 16'h0021; 
        10'b0001110010: data <= 16'h004a; 
        10'b0001110011: data <= 16'h004a; 
        10'b0001110100: data <= 16'h0008; 
        10'b0001110101: data <= 16'h000f; 
        10'b0001110110: data <= 16'h0041; 
        10'b0001110111: data <= 16'h0029; 
        10'b0001111000: data <= 16'h0010; 
        10'b0001111001: data <= 16'hffbc; 
        10'b0001111010: data <= 16'h0006; 
        10'b0001111011: data <= 16'h0018; 
        10'b0001111100: data <= 16'h0025; 
        10'b0001111101: data <= 16'h0042; 
        10'b0001111110: data <= 16'h004d; 
        10'b0001111111: data <= 16'h009e; 
        10'b0010000000: data <= 16'h002b; 
        10'b0010000001: data <= 16'hffdf; 
        10'b0010000010: data <= 16'hffdc; 
        10'b0010000011: data <= 16'h0019; 
        10'b0010000100: data <= 16'h0058; 
        10'b0010000101: data <= 16'h0062; 
        10'b0010000110: data <= 16'h0062; 
        10'b0010000111: data <= 16'h0072; 
        10'b0010001000: data <= 16'h003c; 
        10'b0010001001: data <= 16'h001c; 
        10'b0010001010: data <= 16'h0019; 
        10'b0010001011: data <= 16'h001b; 
        10'b0010001100: data <= 16'h000a; 
        10'b0010001101: data <= 16'h0040; 
        10'b0010001110: data <= 16'h000c; 
        10'b0010001111: data <= 16'h002d; 
        10'b0010010000: data <= 16'h000b; 
        10'b0010010001: data <= 16'h002b; 
        10'b0010010010: data <= 16'h000d; 
        10'b0010010011: data <= 16'hffef; 
        10'b0010010100: data <= 16'hff71; 
        10'b0010010101: data <= 16'hff70; 
        10'b0010010110: data <= 16'hffbe; 
        10'b0010010111: data <= 16'h0001; 
        10'b0010011000: data <= 16'h0036; 
        10'b0010011001: data <= 16'h003d; 
        10'b0010011010: data <= 16'h006a; 
        10'b0010011011: data <= 16'h0052; 
        10'b0010011100: data <= 16'h0031; 
        10'b0010011101: data <= 16'hffb0; 
        10'b0010011110: data <= 16'hfff8; 
        10'b0010011111: data <= 16'h0011; 
        10'b0010100000: data <= 16'h004e; 
        10'b0010100001: data <= 16'h007e; 
        10'b0010100010: data <= 16'h00d1; 
        10'b0010100011: data <= 16'h0082; 
        10'b0010100100: data <= 16'h006b; 
        10'b0010100101: data <= 16'hffe4; 
        10'b0010100110: data <= 16'h001e; 
        10'b0010100111: data <= 16'h0010; 
        10'b0010101000: data <= 16'h000e; 
        10'b0010101001: data <= 16'h002e; 
        10'b0010101010: data <= 16'h0009; 
        10'b0010101011: data <= 16'h0024; 
        10'b0010101100: data <= 16'h0008; 
        10'b0010101101: data <= 16'hffeb; 
        10'b0010101110: data <= 16'hffb2; 
        10'b0010101111: data <= 16'hffb2; 
        10'b0010110000: data <= 16'hff4e; 
        10'b0010110001: data <= 16'hff29; 
        10'b0010110010: data <= 16'hff79; 
        10'b0010110011: data <= 16'hffe0; 
        10'b0010110100: data <= 16'hffdf; 
        10'b0010110101: data <= 16'hffbc; 
        10'b0010110110: data <= 16'hffe1; 
        10'b0010110111: data <= 16'hff65; 
        10'b0010111000: data <= 16'hff5a; 
        10'b0010111001: data <= 16'hff58; 
        10'b0010111010: data <= 16'hffba; 
        10'b0010111011: data <= 16'hffcc; 
        10'b0010111100: data <= 16'h004e; 
        10'b0010111101: data <= 16'h0081; 
        10'b0010111110: data <= 16'h0078; 
        10'b0010111111: data <= 16'h0065; 
        10'b0011000000: data <= 16'h001a; 
        10'b0011000001: data <= 16'hffeb; 
        10'b0011000010: data <= 16'h0002; 
        10'b0011000011: data <= 16'h0026; 
        10'b0011000100: data <= 16'h001f; 
        10'b0011000101: data <= 16'h0011; 
        10'b0011000110: data <= 16'h0015; 
        10'b0011000111: data <= 16'h0005; 
        10'b0011001000: data <= 16'h0033; 
        10'b0011001001: data <= 16'hfff5; 
        10'b0011001010: data <= 16'hffb5; 
        10'b0011001011: data <= 16'hff66; 
        10'b0011001100: data <= 16'hff0f; 
        10'b0011001101: data <= 16'hfece; 
        10'b0011001110: data <= 16'hff30; 
        10'b0011001111: data <= 16'hffa5; 
        10'b0011010000: data <= 16'hffad; 
        10'b0011010001: data <= 16'hff88; 
        10'b0011010010: data <= 16'hff6c; 
        10'b0011010011: data <= 16'hff1a; 
        10'b0011010100: data <= 16'hff37; 
        10'b0011010101: data <= 16'hff43; 
        10'b0011010110: data <= 16'hff56; 
        10'b0011010111: data <= 16'hfffa; 
        10'b0011011000: data <= 16'h0024; 
        10'b0011011001: data <= 16'h0016; 
        10'b0011011010: data <= 16'h0015; 
        10'b0011011011: data <= 16'hffbf; 
        10'b0011011100: data <= 16'hffa8; 
        10'b0011011101: data <= 16'hffdd; 
        10'b0011011110: data <= 16'h001d; 
        10'b0011011111: data <= 16'h0021; 
        10'b0011100000: data <= 16'h0025; 
        10'b0011100001: data <= 16'h001f; 
        10'b0011100010: data <= 16'h001f; 
        10'b0011100011: data <= 16'h0041; 
        10'b0011100100: data <= 16'h0015; 
        10'b0011100101: data <= 16'hfffe; 
        10'b0011100110: data <= 16'hffa7; 
        10'b0011100111: data <= 16'hff78; 
        10'b0011101000: data <= 16'hfee8; 
        10'b0011101001: data <= 16'hfed0; 
        10'b0011101010: data <= 16'hfede; 
        10'b0011101011: data <= 16'hff64; 
        10'b0011101100: data <= 16'hffb8; 
        10'b0011101101: data <= 16'hffa8; 
        10'b0011101110: data <= 16'hffb8; 
        10'b0011101111: data <= 16'h001f; 
        10'b0011110000: data <= 16'hff81; 
        10'b0011110001: data <= 16'hffd5; 
        10'b0011110010: data <= 16'hfff9; 
        10'b0011110011: data <= 16'h0011; 
        10'b0011110100: data <= 16'hffa0; 
        10'b0011110101: data <= 16'hffa3; 
        10'b0011110110: data <= 16'hff6c; 
        10'b0011110111: data <= 16'hff3d; 
        10'b0011111000: data <= 16'hff65; 
        10'b0011111001: data <= 16'hffda; 
        10'b0011111010: data <= 16'h003a; 
        10'b0011111011: data <= 16'h004c; 
        10'b0011111100: data <= 16'h004d; 
        10'b0011111101: data <= 16'h0012; 
        10'b0011111110: data <= 16'h001f; 
        10'b0011111111: data <= 16'h001b; 
        10'b0100000000: data <= 16'hfffb; 
        10'b0100000001: data <= 16'hfff8; 
        10'b0100000010: data <= 16'hff8e; 
        10'b0100000011: data <= 16'hff94; 
        10'b0100000100: data <= 16'hff3f; 
        10'b0100000101: data <= 16'hfeda; 
        10'b0100000110: data <= 16'hfef3; 
        10'b0100000111: data <= 16'hff96; 
        10'b0100001000: data <= 16'hffb0; 
        10'b0100001001: data <= 16'h003c; 
        10'b0100001010: data <= 16'h00be; 
        10'b0100001011: data <= 16'h0111; 
        10'b0100001100: data <= 16'h0065; 
        10'b0100001101: data <= 16'hfff9; 
        10'b0100001110: data <= 16'hffd2; 
        10'b0100001111: data <= 16'hff47; 
        10'b0100010000: data <= 16'hff1d; 
        10'b0100010001: data <= 16'hff20; 
        10'b0100010010: data <= 16'hfee5; 
        10'b0100010011: data <= 16'hff0b; 
        10'b0100010100: data <= 16'hff7d; 
        10'b0100010101: data <= 16'h000f; 
        10'b0100010110: data <= 16'h003f; 
        10'b0100010111: data <= 16'h002e; 
        10'b0100011000: data <= 16'h0046; 
        10'b0100011001: data <= 16'h004d; 
        10'b0100011010: data <= 16'h0040; 
        10'b0100011011: data <= 16'h0008; 
        10'b0100011100: data <= 16'h0034; 
        10'b0100011101: data <= 16'hffc3; 
        10'b0100011110: data <= 16'hff94; 
        10'b0100011111: data <= 16'hffce; 
        10'b0100100000: data <= 16'hff6a; 
        10'b0100100001: data <= 16'hff68; 
        10'b0100100010: data <= 16'hff91; 
        10'b0100100011: data <= 16'hffb6; 
        10'b0100100100: data <= 16'hffce; 
        10'b0100100101: data <= 16'h0098; 
        10'b0100100110: data <= 16'h01ec; 
        10'b0100100111: data <= 16'h0207; 
        10'b0100101000: data <= 16'h00f7; 
        10'b0100101001: data <= 16'hfffb; 
        10'b0100101010: data <= 16'hff6c; 
        10'b0100101011: data <= 16'hff4e; 
        10'b0100101100: data <= 16'hff29; 
        10'b0100101101: data <= 16'hff3e; 
        10'b0100101110: data <= 16'hff49; 
        10'b0100101111: data <= 16'hff8e; 
        10'b0100110000: data <= 16'hffda; 
        10'b0100110001: data <= 16'hfff9; 
        10'b0100110010: data <= 16'h0042; 
        10'b0100110011: data <= 16'h001b; 
        10'b0100110100: data <= 16'h000d; 
        10'b0100110101: data <= 16'h000c; 
        10'b0100110110: data <= 16'h0035; 
        10'b0100110111: data <= 16'h0039; 
        10'b0100111000: data <= 16'h0000; 
        10'b0100111001: data <= 16'hffef; 
        10'b0100111010: data <= 16'hfff7; 
        10'b0100111011: data <= 16'hffa2; 
        10'b0100111100: data <= 16'hffc4; 
        10'b0100111101: data <= 16'hffa3; 
        10'b0100111110: data <= 16'hff77; 
        10'b0100111111: data <= 16'hff30; 
        10'b0101000000: data <= 16'hffe8; 
        10'b0101000001: data <= 16'h0104; 
        10'b0101000010: data <= 16'h0251; 
        10'b0101000011: data <= 16'h0274; 
        10'b0101000100: data <= 16'h00e9; 
        10'b0101000101: data <= 16'hffcd; 
        10'b0101000110: data <= 16'hffd1; 
        10'b0101000111: data <= 16'hff84; 
        10'b0101001000: data <= 16'hff7d; 
        10'b0101001001: data <= 16'hff86; 
        10'b0101001010: data <= 16'hff8f; 
        10'b0101001011: data <= 16'hffcb; 
        10'b0101001100: data <= 16'hffea; 
        10'b0101001101: data <= 16'h0034; 
        10'b0101001110: data <= 16'h0049; 
        10'b0101001111: data <= 16'h0033; 
        10'b0101010000: data <= 16'h0008; 
        10'b0101010001: data <= 16'h0046; 
        10'b0101010010: data <= 16'h0022; 
        10'b0101010011: data <= 16'h0017; 
        10'b0101010100: data <= 16'h0048; 
        10'b0101010101: data <= 16'hfff2; 
        10'b0101010110: data <= 16'hffea; 
        10'b0101010111: data <= 16'hffe1; 
        10'b0101011000: data <= 16'hffa7; 
        10'b0101011001: data <= 16'hff8b; 
        10'b0101011010: data <= 16'hff08; 
        10'b0101011011: data <= 16'hfea5; 
        10'b0101011100: data <= 16'hfff5; 
        10'b0101011101: data <= 16'h0108; 
        10'b0101011110: data <= 16'h02ba; 
        10'b0101011111: data <= 16'h01e4; 
        10'b0101100000: data <= 16'h0060; 
        10'b0101100001: data <= 16'h0033; 
        10'b0101100010: data <= 16'hffe2; 
        10'b0101100011: data <= 16'hff73; 
        10'b0101100100: data <= 16'hffa7; 
        10'b0101100101: data <= 16'hffd5; 
        10'b0101100110: data <= 16'hffe8; 
        10'b0101100111: data <= 16'hffe2; 
        10'b0101101000: data <= 16'h0005; 
        10'b0101101001: data <= 16'h0047; 
        10'b0101101010: data <= 16'h000b; 
        10'b0101101011: data <= 16'h0032; 
        10'b0101101100: data <= 16'h0007; 
        10'b0101101101: data <= 16'h0030; 
        10'b0101101110: data <= 16'h002c; 
        10'b0101101111: data <= 16'h002f; 
        10'b0101110000: data <= 16'h004f; 
        10'b0101110001: data <= 16'h0000; 
        10'b0101110010: data <= 16'h0007; 
        10'b0101110011: data <= 16'hffdd; 
        10'b0101110100: data <= 16'hffd0; 
        10'b0101110101: data <= 16'hff3d; 
        10'b0101110110: data <= 16'hfe63; 
        10'b0101110111: data <= 16'hfe5d; 
        10'b0101111000: data <= 16'h0001; 
        10'b0101111001: data <= 16'h00dc; 
        10'b0101111010: data <= 16'h023f; 
        10'b0101111011: data <= 16'h0145; 
        10'b0101111100: data <= 16'h0056; 
        10'b0101111101: data <= 16'h002a; 
        10'b0101111110: data <= 16'hff7d; 
        10'b0101111111: data <= 16'hff41; 
        10'b0110000000: data <= 16'hffbb; 
        10'b0110000001: data <= 16'hffe8; 
        10'b0110000010: data <= 16'hffe7; 
        10'b0110000011: data <= 16'hfff7; 
        10'b0110000100: data <= 16'h0020; 
        10'b0110000101: data <= 16'h0030; 
        10'b0110000110: data <= 16'h0045; 
        10'b0110000111: data <= 16'h002d; 
        10'b0110001000: data <= 16'h0023; 
        10'b0110001001: data <= 16'h004b; 
        10'b0110001010: data <= 16'h002a; 
        10'b0110001011: data <= 16'h003c; 
        10'b0110001100: data <= 16'h003c; 
        10'b0110001101: data <= 16'h0000; 
        10'b0110001110: data <= 16'h000a; 
        10'b0110001111: data <= 16'hffe9; 
        10'b0110010000: data <= 16'hff7f; 
        10'b0110010001: data <= 16'hff23; 
        10'b0110010010: data <= 16'hfe64; 
        10'b0110010011: data <= 16'hfec8; 
        10'b0110010100: data <= 16'hfff9; 
        10'b0110010101: data <= 16'h00df; 
        10'b0110010110: data <= 16'h01eb; 
        10'b0110010111: data <= 16'h013c; 
        10'b0110011000: data <= 16'h005e; 
        10'b0110011001: data <= 16'hff51; 
        10'b0110011010: data <= 16'hff12; 
        10'b0110011011: data <= 16'hff4c; 
        10'b0110011100: data <= 16'hff95; 
        10'b0110011101: data <= 16'hffe1; 
        10'b0110011110: data <= 16'hffde; 
        10'b0110011111: data <= 16'hffe9; 
        10'b0110100000: data <= 16'h0035; 
        10'b0110100001: data <= 16'h0008; 
        10'b0110100010: data <= 16'h000f; 
        10'b0110100011: data <= 16'h002b; 
        10'b0110100100: data <= 16'h004f; 
        10'b0110100101: data <= 16'h000d; 
        10'b0110100110: data <= 16'h0033; 
        10'b0110100111: data <= 16'h0020; 
        10'b0110101000: data <= 16'h0012; 
        10'b0110101001: data <= 16'h002e; 
        10'b0110101010: data <= 16'hffd3; 
        10'b0110101011: data <= 16'hffcd; 
        10'b0110101100: data <= 16'hffaf; 
        10'b0110101101: data <= 16'hff0e; 
        10'b0110101110: data <= 16'hfef1; 
        10'b0110101111: data <= 16'hffbc; 
        10'b0110110000: data <= 16'h0064; 
        10'b0110110001: data <= 16'h013a; 
        10'b0110110010: data <= 16'h020d; 
        10'b0110110011: data <= 16'h00ba; 
        10'b0110110100: data <= 16'h0022; 
        10'b0110110101: data <= 16'hfeb5; 
        10'b0110110110: data <= 16'hfedb; 
        10'b0110110111: data <= 16'hff4d; 
        10'b0110111000: data <= 16'hff94; 
        10'b0110111001: data <= 16'hffb3; 
        10'b0110111010: data <= 16'hffec; 
        10'b0110111011: data <= 16'h0006; 
        10'b0110111100: data <= 16'h001c; 
        10'b0110111101: data <= 16'h0024; 
        10'b0110111110: data <= 16'h004a; 
        10'b0110111111: data <= 16'h000c; 
        10'b0111000000: data <= 16'h004d; 
        10'b0111000001: data <= 16'h0026; 
        10'b0111000010: data <= 16'h0046; 
        10'b0111000011: data <= 16'h002b; 
        10'b0111000100: data <= 16'h0017; 
        10'b0111000101: data <= 16'hffe1; 
        10'b0111000110: data <= 16'hffb9; 
        10'b0111000111: data <= 16'hffb3; 
        10'b0111001000: data <= 16'hff45; 
        10'b0111001001: data <= 16'hff90; 
        10'b0111001010: data <= 16'hffa7; 
        10'b0111001011: data <= 16'hffce; 
        10'b0111001100: data <= 16'hfff3; 
        10'b0111001101: data <= 16'h019d; 
        10'b0111001110: data <= 16'h01f0; 
        10'b0111001111: data <= 16'h001c; 
        10'b0111010000: data <= 16'hff67; 
        10'b0111010001: data <= 16'hfe9a; 
        10'b0111010010: data <= 16'hfed8; 
        10'b0111010011: data <= 16'hff42; 
        10'b0111010100: data <= 16'hff6f; 
        10'b0111010101: data <= 16'hffc2; 
        10'b0111010110: data <= 16'hffc1; 
        10'b0111010111: data <= 16'h0001; 
        10'b0111011000: data <= 16'hffe4; 
        10'b0111011001: data <= 16'h0004; 
        10'b0111011010: data <= 16'h0013; 
        10'b0111011011: data <= 16'h0028; 
        10'b0111011100: data <= 16'h0020; 
        10'b0111011101: data <= 16'h004c; 
        10'b0111011110: data <= 16'h0011; 
        10'b0111011111: data <= 16'h004b; 
        10'b0111100000: data <= 16'h0037; 
        10'b0111100001: data <= 16'hffd4; 
        10'b0111100010: data <= 16'hff63; 
        10'b0111100011: data <= 16'hff56; 
        10'b0111100100: data <= 16'hff86; 
        10'b0111100101: data <= 16'hffb2; 
        10'b0111100110: data <= 16'h0038; 
        10'b0111100111: data <= 16'h0001; 
        10'b0111101000: data <= 16'h0087; 
        10'b0111101001: data <= 16'h01d9; 
        10'b0111101010: data <= 16'h0196; 
        10'b0111101011: data <= 16'hffae; 
        10'b0111101100: data <= 16'hfee6; 
        10'b0111101101: data <= 16'hfe99; 
        10'b0111101110: data <= 16'hfeda; 
        10'b0111101111: data <= 16'hff46; 
        10'b0111110000: data <= 16'hffba; 
        10'b0111110001: data <= 16'hffdd; 
        10'b0111110010: data <= 16'hffe7; 
        10'b0111110011: data <= 16'hffde; 
        10'b0111110100: data <= 16'hffc6; 
        10'b0111110101: data <= 16'h0011; 
        10'b0111110110: data <= 16'h002c; 
        10'b0111110111: data <= 16'h0034; 
        10'b0111111000: data <= 16'h002f; 
        10'b0111111001: data <= 16'h002b; 
        10'b0111111010: data <= 16'h001b; 
        10'b0111111011: data <= 16'h003f; 
        10'b0111111100: data <= 16'h0023; 
        10'b0111111101: data <= 16'hffc2; 
        10'b0111111110: data <= 16'hff59; 
        10'b0111111111: data <= 16'hff5a; 
        10'b1000000000: data <= 16'hffc2; 
        10'b1000000001: data <= 16'h0040; 
        10'b1000000010: data <= 16'h0035; 
        10'b1000000011: data <= 16'h0054; 
        10'b1000000100: data <= 16'h00dc; 
        10'b1000000101: data <= 16'h0161; 
        10'b1000000110: data <= 16'h00f4; 
        10'b1000000111: data <= 16'hff5f; 
        10'b1000001000: data <= 16'hfef8; 
        10'b1000001001: data <= 16'hff1e; 
        10'b1000001010: data <= 16'hff3f; 
        10'b1000001011: data <= 16'hff7f; 
        10'b1000001100: data <= 16'hffc0; 
        10'b1000001101: data <= 16'hff94; 
        10'b1000001110: data <= 16'hffd0; 
        10'b1000001111: data <= 16'hffb7; 
        10'b1000010000: data <= 16'hffd3; 
        10'b1000010001: data <= 16'h0029; 
        10'b1000010010: data <= 16'h0046; 
        10'b1000010011: data <= 16'h0048; 
        10'b1000010100: data <= 16'h004a; 
        10'b1000010101: data <= 16'h0034; 
        10'b1000010110: data <= 16'h0036; 
        10'b1000010111: data <= 16'h003c; 
        10'b1000011000: data <= 16'h0007; 
        10'b1000011001: data <= 16'hffa3; 
        10'b1000011010: data <= 16'hff30; 
        10'b1000011011: data <= 16'hff74; 
        10'b1000011100: data <= 16'hffc7; 
        10'b1000011101: data <= 16'h0021; 
        10'b1000011110: data <= 16'h0011; 
        10'b1000011111: data <= 16'h000b; 
        10'b1000100000: data <= 16'h001d; 
        10'b1000100001: data <= 16'h00a3; 
        10'b1000100010: data <= 16'h0024; 
        10'b1000100011: data <= 16'hff7b; 
        10'b1000100100: data <= 16'hff91; 
        10'b1000100101: data <= 16'hffa0; 
        10'b1000100110: data <= 16'hff87; 
        10'b1000100111: data <= 16'hffa2; 
        10'b1000101000: data <= 16'hff77; 
        10'b1000101001: data <= 16'hff8e; 
        10'b1000101010: data <= 16'hffbb; 
        10'b1000101011: data <= 16'hffc3; 
        10'b1000101100: data <= 16'h0003; 
        10'b1000101101: data <= 16'h0017; 
        10'b1000101110: data <= 16'h001a; 
        10'b1000101111: data <= 16'h000a; 
        10'b1000110000: data <= 16'h000c; 
        10'b1000110001: data <= 16'h004e; 
        10'b1000110010: data <= 16'h002a; 
        10'b1000110011: data <= 16'h001b; 
        10'b1000110100: data <= 16'hffeb; 
        10'b1000110101: data <= 16'hffbe; 
        10'b1000110110: data <= 16'hfff4; 
        10'b1000110111: data <= 16'hffd2; 
        10'b1000111000: data <= 16'hffff; 
        10'b1000111001: data <= 16'h0013; 
        10'b1000111010: data <= 16'hffcd; 
        10'b1000111011: data <= 16'hffee; 
        10'b1000111100: data <= 16'hffad; 
        10'b1000111101: data <= 16'hffe4; 
        10'b1000111110: data <= 16'hffeb; 
        10'b1000111111: data <= 16'h0005; 
        10'b1001000000: data <= 16'h004f; 
        10'b1001000001: data <= 16'h001c; 
        10'b1001000010: data <= 16'hffe2; 
        10'b1001000011: data <= 16'hff91; 
        10'b1001000100: data <= 16'hff77; 
        10'b1001000101: data <= 16'hff82; 
        10'b1001000110: data <= 16'hff9d; 
        10'b1001000111: data <= 16'hffea; 
        10'b1001001000: data <= 16'h000a; 
        10'b1001001001: data <= 16'h003f; 
        10'b1001001010: data <= 16'h0019; 
        10'b1001001011: data <= 16'h004e; 
        10'b1001001100: data <= 16'h0037; 
        10'b1001001101: data <= 16'h001d; 
        10'b1001001110: data <= 16'h002d; 
        10'b1001001111: data <= 16'h0036; 
        10'b1001010000: data <= 16'h002b; 
        10'b1001010001: data <= 16'h0074; 
        10'b1001010010: data <= 16'h0060; 
        10'b1001010011: data <= 16'h002d; 
        10'b1001010100: data <= 16'h0008; 
        10'b1001010101: data <= 16'hffdf; 
        10'b1001010110: data <= 16'h0001; 
        10'b1001010111: data <= 16'hffbd; 
        10'b1001011000: data <= 16'hff67; 
        10'b1001011001: data <= 16'hff52; 
        10'b1001011010: data <= 16'hfff0; 
        10'b1001011011: data <= 16'h0034; 
        10'b1001011100: data <= 16'h0054; 
        10'b1001011101: data <= 16'h005f; 
        10'b1001011110: data <= 16'h0042; 
        10'b1001011111: data <= 16'hff91; 
        10'b1001100000: data <= 16'hff93; 
        10'b1001100001: data <= 16'hff84; 
        10'b1001100010: data <= 16'hffab; 
        10'b1001100011: data <= 16'hffcf; 
        10'b1001100100: data <= 16'h000b; 
        10'b1001100101: data <= 16'h0022; 
        10'b1001100110: data <= 16'h0007; 
        10'b1001100111: data <= 16'h000a; 
        10'b1001101000: data <= 16'h002b; 
        10'b1001101001: data <= 16'h002c; 
        10'b1001101010: data <= 16'h0032; 
        10'b1001101011: data <= 16'h000a; 
        10'b1001101100: data <= 16'h0065; 
        10'b1001101101: data <= 16'h00e1; 
        10'b1001101110: data <= 16'h00e9; 
        10'b1001101111: data <= 16'h008d; 
        10'b1001110000: data <= 16'h0013; 
        10'b1001110001: data <= 16'hfff0; 
        10'b1001110010: data <= 16'hffcb; 
        10'b1001110011: data <= 16'hff22; 
        10'b1001110100: data <= 16'hfe97; 
        10'b1001110101: data <= 16'hfeec; 
        10'b1001110110: data <= 16'h0001; 
        10'b1001110111: data <= 16'h0036; 
        10'b1001111000: data <= 16'h00cf; 
        10'b1001111001: data <= 16'h0153; 
        10'b1001111010: data <= 16'h0094; 
        10'b1001111011: data <= 16'h001f; 
        10'b1001111100: data <= 16'hffb4; 
        10'b1001111101: data <= 16'hffc5; 
        10'b1001111110: data <= 16'hfffb; 
        10'b1001111111: data <= 16'h000a; 
        10'b1010000000: data <= 16'h0005; 
        10'b1010000001: data <= 16'h0021; 
        10'b1010000010: data <= 16'h004b; 
        10'b1010000011: data <= 16'h0024; 
        10'b1010000100: data <= 16'h0046; 
        10'b1010000101: data <= 16'h002c; 
        10'b1010000110: data <= 16'h0038; 
        10'b1010000111: data <= 16'h001f; 
        10'b1010001000: data <= 16'h005a; 
        10'b1010001001: data <= 16'h00c2; 
        10'b1010001010: data <= 16'h00ce; 
        10'b1010001011: data <= 16'h005f; 
        10'b1010001100: data <= 16'h001a; 
        10'b1010001101: data <= 16'hffd0; 
        10'b1010001110: data <= 16'hffdf; 
        10'b1010001111: data <= 16'hff82; 
        10'b1010010000: data <= 16'hffa8; 
        10'b1010010001: data <= 16'hffb2; 
        10'b1010010010: data <= 16'hff97; 
        10'b1010010011: data <= 16'h0029; 
        10'b1010010100: data <= 16'h00f1; 
        10'b1010010101: data <= 16'h0122; 
        10'b1010010110: data <= 16'h0082; 
        10'b1010010111: data <= 16'hffe9; 
        10'b1010011000: data <= 16'hffc9; 
        10'b1010011001: data <= 16'hffaa; 
        10'b1010011010: data <= 16'hffe2; 
        10'b1010011011: data <= 16'hffe5; 
        10'b1010011100: data <= 16'h0011; 
        10'b1010011101: data <= 16'h0009; 
        10'b1010011110: data <= 16'h0010; 
        10'b1010011111: data <= 16'h0008; 
        10'b1010100000: data <= 16'h0011; 
        10'b1010100001: data <= 16'h000b; 
        10'b1010100010: data <= 16'h001c; 
        10'b1010100011: data <= 16'h0009; 
        10'b1010100100: data <= 16'h002c; 
        10'b1010100101: data <= 16'h0056; 
        10'b1010100110: data <= 16'h0058; 
        10'b1010100111: data <= 16'hffe3; 
        10'b1010101000: data <= 16'hff80; 
        10'b1010101001: data <= 16'hff7f; 
        10'b1010101010: data <= 16'hff1d; 
        10'b1010101011: data <= 16'hff27; 
        10'b1010101100: data <= 16'hff3d; 
        10'b1010101101: data <= 16'hff59; 
        10'b1010101110: data <= 16'hff5a; 
        10'b1010101111: data <= 16'hff5a; 
        10'b1010110000: data <= 16'hffd0; 
        10'b1010110001: data <= 16'h0014; 
        10'b1010110010: data <= 16'h0025; 
        10'b1010110011: data <= 16'h0035; 
        10'b1010110100: data <= 16'h002d; 
        10'b1010110101: data <= 16'h000b; 
        10'b1010110110: data <= 16'h0017; 
        10'b1010110111: data <= 16'h003e; 
        10'b1010111000: data <= 16'h0013; 
        10'b1010111001: data <= 16'h001e; 
        10'b1010111010: data <= 16'h003b; 
        10'b1010111011: data <= 16'h0013; 
        10'b1010111100: data <= 16'h004c; 
        10'b1010111101: data <= 16'h0018; 
        10'b1010111110: data <= 16'h001d; 
        10'b1010111111: data <= 16'h0029; 
        10'b1011000000: data <= 16'h003b; 
        10'b1011000001: data <= 16'h0035; 
        10'b1011000010: data <= 16'h0001; 
        10'b1011000011: data <= 16'hffdf; 
        10'b1011000100: data <= 16'hfff3; 
        10'b1011000101: data <= 16'hffe2; 
        10'b1011000110: data <= 16'hff81; 
        10'b1011000111: data <= 16'hff66; 
        10'b1011001000: data <= 16'hff8e; 
        10'b1011001001: data <= 16'hff60; 
        10'b1011001010: data <= 16'hff9e; 
        10'b1011001011: data <= 16'hff84; 
        10'b1011001100: data <= 16'hffb9; 
        10'b1011001101: data <= 16'hfff3; 
        10'b1011001110: data <= 16'h0019; 
        10'b1011001111: data <= 16'h0033; 
        10'b1011010000: data <= 16'h0005; 
        10'b1011010001: data <= 16'h002e; 
        10'b1011010010: data <= 16'h001c; 
        10'b1011010011: data <= 16'h0042; 
        10'b1011010100: data <= 16'h0011; 
        10'b1011010101: data <= 16'h0014; 
        10'b1011010110: data <= 16'h001c; 
        10'b1011010111: data <= 16'h0018; 
        10'b1011011000: data <= 16'h001c; 
        10'b1011011001: data <= 16'h0036; 
        10'b1011011010: data <= 16'h0030; 
        10'b1011011011: data <= 16'h000f; 
        10'b1011011100: data <= 16'h0034; 
        10'b1011011101: data <= 16'h0045; 
        10'b1011011110: data <= 16'h002f; 
        10'b1011011111: data <= 16'h002b; 
        10'b1011100000: data <= 16'h003d; 
        10'b1011100001: data <= 16'h0034; 
        10'b1011100010: data <= 16'h0007; 
        10'b1011100011: data <= 16'h002a; 
        10'b1011100100: data <= 16'h0026; 
        10'b1011100101: data <= 16'h0016; 
        10'b1011100110: data <= 16'hffff; 
        10'b1011100111: data <= 16'h0014; 
        10'b1011101000: data <= 16'h002d; 
        10'b1011101001: data <= 16'h0046; 
        10'b1011101010: data <= 16'h0033; 
        10'b1011101011: data <= 16'h0008; 
        10'b1011101100: data <= 16'h0030; 
        10'b1011101101: data <= 16'h002d; 
        10'b1011101110: data <= 16'h002b; 
        10'b1011101111: data <= 16'h0014; 
        10'b1011110000: data <= 16'h0012; 
        10'b1011110001: data <= 16'h0034; 
        10'b1011110010: data <= 16'h0047; 
        10'b1011110011: data <= 16'h003a; 
        10'b1011110100: data <= 16'h003a; 
        10'b1011110101: data <= 16'h0049; 
        10'b1011110110: data <= 16'h000c; 
        10'b1011110111: data <= 16'h0028; 
        10'b1011111000: data <= 16'h004d; 
        10'b1011111001: data <= 16'h003d; 
        10'b1011111010: data <= 16'h0045; 
        10'b1011111011: data <= 16'h0040; 
        10'b1011111100: data <= 16'h0045; 
        10'b1011111101: data <= 16'h0021; 
        10'b1011111110: data <= 16'h003d; 
        10'b1011111111: data <= 16'h003f; 
        10'b1100000000: data <= 16'h0006; 
        10'b1100000001: data <= 16'h000d; 
        10'b1100000010: data <= 16'h004b; 
        10'b1100000011: data <= 16'h0031; 
        10'b1100000100: data <= 16'h002d; 
        10'b1100000101: data <= 16'h0007; 
        10'b1100000110: data <= 16'h0021; 
        10'b1100000111: data <= 16'h000e; 
        10'b1100001000: data <= 16'h000d; 
        10'b1100001001: data <= 16'h0019; 
        10'b1100001010: data <= 16'h002c; 
        10'b1100001011: data <= 16'h0040; 
        10'b1100001100: data <= 16'h0047; 
        10'b1100001101: data <= 16'h0045; 
        10'b1100001110: data <= 16'h0044; 
        10'b1100001111: data <= 16'h0017; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 11) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 17'h00080; 
        10'b0000000001: data <= 17'h0003d; 
        10'b0000000010: data <= 17'h00044; 
        10'b0000000011: data <= 17'h0001c; 
        10'b0000000100: data <= 17'h0006c; 
        10'b0000000101: data <= 17'h00069; 
        10'b0000000110: data <= 17'h00074; 
        10'b0000000111: data <= 17'h0001d; 
        10'b0000001000: data <= 17'h00065; 
        10'b0000001001: data <= 17'h0001f; 
        10'b0000001010: data <= 17'h00060; 
        10'b0000001011: data <= 17'h0004e; 
        10'b0000001100: data <= 17'h0006d; 
        10'b0000001101: data <= 17'h00091; 
        10'b0000001110: data <= 17'h0007f; 
        10'b0000001111: data <= 17'h00057; 
        10'b0000010000: data <= 17'h00059; 
        10'b0000010001: data <= 17'h0001f; 
        10'b0000010010: data <= 17'h00095; 
        10'b0000010011: data <= 17'h00094; 
        10'b0000010100: data <= 17'h00054; 
        10'b0000010101: data <= 17'h0006c; 
        10'b0000010110: data <= 17'h00054; 
        10'b0000010111: data <= 17'h00082; 
        10'b0000011000: data <= 17'h00031; 
        10'b0000011001: data <= 17'h00089; 
        10'b0000011010: data <= 17'h00054; 
        10'b0000011011: data <= 17'h00079; 
        10'b0000011100: data <= 17'h00010; 
        10'b0000011101: data <= 17'h00080; 
        10'b0000011110: data <= 17'h00026; 
        10'b0000011111: data <= 17'h0005b; 
        10'b0000100000: data <= 17'h00052; 
        10'b0000100001: data <= 17'h00020; 
        10'b0000100010: data <= 17'h0002e; 
        10'b0000100011: data <= 17'h00079; 
        10'b0000100100: data <= 17'h00074; 
        10'b0000100101: data <= 17'h0005e; 
        10'b0000100110: data <= 17'h0005d; 
        10'b0000100111: data <= 17'h00045; 
        10'b0000101000: data <= 17'h0006f; 
        10'b0000101001: data <= 17'h0007d; 
        10'b0000101010: data <= 17'h000a2; 
        10'b0000101011: data <= 17'h00050; 
        10'b0000101100: data <= 17'h00041; 
        10'b0000101101: data <= 17'h00082; 
        10'b0000101110: data <= 17'h00057; 
        10'b0000101111: data <= 17'h0003b; 
        10'b0000110000: data <= 17'h0008d; 
        10'b0000110001: data <= 17'h00087; 
        10'b0000110010: data <= 17'h00037; 
        10'b0000110011: data <= 17'h00091; 
        10'b0000110100: data <= 17'h0009b; 
        10'b0000110101: data <= 17'h00052; 
        10'b0000110110: data <= 17'h00084; 
        10'b0000110111: data <= 17'h0006a; 
        10'b0000111000: data <= 17'h00083; 
        10'b0000111001: data <= 17'h00062; 
        10'b0000111010: data <= 17'h0009d; 
        10'b0000111011: data <= 17'h0001e; 
        10'b0000111100: data <= 17'h0001d; 
        10'b0000111101: data <= 17'h00067; 
        10'b0000111110: data <= 17'h0004c; 
        10'b0000111111: data <= 17'h00049; 
        10'b0001000000: data <= 17'h00031; 
        10'b0001000001: data <= 17'h00056; 
        10'b0001000010: data <= 17'h00002; 
        10'b0001000011: data <= 17'h0002b; 
        10'b0001000100: data <= 17'h00006; 
        10'b0001000101: data <= 17'h00026; 
        10'b0001000110: data <= 17'h0004f; 
        10'b0001000111: data <= 17'h00080; 
        10'b0001001000: data <= 17'h00061; 
        10'b0001001001: data <= 17'h00000; 
        10'b0001001010: data <= 17'h0005f; 
        10'b0001001011: data <= 17'h00039; 
        10'b0001001100: data <= 17'h0007d; 
        10'b0001001101: data <= 17'h00036; 
        10'b0001001110: data <= 17'h0008a; 
        10'b0001001111: data <= 17'h00064; 
        10'b0001010000: data <= 17'h0006c; 
        10'b0001010001: data <= 17'h00012; 
        10'b0001010010: data <= 17'h00075; 
        10'b0001010011: data <= 17'h00078; 
        10'b0001010100: data <= 17'h0002f; 
        10'b0001010101: data <= 17'h00034; 
        10'b0001010110: data <= 17'h00058; 
        10'b0001010111: data <= 17'h00048; 
        10'b0001011000: data <= 17'h00093; 
        10'b0001011001: data <= 17'h0004d; 
        10'b0001011010: data <= 17'h00011; 
        10'b0001011011: data <= 17'h00090; 
        10'b0001011100: data <= 17'h1fff0; 
        10'b0001011101: data <= 17'h1ffe3; 
        10'b0001011110: data <= 17'h1ffe4; 
        10'b0001011111: data <= 17'h1ffb0; 
        10'b0001100000: data <= 17'h1ffe4; 
        10'b0001100001: data <= 17'h0000b; 
        10'b0001100010: data <= 17'h0003c; 
        10'b0001100011: data <= 17'h00078; 
        10'b0001100100: data <= 17'h1ffc5; 
        10'b0001100101: data <= 17'h1ffea; 
        10'b0001100110: data <= 17'h1fffd; 
        10'b0001100111: data <= 17'h1ffa4; 
        10'b0001101000: data <= 17'h1fff6; 
        10'b0001101001: data <= 17'h00026; 
        10'b0001101010: data <= 17'h00060; 
        10'b0001101011: data <= 17'h0005e; 
        10'b0001101100: data <= 17'h1ffef; 
        10'b0001101101: data <= 17'h00085; 
        10'b0001101110: data <= 17'h00032; 
        10'b0001101111: data <= 17'h0008c; 
        10'b0001110000: data <= 17'h0006c; 
        10'b0001110001: data <= 17'h00041; 
        10'b0001110010: data <= 17'h00095; 
        10'b0001110011: data <= 17'h00093; 
        10'b0001110100: data <= 17'h00010; 
        10'b0001110101: data <= 17'h0001d; 
        10'b0001110110: data <= 17'h00082; 
        10'b0001110111: data <= 17'h00053; 
        10'b0001111000: data <= 17'h0001f; 
        10'b0001111001: data <= 17'h1ff78; 
        10'b0001111010: data <= 17'h0000c; 
        10'b0001111011: data <= 17'h00030; 
        10'b0001111100: data <= 17'h0004a; 
        10'b0001111101: data <= 17'h00084; 
        10'b0001111110: data <= 17'h0009b; 
        10'b0001111111: data <= 17'h0013d; 
        10'b0010000000: data <= 17'h00057; 
        10'b0010000001: data <= 17'h1ffbd; 
        10'b0010000010: data <= 17'h1ffb7; 
        10'b0010000011: data <= 17'h00031; 
        10'b0010000100: data <= 17'h000af; 
        10'b0010000101: data <= 17'h000c4; 
        10'b0010000110: data <= 17'h000c3; 
        10'b0010000111: data <= 17'h000e5; 
        10'b0010001000: data <= 17'h00078; 
        10'b0010001001: data <= 17'h00039; 
        10'b0010001010: data <= 17'h00032; 
        10'b0010001011: data <= 17'h00037; 
        10'b0010001100: data <= 17'h00014; 
        10'b0010001101: data <= 17'h00080; 
        10'b0010001110: data <= 17'h00019; 
        10'b0010001111: data <= 17'h0005a; 
        10'b0010010000: data <= 17'h00017; 
        10'b0010010001: data <= 17'h00056; 
        10'b0010010010: data <= 17'h0001a; 
        10'b0010010011: data <= 17'h1ffdf; 
        10'b0010010100: data <= 17'h1fee3; 
        10'b0010010101: data <= 17'h1fee0; 
        10'b0010010110: data <= 17'h1ff7c; 
        10'b0010010111: data <= 17'h00002; 
        10'b0010011000: data <= 17'h0006c; 
        10'b0010011001: data <= 17'h0007a; 
        10'b0010011010: data <= 17'h000d3; 
        10'b0010011011: data <= 17'h000a4; 
        10'b0010011100: data <= 17'h00061; 
        10'b0010011101: data <= 17'h1ff60; 
        10'b0010011110: data <= 17'h1fff0; 
        10'b0010011111: data <= 17'h00021; 
        10'b0010100000: data <= 17'h0009c; 
        10'b0010100001: data <= 17'h000fb; 
        10'b0010100010: data <= 17'h001a2; 
        10'b0010100011: data <= 17'h00105; 
        10'b0010100100: data <= 17'h000d6; 
        10'b0010100101: data <= 17'h1ffc9; 
        10'b0010100110: data <= 17'h0003b; 
        10'b0010100111: data <= 17'h00021; 
        10'b0010101000: data <= 17'h0001b; 
        10'b0010101001: data <= 17'h0005d; 
        10'b0010101010: data <= 17'h00011; 
        10'b0010101011: data <= 17'h00048; 
        10'b0010101100: data <= 17'h00011; 
        10'b0010101101: data <= 17'h1ffd5; 
        10'b0010101110: data <= 17'h1ff63; 
        10'b0010101111: data <= 17'h1ff65; 
        10'b0010110000: data <= 17'h1fe9b; 
        10'b0010110001: data <= 17'h1fe51; 
        10'b0010110010: data <= 17'h1fef2; 
        10'b0010110011: data <= 17'h1ffc1; 
        10'b0010110100: data <= 17'h1ffbe; 
        10'b0010110101: data <= 17'h1ff79; 
        10'b0010110110: data <= 17'h1ffc2; 
        10'b0010110111: data <= 17'h1fecb; 
        10'b0010111000: data <= 17'h1feb3; 
        10'b0010111001: data <= 17'h1feb1; 
        10'b0010111010: data <= 17'h1ff74; 
        10'b0010111011: data <= 17'h1ff98; 
        10'b0010111100: data <= 17'h0009d; 
        10'b0010111101: data <= 17'h00102; 
        10'b0010111110: data <= 17'h000ef; 
        10'b0010111111: data <= 17'h000ca; 
        10'b0011000000: data <= 17'h00034; 
        10'b0011000001: data <= 17'h1ffd5; 
        10'b0011000010: data <= 17'h00004; 
        10'b0011000011: data <= 17'h0004c; 
        10'b0011000100: data <= 17'h0003d; 
        10'b0011000101: data <= 17'h00022; 
        10'b0011000110: data <= 17'h0002b; 
        10'b0011000111: data <= 17'h0000a; 
        10'b0011001000: data <= 17'h00065; 
        10'b0011001001: data <= 17'h1ffea; 
        10'b0011001010: data <= 17'h1ff6a; 
        10'b0011001011: data <= 17'h1fecc; 
        10'b0011001100: data <= 17'h1fe1f; 
        10'b0011001101: data <= 17'h1fd9b; 
        10'b0011001110: data <= 17'h1fe60; 
        10'b0011001111: data <= 17'h1ff4a; 
        10'b0011010000: data <= 17'h1ff5a; 
        10'b0011010001: data <= 17'h1ff11; 
        10'b0011010010: data <= 17'h1fed8; 
        10'b0011010011: data <= 17'h1fe34; 
        10'b0011010100: data <= 17'h1fe6e; 
        10'b0011010101: data <= 17'h1fe87; 
        10'b0011010110: data <= 17'h1feac; 
        10'b0011010111: data <= 17'h1fff4; 
        10'b0011011000: data <= 17'h00047; 
        10'b0011011001: data <= 17'h0002c; 
        10'b0011011010: data <= 17'h0002a; 
        10'b0011011011: data <= 17'h1ff7f; 
        10'b0011011100: data <= 17'h1ff4f; 
        10'b0011011101: data <= 17'h1ffb9; 
        10'b0011011110: data <= 17'h00039; 
        10'b0011011111: data <= 17'h00043; 
        10'b0011100000: data <= 17'h0004a; 
        10'b0011100001: data <= 17'h0003f; 
        10'b0011100010: data <= 17'h0003e; 
        10'b0011100011: data <= 17'h00083; 
        10'b0011100100: data <= 17'h0002a; 
        10'b0011100101: data <= 17'h1fffc; 
        10'b0011100110: data <= 17'h1ff4d; 
        10'b0011100111: data <= 17'h1fef1; 
        10'b0011101000: data <= 17'h1fdcf; 
        10'b0011101001: data <= 17'h1fd9f; 
        10'b0011101010: data <= 17'h1fdbc; 
        10'b0011101011: data <= 17'h1fec8; 
        10'b0011101100: data <= 17'h1ff71; 
        10'b0011101101: data <= 17'h1ff50; 
        10'b0011101110: data <= 17'h1ff70; 
        10'b0011101111: data <= 17'h0003f; 
        10'b0011110000: data <= 17'h1ff01; 
        10'b0011110001: data <= 17'h1ffaa; 
        10'b0011110010: data <= 17'h1fff2; 
        10'b0011110011: data <= 17'h00021; 
        10'b0011110100: data <= 17'h1ff40; 
        10'b0011110101: data <= 17'h1ff47; 
        10'b0011110110: data <= 17'h1fed7; 
        10'b0011110111: data <= 17'h1fe7a; 
        10'b0011111000: data <= 17'h1feca; 
        10'b0011111001: data <= 17'h1ffb4; 
        10'b0011111010: data <= 17'h00073; 
        10'b0011111011: data <= 17'h00098; 
        10'b0011111100: data <= 17'h0009a; 
        10'b0011111101: data <= 17'h00023; 
        10'b0011111110: data <= 17'h0003f; 
        10'b0011111111: data <= 17'h00036; 
        10'b0100000000: data <= 17'h1fff6; 
        10'b0100000001: data <= 17'h1ffef; 
        10'b0100000010: data <= 17'h1ff1c; 
        10'b0100000011: data <= 17'h1ff28; 
        10'b0100000100: data <= 17'h1fe7e; 
        10'b0100000101: data <= 17'h1fdb4; 
        10'b0100000110: data <= 17'h1fde5; 
        10'b0100000111: data <= 17'h1ff2b; 
        10'b0100001000: data <= 17'h1ff61; 
        10'b0100001001: data <= 17'h00079; 
        10'b0100001010: data <= 17'h0017d; 
        10'b0100001011: data <= 17'h00221; 
        10'b0100001100: data <= 17'h000ca; 
        10'b0100001101: data <= 17'h1fff2; 
        10'b0100001110: data <= 17'h1ffa5; 
        10'b0100001111: data <= 17'h1fe8e; 
        10'b0100010000: data <= 17'h1fe39; 
        10'b0100010001: data <= 17'h1fe3f; 
        10'b0100010010: data <= 17'h1fdcb; 
        10'b0100010011: data <= 17'h1fe16; 
        10'b0100010100: data <= 17'h1fef9; 
        10'b0100010101: data <= 17'h0001f; 
        10'b0100010110: data <= 17'h0007f; 
        10'b0100010111: data <= 17'h0005c; 
        10'b0100011000: data <= 17'h0008c; 
        10'b0100011001: data <= 17'h0009b; 
        10'b0100011010: data <= 17'h00080; 
        10'b0100011011: data <= 17'h00011; 
        10'b0100011100: data <= 17'h00069; 
        10'b0100011101: data <= 17'h1ff87; 
        10'b0100011110: data <= 17'h1ff29; 
        10'b0100011111: data <= 17'h1ff9c; 
        10'b0100100000: data <= 17'h1fed5; 
        10'b0100100001: data <= 17'h1fed0; 
        10'b0100100010: data <= 17'h1ff22; 
        10'b0100100011: data <= 17'h1ff6c; 
        10'b0100100100: data <= 17'h1ff9c; 
        10'b0100100101: data <= 17'h00130; 
        10'b0100100110: data <= 17'h003d8; 
        10'b0100100111: data <= 17'h0040f; 
        10'b0100101000: data <= 17'h001ed; 
        10'b0100101001: data <= 17'h1fff5; 
        10'b0100101010: data <= 17'h1fed9; 
        10'b0100101011: data <= 17'h1fe9c; 
        10'b0100101100: data <= 17'h1fe51; 
        10'b0100101101: data <= 17'h1fe7b; 
        10'b0100101110: data <= 17'h1fe92; 
        10'b0100101111: data <= 17'h1ff1d; 
        10'b0100110000: data <= 17'h1ffb4; 
        10'b0100110001: data <= 17'h1fff3; 
        10'b0100110010: data <= 17'h00084; 
        10'b0100110011: data <= 17'h00036; 
        10'b0100110100: data <= 17'h0001a; 
        10'b0100110101: data <= 17'h00018; 
        10'b0100110110: data <= 17'h0006b; 
        10'b0100110111: data <= 17'h00072; 
        10'b0100111000: data <= 17'h00000; 
        10'b0100111001: data <= 17'h1ffde; 
        10'b0100111010: data <= 17'h1ffee; 
        10'b0100111011: data <= 17'h1ff45; 
        10'b0100111100: data <= 17'h1ff87; 
        10'b0100111101: data <= 17'h1ff45; 
        10'b0100111110: data <= 17'h1feed; 
        10'b0100111111: data <= 17'h1fe61; 
        10'b0101000000: data <= 17'h1ffd0; 
        10'b0101000001: data <= 17'h00208; 
        10'b0101000010: data <= 17'h004a2; 
        10'b0101000011: data <= 17'h004e9; 
        10'b0101000100: data <= 17'h001d2; 
        10'b0101000101: data <= 17'h1ff9a; 
        10'b0101000110: data <= 17'h1ffa2; 
        10'b0101000111: data <= 17'h1ff08; 
        10'b0101001000: data <= 17'h1fefa; 
        10'b0101001001: data <= 17'h1ff0d; 
        10'b0101001010: data <= 17'h1ff1f; 
        10'b0101001011: data <= 17'h1ff97; 
        10'b0101001100: data <= 17'h1ffd3; 
        10'b0101001101: data <= 17'h00068; 
        10'b0101001110: data <= 17'h00092; 
        10'b0101001111: data <= 17'h00067; 
        10'b0101010000: data <= 17'h00010; 
        10'b0101010001: data <= 17'h0008c; 
        10'b0101010010: data <= 17'h00043; 
        10'b0101010011: data <= 17'h0002d; 
        10'b0101010100: data <= 17'h0008f; 
        10'b0101010101: data <= 17'h1ffe5; 
        10'b0101010110: data <= 17'h1ffd4; 
        10'b0101010111: data <= 17'h1ffc2; 
        10'b0101011000: data <= 17'h1ff4e; 
        10'b0101011001: data <= 17'h1ff16; 
        10'b0101011010: data <= 17'h1fe11; 
        10'b0101011011: data <= 17'h1fd49; 
        10'b0101011100: data <= 17'h1ffea; 
        10'b0101011101: data <= 17'h00210; 
        10'b0101011110: data <= 17'h00574; 
        10'b0101011111: data <= 17'h003c8; 
        10'b0101100000: data <= 17'h000c0; 
        10'b0101100001: data <= 17'h00065; 
        10'b0101100010: data <= 17'h1ffc4; 
        10'b0101100011: data <= 17'h1fee5; 
        10'b0101100100: data <= 17'h1ff4d; 
        10'b0101100101: data <= 17'h1ffa9; 
        10'b0101100110: data <= 17'h1ffcf; 
        10'b0101100111: data <= 17'h1ffc4; 
        10'b0101101000: data <= 17'h00009; 
        10'b0101101001: data <= 17'h0008e; 
        10'b0101101010: data <= 17'h00015; 
        10'b0101101011: data <= 17'h00064; 
        10'b0101101100: data <= 17'h0000e; 
        10'b0101101101: data <= 17'h0005f; 
        10'b0101101110: data <= 17'h00059; 
        10'b0101101111: data <= 17'h0005f; 
        10'b0101110000: data <= 17'h0009e; 
        10'b0101110001: data <= 17'h00001; 
        10'b0101110010: data <= 17'h0000d; 
        10'b0101110011: data <= 17'h1ffb9; 
        10'b0101110100: data <= 17'h1ffa1; 
        10'b0101110101: data <= 17'h1fe7a; 
        10'b0101110110: data <= 17'h1fcc6; 
        10'b0101110111: data <= 17'h1fcba; 
        10'b0101111000: data <= 17'h00001; 
        10'b0101111001: data <= 17'h001b8; 
        10'b0101111010: data <= 17'h0047f; 
        10'b0101111011: data <= 17'h0028a; 
        10'b0101111100: data <= 17'h000ac; 
        10'b0101111101: data <= 17'h00053; 
        10'b0101111110: data <= 17'h1fef9; 
        10'b0101111111: data <= 17'h1fe82; 
        10'b0110000000: data <= 17'h1ff75; 
        10'b0110000001: data <= 17'h1ffcf; 
        10'b0110000010: data <= 17'h1ffcd; 
        10'b0110000011: data <= 17'h1ffee; 
        10'b0110000100: data <= 17'h00040; 
        10'b0110000101: data <= 17'h00060; 
        10'b0110000110: data <= 17'h0008b; 
        10'b0110000111: data <= 17'h0005a; 
        10'b0110001000: data <= 17'h00046; 
        10'b0110001001: data <= 17'h00096; 
        10'b0110001010: data <= 17'h00054; 
        10'b0110001011: data <= 17'h00078; 
        10'b0110001100: data <= 17'h00078; 
        10'b0110001101: data <= 17'h00000; 
        10'b0110001110: data <= 17'h00015; 
        10'b0110001111: data <= 17'h1ffd2; 
        10'b0110010000: data <= 17'h1fefe; 
        10'b0110010001: data <= 17'h1fe46; 
        10'b0110010010: data <= 17'h1fcc9; 
        10'b0110010011: data <= 17'h1fd8f; 
        10'b0110010100: data <= 17'h1fff2; 
        10'b0110010101: data <= 17'h001bf; 
        10'b0110010110: data <= 17'h003d5; 
        10'b0110010111: data <= 17'h00278; 
        10'b0110011000: data <= 17'h000bd; 
        10'b0110011001: data <= 17'h1fea1; 
        10'b0110011010: data <= 17'h1fe25; 
        10'b0110011011: data <= 17'h1fe97; 
        10'b0110011100: data <= 17'h1ff2b; 
        10'b0110011101: data <= 17'h1ffc2; 
        10'b0110011110: data <= 17'h1ffbd; 
        10'b0110011111: data <= 17'h1ffd2; 
        10'b0110100000: data <= 17'h0006b; 
        10'b0110100001: data <= 17'h00010; 
        10'b0110100010: data <= 17'h0001e; 
        10'b0110100011: data <= 17'h00055; 
        10'b0110100100: data <= 17'h0009f; 
        10'b0110100101: data <= 17'h0001a; 
        10'b0110100110: data <= 17'h00066; 
        10'b0110100111: data <= 17'h00041; 
        10'b0110101000: data <= 17'h00024; 
        10'b0110101001: data <= 17'h0005c; 
        10'b0110101010: data <= 17'h1ffa6; 
        10'b0110101011: data <= 17'h1ff99; 
        10'b0110101100: data <= 17'h1ff5e; 
        10'b0110101101: data <= 17'h1fe1c; 
        10'b0110101110: data <= 17'h1fde1; 
        10'b0110101111: data <= 17'h1ff77; 
        10'b0110110000: data <= 17'h000c7; 
        10'b0110110001: data <= 17'h00274; 
        10'b0110110010: data <= 17'h0041a; 
        10'b0110110011: data <= 17'h00173; 
        10'b0110110100: data <= 17'h00044; 
        10'b0110110101: data <= 17'h1fd6b; 
        10'b0110110110: data <= 17'h1fdb6; 
        10'b0110110111: data <= 17'h1fe99; 
        10'b0110111000: data <= 17'h1ff28; 
        10'b0110111001: data <= 17'h1ff65; 
        10'b0110111010: data <= 17'h1ffd9; 
        10'b0110111011: data <= 17'h0000c; 
        10'b0110111100: data <= 17'h00038; 
        10'b0110111101: data <= 17'h00048; 
        10'b0110111110: data <= 17'h00094; 
        10'b0110111111: data <= 17'h00019; 
        10'b0111000000: data <= 17'h0009a; 
        10'b0111000001: data <= 17'h0004b; 
        10'b0111000010: data <= 17'h0008c; 
        10'b0111000011: data <= 17'h00056; 
        10'b0111000100: data <= 17'h0002d; 
        10'b0111000101: data <= 17'h1ffc2; 
        10'b0111000110: data <= 17'h1ff71; 
        10'b0111000111: data <= 17'h1ff67; 
        10'b0111001000: data <= 17'h1fe89; 
        10'b0111001001: data <= 17'h1ff20; 
        10'b0111001010: data <= 17'h1ff4d; 
        10'b0111001011: data <= 17'h1ff9d; 
        10'b0111001100: data <= 17'h1ffe7; 
        10'b0111001101: data <= 17'h0033a; 
        10'b0111001110: data <= 17'h003df; 
        10'b0111001111: data <= 17'h00039; 
        10'b0111010000: data <= 17'h1fecd; 
        10'b0111010001: data <= 17'h1fd35; 
        10'b0111010010: data <= 17'h1fdb0; 
        10'b0111010011: data <= 17'h1fe83; 
        10'b0111010100: data <= 17'h1fedf; 
        10'b0111010101: data <= 17'h1ff85; 
        10'b0111010110: data <= 17'h1ff83; 
        10'b0111010111: data <= 17'h00002; 
        10'b0111011000: data <= 17'h1ffc9; 
        10'b0111011001: data <= 17'h00009; 
        10'b0111011010: data <= 17'h00026; 
        10'b0111011011: data <= 17'h00050; 
        10'b0111011100: data <= 17'h00040; 
        10'b0111011101: data <= 17'h00098; 
        10'b0111011110: data <= 17'h00022; 
        10'b0111011111: data <= 17'h00096; 
        10'b0111100000: data <= 17'h0006f; 
        10'b0111100001: data <= 17'h1ffa9; 
        10'b0111100010: data <= 17'h1fec6; 
        10'b0111100011: data <= 17'h1feac; 
        10'b0111100100: data <= 17'h1ff0d; 
        10'b0111100101: data <= 17'h1ff64; 
        10'b0111100110: data <= 17'h00070; 
        10'b0111100111: data <= 17'h00001; 
        10'b0111101000: data <= 17'h0010e; 
        10'b0111101001: data <= 17'h003b2; 
        10'b0111101010: data <= 17'h0032c; 
        10'b0111101011: data <= 17'h1ff5b; 
        10'b0111101100: data <= 17'h1fdcc; 
        10'b0111101101: data <= 17'h1fd32; 
        10'b0111101110: data <= 17'h1fdb4; 
        10'b0111101111: data <= 17'h1fe8c; 
        10'b0111110000: data <= 17'h1ff74; 
        10'b0111110001: data <= 17'h1ffba; 
        10'b0111110010: data <= 17'h1ffce; 
        10'b0111110011: data <= 17'h1ffbd; 
        10'b0111110100: data <= 17'h1ff8c; 
        10'b0111110101: data <= 17'h00021; 
        10'b0111110110: data <= 17'h00058; 
        10'b0111110111: data <= 17'h00067; 
        10'b0111111000: data <= 17'h0005e; 
        10'b0111111001: data <= 17'h00056; 
        10'b0111111010: data <= 17'h00035; 
        10'b0111111011: data <= 17'h0007d; 
        10'b0111111100: data <= 17'h00045; 
        10'b0111111101: data <= 17'h1ff84; 
        10'b0111111110: data <= 17'h1feb1; 
        10'b0111111111: data <= 17'h1feb4; 
        10'b1000000000: data <= 17'h1ff83; 
        10'b1000000001: data <= 17'h0007f; 
        10'b1000000010: data <= 17'h00069; 
        10'b1000000011: data <= 17'h000a8; 
        10'b1000000100: data <= 17'h001b7; 
        10'b1000000101: data <= 17'h002c3; 
        10'b1000000110: data <= 17'h001e9; 
        10'b1000000111: data <= 17'h1febf; 
        10'b1000001000: data <= 17'h1fdf0; 
        10'b1000001001: data <= 17'h1fe3c; 
        10'b1000001010: data <= 17'h1fe7e; 
        10'b1000001011: data <= 17'h1fefd; 
        10'b1000001100: data <= 17'h1ff81; 
        10'b1000001101: data <= 17'h1ff29; 
        10'b1000001110: data <= 17'h1ffa1; 
        10'b1000001111: data <= 17'h1ff6d; 
        10'b1000010000: data <= 17'h1ffa6; 
        10'b1000010001: data <= 17'h00051; 
        10'b1000010010: data <= 17'h0008d; 
        10'b1000010011: data <= 17'h00090; 
        10'b1000010100: data <= 17'h00094; 
        10'b1000010101: data <= 17'h00068; 
        10'b1000010110: data <= 17'h0006c; 
        10'b1000010111: data <= 17'h00078; 
        10'b1000011000: data <= 17'h0000e; 
        10'b1000011001: data <= 17'h1ff46; 
        10'b1000011010: data <= 17'h1fe60; 
        10'b1000011011: data <= 17'h1fee8; 
        10'b1000011100: data <= 17'h1ff8e; 
        10'b1000011101: data <= 17'h00042; 
        10'b1000011110: data <= 17'h00021; 
        10'b1000011111: data <= 17'h00017; 
        10'b1000100000: data <= 17'h0003a; 
        10'b1000100001: data <= 17'h00146; 
        10'b1000100010: data <= 17'h00048; 
        10'b1000100011: data <= 17'h1fef6; 
        10'b1000100100: data <= 17'h1ff23; 
        10'b1000100101: data <= 17'h1ff3f; 
        10'b1000100110: data <= 17'h1ff0e; 
        10'b1000100111: data <= 17'h1ff44; 
        10'b1000101000: data <= 17'h1feed; 
        10'b1000101001: data <= 17'h1ff1b; 
        10'b1000101010: data <= 17'h1ff76; 
        10'b1000101011: data <= 17'h1ff86; 
        10'b1000101100: data <= 17'h00007; 
        10'b1000101101: data <= 17'h0002f; 
        10'b1000101110: data <= 17'h00033; 
        10'b1000101111: data <= 17'h00014; 
        10'b1000110000: data <= 17'h00018; 
        10'b1000110001: data <= 17'h0009b; 
        10'b1000110010: data <= 17'h00054; 
        10'b1000110011: data <= 17'h00036; 
        10'b1000110100: data <= 17'h1ffd6; 
        10'b1000110101: data <= 17'h1ff7c; 
        10'b1000110110: data <= 17'h1ffe7; 
        10'b1000110111: data <= 17'h1ffa5; 
        10'b1000111000: data <= 17'h1fffe; 
        10'b1000111001: data <= 17'h00027; 
        10'b1000111010: data <= 17'h1ff9a; 
        10'b1000111011: data <= 17'h1ffdb; 
        10'b1000111100: data <= 17'h1ff59; 
        10'b1000111101: data <= 17'h1ffc7; 
        10'b1000111110: data <= 17'h1ffd6; 
        10'b1000111111: data <= 17'h0000b; 
        10'b1001000000: data <= 17'h0009e; 
        10'b1001000001: data <= 17'h00039; 
        10'b1001000010: data <= 17'h1ffc4; 
        10'b1001000011: data <= 17'h1ff22; 
        10'b1001000100: data <= 17'h1feef; 
        10'b1001000101: data <= 17'h1ff03; 
        10'b1001000110: data <= 17'h1ff39; 
        10'b1001000111: data <= 17'h1ffd3; 
        10'b1001001000: data <= 17'h00015; 
        10'b1001001001: data <= 17'h0007f; 
        10'b1001001010: data <= 17'h00033; 
        10'b1001001011: data <= 17'h0009c; 
        10'b1001001100: data <= 17'h0006f; 
        10'b1001001101: data <= 17'h0003a; 
        10'b1001001110: data <= 17'h0005b; 
        10'b1001001111: data <= 17'h0006d; 
        10'b1001010000: data <= 17'h00056; 
        10'b1001010001: data <= 17'h000e9; 
        10'b1001010010: data <= 17'h000bf; 
        10'b1001010011: data <= 17'h0005a; 
        10'b1001010100: data <= 17'h0000f; 
        10'b1001010101: data <= 17'h1ffbe; 
        10'b1001010110: data <= 17'h00003; 
        10'b1001010111: data <= 17'h1ff7a; 
        10'b1001011000: data <= 17'h1fecf; 
        10'b1001011001: data <= 17'h1fea4; 
        10'b1001011010: data <= 17'h1ffe1; 
        10'b1001011011: data <= 17'h00069; 
        10'b1001011100: data <= 17'h000a7; 
        10'b1001011101: data <= 17'h000be; 
        10'b1001011110: data <= 17'h00083; 
        10'b1001011111: data <= 17'h1ff23; 
        10'b1001100000: data <= 17'h1ff26; 
        10'b1001100001: data <= 17'h1ff08; 
        10'b1001100010: data <= 17'h1ff55; 
        10'b1001100011: data <= 17'h1ff9d; 
        10'b1001100100: data <= 17'h00016; 
        10'b1001100101: data <= 17'h00043; 
        10'b1001100110: data <= 17'h0000d; 
        10'b1001100111: data <= 17'h00013; 
        10'b1001101000: data <= 17'h00056; 
        10'b1001101001: data <= 17'h00058; 
        10'b1001101010: data <= 17'h00063; 
        10'b1001101011: data <= 17'h00014; 
        10'b1001101100: data <= 17'h000ca; 
        10'b1001101101: data <= 17'h001c2; 
        10'b1001101110: data <= 17'h001d3; 
        10'b1001101111: data <= 17'h0011a; 
        10'b1001110000: data <= 17'h00026; 
        10'b1001110001: data <= 17'h1ffe1; 
        10'b1001110010: data <= 17'h1ff95; 
        10'b1001110011: data <= 17'h1fe43; 
        10'b1001110100: data <= 17'h1fd2e; 
        10'b1001110101: data <= 17'h1fdd8; 
        10'b1001110110: data <= 17'h00002; 
        10'b1001110111: data <= 17'h0006c; 
        10'b1001111000: data <= 17'h0019e; 
        10'b1001111001: data <= 17'h002a6; 
        10'b1001111010: data <= 17'h00129; 
        10'b1001111011: data <= 17'h0003e; 
        10'b1001111100: data <= 17'h1ff67; 
        10'b1001111101: data <= 17'h1ff89; 
        10'b1001111110: data <= 17'h1fff5; 
        10'b1001111111: data <= 17'h00014; 
        10'b1010000000: data <= 17'h0000a; 
        10'b1010000001: data <= 17'h00042; 
        10'b1010000010: data <= 17'h00096; 
        10'b1010000011: data <= 17'h00048; 
        10'b1010000100: data <= 17'h0008c; 
        10'b1010000101: data <= 17'h00057; 
        10'b1010000110: data <= 17'h00070; 
        10'b1010000111: data <= 17'h0003e; 
        10'b1010001000: data <= 17'h000b4; 
        10'b1010001001: data <= 17'h00183; 
        10'b1010001010: data <= 17'h0019d; 
        10'b1010001011: data <= 17'h000bd; 
        10'b1010001100: data <= 17'h00034; 
        10'b1010001101: data <= 17'h1ffa0; 
        10'b1010001110: data <= 17'h1ffbf; 
        10'b1010001111: data <= 17'h1ff05; 
        10'b1010010000: data <= 17'h1ff50; 
        10'b1010010001: data <= 17'h1ff63; 
        10'b1010010010: data <= 17'h1ff2e; 
        10'b1010010011: data <= 17'h00052; 
        10'b1010010100: data <= 17'h001e1; 
        10'b1010010101: data <= 17'h00244; 
        10'b1010010110: data <= 17'h00105; 
        10'b1010010111: data <= 17'h1ffd2; 
        10'b1010011000: data <= 17'h1ff91; 
        10'b1010011001: data <= 17'h1ff54; 
        10'b1010011010: data <= 17'h1ffc5; 
        10'b1010011011: data <= 17'h1ffca; 
        10'b1010011100: data <= 17'h00022; 
        10'b1010011101: data <= 17'h00011; 
        10'b1010011110: data <= 17'h00020; 
        10'b1010011111: data <= 17'h00010; 
        10'b1010100000: data <= 17'h00022; 
        10'b1010100001: data <= 17'h00016; 
        10'b1010100010: data <= 17'h00039; 
        10'b1010100011: data <= 17'h00012; 
        10'b1010100100: data <= 17'h00058; 
        10'b1010100101: data <= 17'h000ab; 
        10'b1010100110: data <= 17'h000b1; 
        10'b1010100111: data <= 17'h1ffc7; 
        10'b1010101000: data <= 17'h1feff; 
        10'b1010101001: data <= 17'h1fefe; 
        10'b1010101010: data <= 17'h1fe3b; 
        10'b1010101011: data <= 17'h1fe4e; 
        10'b1010101100: data <= 17'h1fe7b; 
        10'b1010101101: data <= 17'h1feb2; 
        10'b1010101110: data <= 17'h1feb4; 
        10'b1010101111: data <= 17'h1feb3; 
        10'b1010110000: data <= 17'h1ffa0; 
        10'b1010110001: data <= 17'h00028; 
        10'b1010110010: data <= 17'h00049; 
        10'b1010110011: data <= 17'h0006a; 
        10'b1010110100: data <= 17'h00059; 
        10'b1010110101: data <= 17'h00016; 
        10'b1010110110: data <= 17'h0002e; 
        10'b1010110111: data <= 17'h0007c; 
        10'b1010111000: data <= 17'h00025; 
        10'b1010111001: data <= 17'h0003d; 
        10'b1010111010: data <= 17'h00075; 
        10'b1010111011: data <= 17'h00027; 
        10'b1010111100: data <= 17'h00098; 
        10'b1010111101: data <= 17'h00030; 
        10'b1010111110: data <= 17'h0003a; 
        10'b1010111111: data <= 17'h00052; 
        10'b1011000000: data <= 17'h00075; 
        10'b1011000001: data <= 17'h0006b; 
        10'b1011000010: data <= 17'h00002; 
        10'b1011000011: data <= 17'h1ffbe; 
        10'b1011000100: data <= 17'h1ffe6; 
        10'b1011000101: data <= 17'h1ffc3; 
        10'b1011000110: data <= 17'h1ff03; 
        10'b1011000111: data <= 17'h1fecb; 
        10'b1011001000: data <= 17'h1ff1c; 
        10'b1011001001: data <= 17'h1fec0; 
        10'b1011001010: data <= 17'h1ff3c; 
        10'b1011001011: data <= 17'h1ff08; 
        10'b1011001100: data <= 17'h1ff71; 
        10'b1011001101: data <= 17'h1ffe6; 
        10'b1011001110: data <= 17'h00031; 
        10'b1011001111: data <= 17'h00066; 
        10'b1011010000: data <= 17'h0000a; 
        10'b1011010001: data <= 17'h0005d; 
        10'b1011010010: data <= 17'h00037; 
        10'b1011010011: data <= 17'h00085; 
        10'b1011010100: data <= 17'h00021; 
        10'b1011010101: data <= 17'h00028; 
        10'b1011010110: data <= 17'h00039; 
        10'b1011010111: data <= 17'h00031; 
        10'b1011011000: data <= 17'h00038; 
        10'b1011011001: data <= 17'h0006b; 
        10'b1011011010: data <= 17'h00060; 
        10'b1011011011: data <= 17'h0001d; 
        10'b1011011100: data <= 17'h00067; 
        10'b1011011101: data <= 17'h00089; 
        10'b1011011110: data <= 17'h0005d; 
        10'b1011011111: data <= 17'h00056; 
        10'b1011100000: data <= 17'h0007b; 
        10'b1011100001: data <= 17'h00068; 
        10'b1011100010: data <= 17'h0000e; 
        10'b1011100011: data <= 17'h00055; 
        10'b1011100100: data <= 17'h0004d; 
        10'b1011100101: data <= 17'h0002d; 
        10'b1011100110: data <= 17'h1fffd; 
        10'b1011100111: data <= 17'h00028; 
        10'b1011101000: data <= 17'h0005a; 
        10'b1011101001: data <= 17'h0008b; 
        10'b1011101010: data <= 17'h00067; 
        10'b1011101011: data <= 17'h00010; 
        10'b1011101100: data <= 17'h00060; 
        10'b1011101101: data <= 17'h0005a; 
        10'b1011101110: data <= 17'h00056; 
        10'b1011101111: data <= 17'h00029; 
        10'b1011110000: data <= 17'h00024; 
        10'b1011110001: data <= 17'h00068; 
        10'b1011110010: data <= 17'h0008e; 
        10'b1011110011: data <= 17'h00073; 
        10'b1011110100: data <= 17'h00074; 
        10'b1011110101: data <= 17'h00092; 
        10'b1011110110: data <= 17'h00017; 
        10'b1011110111: data <= 17'h00051; 
        10'b1011111000: data <= 17'h0009a; 
        10'b1011111001: data <= 17'h0007a; 
        10'b1011111010: data <= 17'h0008a; 
        10'b1011111011: data <= 17'h00080; 
        10'b1011111100: data <= 17'h0008a; 
        10'b1011111101: data <= 17'h00041; 
        10'b1011111110: data <= 17'h00079; 
        10'b1011111111: data <= 17'h0007e; 
        10'b1100000000: data <= 17'h0000d; 
        10'b1100000001: data <= 17'h0001a; 
        10'b1100000010: data <= 17'h00097; 
        10'b1100000011: data <= 17'h00062; 
        10'b1100000100: data <= 17'h0005b; 
        10'b1100000101: data <= 17'h0000d; 
        10'b1100000110: data <= 17'h00042; 
        10'b1100000111: data <= 17'h0001d; 
        10'b1100001000: data <= 17'h0001b; 
        10'b1100001001: data <= 17'h00031; 
        10'b1100001010: data <= 17'h00059; 
        10'b1100001011: data <= 17'h00080; 
        10'b1100001100: data <= 17'h0008e; 
        10'b1100001101: data <= 17'h0008a; 
        10'b1100001110: data <= 17'h00088; 
        10'b1100001111: data <= 17'h0002e; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 12) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 18'h000ff; 
        10'b0000000001: data <= 18'h0007a; 
        10'b0000000010: data <= 18'h00088; 
        10'b0000000011: data <= 18'h00038; 
        10'b0000000100: data <= 18'h000d8; 
        10'b0000000101: data <= 18'h000d3; 
        10'b0000000110: data <= 18'h000e9; 
        10'b0000000111: data <= 18'h0003a; 
        10'b0000001000: data <= 18'h000cb; 
        10'b0000001001: data <= 18'h0003e; 
        10'b0000001010: data <= 18'h000c1; 
        10'b0000001011: data <= 18'h0009c; 
        10'b0000001100: data <= 18'h000d9; 
        10'b0000001101: data <= 18'h00122; 
        10'b0000001110: data <= 18'h000ff; 
        10'b0000001111: data <= 18'h000af; 
        10'b0000010000: data <= 18'h000b1; 
        10'b0000010001: data <= 18'h0003e; 
        10'b0000010010: data <= 18'h00129; 
        10'b0000010011: data <= 18'h00128; 
        10'b0000010100: data <= 18'h000a9; 
        10'b0000010101: data <= 18'h000d9; 
        10'b0000010110: data <= 18'h000a7; 
        10'b0000010111: data <= 18'h00103; 
        10'b0000011000: data <= 18'h00063; 
        10'b0000011001: data <= 18'h00112; 
        10'b0000011010: data <= 18'h000a7; 
        10'b0000011011: data <= 18'h000f2; 
        10'b0000011100: data <= 18'h0001f; 
        10'b0000011101: data <= 18'h00101; 
        10'b0000011110: data <= 18'h0004c; 
        10'b0000011111: data <= 18'h000b7; 
        10'b0000100000: data <= 18'h000a3; 
        10'b0000100001: data <= 18'h00041; 
        10'b0000100010: data <= 18'h0005b; 
        10'b0000100011: data <= 18'h000f1; 
        10'b0000100100: data <= 18'h000e8; 
        10'b0000100101: data <= 18'h000bc; 
        10'b0000100110: data <= 18'h000ba; 
        10'b0000100111: data <= 18'h00089; 
        10'b0000101000: data <= 18'h000de; 
        10'b0000101001: data <= 18'h000fa; 
        10'b0000101010: data <= 18'h00143; 
        10'b0000101011: data <= 18'h000a1; 
        10'b0000101100: data <= 18'h00082; 
        10'b0000101101: data <= 18'h00104; 
        10'b0000101110: data <= 18'h000af; 
        10'b0000101111: data <= 18'h00077; 
        10'b0000110000: data <= 18'h00119; 
        10'b0000110001: data <= 18'h0010f; 
        10'b0000110010: data <= 18'h0006f; 
        10'b0000110011: data <= 18'h00122; 
        10'b0000110100: data <= 18'h00137; 
        10'b0000110101: data <= 18'h000a5; 
        10'b0000110110: data <= 18'h00109; 
        10'b0000110111: data <= 18'h000d5; 
        10'b0000111000: data <= 18'h00105; 
        10'b0000111001: data <= 18'h000c4; 
        10'b0000111010: data <= 18'h00139; 
        10'b0000111011: data <= 18'h0003d; 
        10'b0000111100: data <= 18'h0003a; 
        10'b0000111101: data <= 18'h000ce; 
        10'b0000111110: data <= 18'h00098; 
        10'b0000111111: data <= 18'h00093; 
        10'b0001000000: data <= 18'h00063; 
        10'b0001000001: data <= 18'h000ad; 
        10'b0001000010: data <= 18'h00004; 
        10'b0001000011: data <= 18'h00057; 
        10'b0001000100: data <= 18'h0000b; 
        10'b0001000101: data <= 18'h0004c; 
        10'b0001000110: data <= 18'h0009f; 
        10'b0001000111: data <= 18'h000ff; 
        10'b0001001000: data <= 18'h000c1; 
        10'b0001001001: data <= 18'h00000; 
        10'b0001001010: data <= 18'h000bf; 
        10'b0001001011: data <= 18'h00072; 
        10'b0001001100: data <= 18'h000fb; 
        10'b0001001101: data <= 18'h0006d; 
        10'b0001001110: data <= 18'h00114; 
        10'b0001001111: data <= 18'h000c9; 
        10'b0001010000: data <= 18'h000d8; 
        10'b0001010001: data <= 18'h00025; 
        10'b0001010010: data <= 18'h000eb; 
        10'b0001010011: data <= 18'h000f0; 
        10'b0001010100: data <= 18'h0005d; 
        10'b0001010101: data <= 18'h00068; 
        10'b0001010110: data <= 18'h000b0; 
        10'b0001010111: data <= 18'h00091; 
        10'b0001011000: data <= 18'h00126; 
        10'b0001011001: data <= 18'h0009b; 
        10'b0001011010: data <= 18'h00022; 
        10'b0001011011: data <= 18'h00120; 
        10'b0001011100: data <= 18'h3ffe0; 
        10'b0001011101: data <= 18'h3ffc6; 
        10'b0001011110: data <= 18'h3ffc8; 
        10'b0001011111: data <= 18'h3ff60; 
        10'b0001100000: data <= 18'h3ffc7; 
        10'b0001100001: data <= 18'h00015; 
        10'b0001100010: data <= 18'h00078; 
        10'b0001100011: data <= 18'h000f0; 
        10'b0001100100: data <= 18'h3ff89; 
        10'b0001100101: data <= 18'h3ffd5; 
        10'b0001100110: data <= 18'h3fffa; 
        10'b0001100111: data <= 18'h3ff47; 
        10'b0001101000: data <= 18'h3ffed; 
        10'b0001101001: data <= 18'h0004c; 
        10'b0001101010: data <= 18'h000c0; 
        10'b0001101011: data <= 18'h000bb; 
        10'b0001101100: data <= 18'h3ffde; 
        10'b0001101101: data <= 18'h0010a; 
        10'b0001101110: data <= 18'h00064; 
        10'b0001101111: data <= 18'h00118; 
        10'b0001110000: data <= 18'h000d8; 
        10'b0001110001: data <= 18'h00083; 
        10'b0001110010: data <= 18'h0012a; 
        10'b0001110011: data <= 18'h00127; 
        10'b0001110100: data <= 18'h00021; 
        10'b0001110101: data <= 18'h0003b; 
        10'b0001110110: data <= 18'h00104; 
        10'b0001110111: data <= 18'h000a5; 
        10'b0001111000: data <= 18'h0003f; 
        10'b0001111001: data <= 18'h3fef0; 
        10'b0001111010: data <= 18'h00019; 
        10'b0001111011: data <= 18'h0005f; 
        10'b0001111100: data <= 18'h00094; 
        10'b0001111101: data <= 18'h00108; 
        10'b0001111110: data <= 18'h00136; 
        10'b0001111111: data <= 18'h0027a; 
        10'b0010000000: data <= 18'h000ad; 
        10'b0010000001: data <= 18'h3ff7b; 
        10'b0010000010: data <= 18'h3ff6f; 
        10'b0010000011: data <= 18'h00062; 
        10'b0010000100: data <= 18'h0015f; 
        10'b0010000101: data <= 18'h00189; 
        10'b0010000110: data <= 18'h00187; 
        10'b0010000111: data <= 18'h001ca; 
        10'b0010001000: data <= 18'h000ef; 
        10'b0010001001: data <= 18'h00071; 
        10'b0010001010: data <= 18'h00063; 
        10'b0010001011: data <= 18'h0006d; 
        10'b0010001100: data <= 18'h00027; 
        10'b0010001101: data <= 18'h00100; 
        10'b0010001110: data <= 18'h00032; 
        10'b0010001111: data <= 18'h000b4; 
        10'b0010010000: data <= 18'h0002d; 
        10'b0010010001: data <= 18'h000ac; 
        10'b0010010010: data <= 18'h00034; 
        10'b0010010011: data <= 18'h3ffbd; 
        10'b0010010100: data <= 18'h3fdc6; 
        10'b0010010101: data <= 18'h3fdc1; 
        10'b0010010110: data <= 18'h3fef8; 
        10'b0010010111: data <= 18'h00003; 
        10'b0010011000: data <= 18'h000d8; 
        10'b0010011001: data <= 18'h000f3; 
        10'b0010011010: data <= 18'h001a7; 
        10'b0010011011: data <= 18'h00148; 
        10'b0010011100: data <= 18'h000c2; 
        10'b0010011101: data <= 18'h3fec1; 
        10'b0010011110: data <= 18'h3ffe0; 
        10'b0010011111: data <= 18'h00043; 
        10'b0010100000: data <= 18'h00138; 
        10'b0010100001: data <= 18'h001f7; 
        10'b0010100010: data <= 18'h00344; 
        10'b0010100011: data <= 18'h0020a; 
        10'b0010100100: data <= 18'h001ab; 
        10'b0010100101: data <= 18'h3ff92; 
        10'b0010100110: data <= 18'h00076; 
        10'b0010100111: data <= 18'h00041; 
        10'b0010101000: data <= 18'h00036; 
        10'b0010101001: data <= 18'h000b9; 
        10'b0010101010: data <= 18'h00022; 
        10'b0010101011: data <= 18'h00090; 
        10'b0010101100: data <= 18'h00022; 
        10'b0010101101: data <= 18'h3ffab; 
        10'b0010101110: data <= 18'h3fec6; 
        10'b0010101111: data <= 18'h3feca; 
        10'b0010110000: data <= 18'h3fd37; 
        10'b0010110001: data <= 18'h3fca2; 
        10'b0010110010: data <= 18'h3fde4; 
        10'b0010110011: data <= 18'h3ff81; 
        10'b0010110100: data <= 18'h3ff7c; 
        10'b0010110101: data <= 18'h3fef1; 
        10'b0010110110: data <= 18'h3ff83; 
        10'b0010110111: data <= 18'h3fd95; 
        10'b0010111000: data <= 18'h3fd67; 
        10'b0010111001: data <= 18'h3fd62; 
        10'b0010111010: data <= 18'h3fee8; 
        10'b0010111011: data <= 18'h3ff31; 
        10'b0010111100: data <= 18'h0013a; 
        10'b0010111101: data <= 18'h00204; 
        10'b0010111110: data <= 18'h001df; 
        10'b0010111111: data <= 18'h00193; 
        10'b0011000000: data <= 18'h00069; 
        10'b0011000001: data <= 18'h3ffaa; 
        10'b0011000010: data <= 18'h00007; 
        10'b0011000011: data <= 18'h00097; 
        10'b0011000100: data <= 18'h0007a; 
        10'b0011000101: data <= 18'h00045; 
        10'b0011000110: data <= 18'h00055; 
        10'b0011000111: data <= 18'h00013; 
        10'b0011001000: data <= 18'h000ca; 
        10'b0011001001: data <= 18'h3ffd5; 
        10'b0011001010: data <= 18'h3fed3; 
        10'b0011001011: data <= 18'h3fd98; 
        10'b0011001100: data <= 18'h3fc3e; 
        10'b0011001101: data <= 18'h3fb37; 
        10'b0011001110: data <= 18'h3fcc0; 
        10'b0011001111: data <= 18'h3fe94; 
        10'b0011010000: data <= 18'h3feb3; 
        10'b0011010001: data <= 18'h3fe21; 
        10'b0011010010: data <= 18'h3fdb0; 
        10'b0011010011: data <= 18'h3fc68; 
        10'b0011010100: data <= 18'h3fcdc; 
        10'b0011010101: data <= 18'h3fd0e; 
        10'b0011010110: data <= 18'h3fd58; 
        10'b0011010111: data <= 18'h3ffe9; 
        10'b0011011000: data <= 18'h0008f; 
        10'b0011011001: data <= 18'h00059; 
        10'b0011011010: data <= 18'h00054; 
        10'b0011011011: data <= 18'h3fefd; 
        10'b0011011100: data <= 18'h3fe9f; 
        10'b0011011101: data <= 18'h3ff73; 
        10'b0011011110: data <= 18'h00073; 
        10'b0011011111: data <= 18'h00086; 
        10'b0011100000: data <= 18'h00095; 
        10'b0011100001: data <= 18'h0007e; 
        10'b0011100010: data <= 18'h0007b; 
        10'b0011100011: data <= 18'h00106; 
        10'b0011100100: data <= 18'h00054; 
        10'b0011100101: data <= 18'h3fff8; 
        10'b0011100110: data <= 18'h3fe9a; 
        10'b0011100111: data <= 18'h3fde1; 
        10'b0011101000: data <= 18'h3fb9f; 
        10'b0011101001: data <= 18'h3fb3e; 
        10'b0011101010: data <= 18'h3fb79; 
        10'b0011101011: data <= 18'h3fd90; 
        10'b0011101100: data <= 18'h3fee2; 
        10'b0011101101: data <= 18'h3fea0; 
        10'b0011101110: data <= 18'h3fee1; 
        10'b0011101111: data <= 18'h0007e; 
        10'b0011110000: data <= 18'h3fe02; 
        10'b0011110001: data <= 18'h3ff53; 
        10'b0011110010: data <= 18'h3ffe3; 
        10'b0011110011: data <= 18'h00042; 
        10'b0011110100: data <= 18'h3fe80; 
        10'b0011110101: data <= 18'h3fe8d; 
        10'b0011110110: data <= 18'h3fdae; 
        10'b0011110111: data <= 18'h3fcf5; 
        10'b0011111000: data <= 18'h3fd94; 
        10'b0011111001: data <= 18'h3ff68; 
        10'b0011111010: data <= 18'h000e7; 
        10'b0011111011: data <= 18'h00130; 
        10'b0011111100: data <= 18'h00133; 
        10'b0011111101: data <= 18'h00047; 
        10'b0011111110: data <= 18'h0007e; 
        10'b0011111111: data <= 18'h0006c; 
        10'b0100000000: data <= 18'h3ffed; 
        10'b0100000001: data <= 18'h3ffde; 
        10'b0100000010: data <= 18'h3fe38; 
        10'b0100000011: data <= 18'h3fe50; 
        10'b0100000100: data <= 18'h3fcfc; 
        10'b0100000101: data <= 18'h3fb67; 
        10'b0100000110: data <= 18'h3fbca; 
        10'b0100000111: data <= 18'h3fe56; 
        10'b0100001000: data <= 18'h3fec2; 
        10'b0100001001: data <= 18'h000f2; 
        10'b0100001010: data <= 18'h002f9; 
        10'b0100001011: data <= 18'h00442; 
        10'b0100001100: data <= 18'h00194; 
        10'b0100001101: data <= 18'h3ffe4; 
        10'b0100001110: data <= 18'h3ff4a; 
        10'b0100001111: data <= 18'h3fd1c; 
        10'b0100010000: data <= 18'h3fc72; 
        10'b0100010001: data <= 18'h3fc7f; 
        10'b0100010010: data <= 18'h3fb95; 
        10'b0100010011: data <= 18'h3fc2c; 
        10'b0100010100: data <= 18'h3fdf2; 
        10'b0100010101: data <= 18'h0003d; 
        10'b0100010110: data <= 18'h000fe; 
        10'b0100010111: data <= 18'h000b8; 
        10'b0100011000: data <= 18'h00118; 
        10'b0100011001: data <= 18'h00136; 
        10'b0100011010: data <= 18'h00100; 
        10'b0100011011: data <= 18'h00022; 
        10'b0100011100: data <= 18'h000d1; 
        10'b0100011101: data <= 18'h3ff0d; 
        10'b0100011110: data <= 18'h3fe51; 
        10'b0100011111: data <= 18'h3ff38; 
        10'b0100100000: data <= 18'h3fda9; 
        10'b0100100001: data <= 18'h3fda1; 
        10'b0100100010: data <= 18'h3fe44; 
        10'b0100100011: data <= 18'h3fed8; 
        10'b0100100100: data <= 18'h3ff38; 
        10'b0100100101: data <= 18'h00260; 
        10'b0100100110: data <= 18'h007b0; 
        10'b0100100111: data <= 18'h0081d; 
        10'b0100101000: data <= 18'h003db; 
        10'b0100101001: data <= 18'h3ffeb; 
        10'b0100101010: data <= 18'h3fdb2; 
        10'b0100101011: data <= 18'h3fd38; 
        10'b0100101100: data <= 18'h3fca2; 
        10'b0100101101: data <= 18'h3fcf7; 
        10'b0100101110: data <= 18'h3fd24; 
        10'b0100101111: data <= 18'h3fe39; 
        10'b0100110000: data <= 18'h3ff68; 
        10'b0100110001: data <= 18'h3ffe6; 
        10'b0100110010: data <= 18'h00107; 
        10'b0100110011: data <= 18'h0006c; 
        10'b0100110100: data <= 18'h00035; 
        10'b0100110101: data <= 18'h0002f; 
        10'b0100110110: data <= 18'h000d5; 
        10'b0100110111: data <= 18'h000e3; 
        10'b0100111000: data <= 18'h00001; 
        10'b0100111001: data <= 18'h3ffbb; 
        10'b0100111010: data <= 18'h3ffdc; 
        10'b0100111011: data <= 18'h3fe8a; 
        10'b0100111100: data <= 18'h3ff0e; 
        10'b0100111101: data <= 18'h3fe8a; 
        10'b0100111110: data <= 18'h3fdda; 
        10'b0100111111: data <= 18'h3fcc2; 
        10'b0101000000: data <= 18'h3ffa1; 
        10'b0101000001: data <= 18'h00410; 
        10'b0101000010: data <= 18'h00944; 
        10'b0101000011: data <= 18'h009d1; 
        10'b0101000100: data <= 18'h003a3; 
        10'b0101000101: data <= 18'h3ff34; 
        10'b0101000110: data <= 18'h3ff45; 
        10'b0101000111: data <= 18'h3fe11; 
        10'b0101001000: data <= 18'h3fdf4; 
        10'b0101001001: data <= 18'h3fe19; 
        10'b0101001010: data <= 18'h3fe3d; 
        10'b0101001011: data <= 18'h3ff2d; 
        10'b0101001100: data <= 18'h3ffa7; 
        10'b0101001101: data <= 18'h000d1; 
        10'b0101001110: data <= 18'h00125; 
        10'b0101001111: data <= 18'h000ce; 
        10'b0101010000: data <= 18'h00020; 
        10'b0101010001: data <= 18'h00118; 
        10'b0101010010: data <= 18'h00086; 
        10'b0101010011: data <= 18'h0005b; 
        10'b0101010100: data <= 18'h0011e; 
        10'b0101010101: data <= 18'h3ffc9; 
        10'b0101010110: data <= 18'h3ffa8; 
        10'b0101010111: data <= 18'h3ff84; 
        10'b0101011000: data <= 18'h3fe9b; 
        10'b0101011001: data <= 18'h3fe2c; 
        10'b0101011010: data <= 18'h3fc22; 
        10'b0101011011: data <= 18'h3fa93; 
        10'b0101011100: data <= 18'h3ffd3; 
        10'b0101011101: data <= 18'h00420; 
        10'b0101011110: data <= 18'h00ae8; 
        10'b0101011111: data <= 18'h00791; 
        10'b0101100000: data <= 18'h0017f; 
        10'b0101100001: data <= 18'h000cb; 
        10'b0101100010: data <= 18'h3ff89; 
        10'b0101100011: data <= 18'h3fdca; 
        10'b0101100100: data <= 18'h3fe9b; 
        10'b0101100101: data <= 18'h3ff53; 
        10'b0101100110: data <= 18'h3ff9e; 
        10'b0101100111: data <= 18'h3ff88; 
        10'b0101101000: data <= 18'h00012; 
        10'b0101101001: data <= 18'h0011c; 
        10'b0101101010: data <= 18'h0002b; 
        10'b0101101011: data <= 18'h000c8; 
        10'b0101101100: data <= 18'h0001d; 
        10'b0101101101: data <= 18'h000be; 
        10'b0101101110: data <= 18'h000b1; 
        10'b0101101111: data <= 18'h000bd; 
        10'b0101110000: data <= 18'h0013b; 
        10'b0101110001: data <= 18'h00002; 
        10'b0101110010: data <= 18'h0001b; 
        10'b0101110011: data <= 18'h3ff73; 
        10'b0101110100: data <= 18'h3ff41; 
        10'b0101110101: data <= 18'h3fcf5; 
        10'b0101110110: data <= 18'h3f98b; 
        10'b0101110111: data <= 18'h3f973; 
        10'b0101111000: data <= 18'h00002; 
        10'b0101111001: data <= 18'h00370; 
        10'b0101111010: data <= 18'h008fd; 
        10'b0101111011: data <= 18'h00514; 
        10'b0101111100: data <= 18'h00158; 
        10'b0101111101: data <= 18'h000a7; 
        10'b0101111110: data <= 18'h3fdf3; 
        10'b0101111111: data <= 18'h3fd05; 
        10'b0110000000: data <= 18'h3feeb; 
        10'b0110000001: data <= 18'h3ff9e; 
        10'b0110000010: data <= 18'h3ff9a; 
        10'b0110000011: data <= 18'h3ffdb; 
        10'b0110000100: data <= 18'h00081; 
        10'b0110000101: data <= 18'h000c0; 
        10'b0110000110: data <= 18'h00115; 
        10'b0110000111: data <= 18'h000b4; 
        10'b0110001000: data <= 18'h0008c; 
        10'b0110001001: data <= 18'h0012c; 
        10'b0110001010: data <= 18'h000a9; 
        10'b0110001011: data <= 18'h000f0; 
        10'b0110001100: data <= 18'h000f1; 
        10'b0110001101: data <= 18'h3ffff; 
        10'b0110001110: data <= 18'h00029; 
        10'b0110001111: data <= 18'h3ffa4; 
        10'b0110010000: data <= 18'h3fdfd; 
        10'b0110010001: data <= 18'h3fc8b; 
        10'b0110010010: data <= 18'h3f991; 
        10'b0110010011: data <= 18'h3fb1e; 
        10'b0110010100: data <= 18'h3ffe4; 
        10'b0110010101: data <= 18'h0037e; 
        10'b0110010110: data <= 18'h007ab; 
        10'b0110010111: data <= 18'h004f0; 
        10'b0110011000: data <= 18'h0017a; 
        10'b0110011001: data <= 18'h3fd43; 
        10'b0110011010: data <= 18'h3fc4a; 
        10'b0110011011: data <= 18'h3fd2f; 
        10'b0110011100: data <= 18'h3fe55; 
        10'b0110011101: data <= 18'h3ff85; 
        10'b0110011110: data <= 18'h3ff7a; 
        10'b0110011111: data <= 18'h3ffa4; 
        10'b0110100000: data <= 18'h000d6; 
        10'b0110100001: data <= 18'h00021; 
        10'b0110100010: data <= 18'h0003b; 
        10'b0110100011: data <= 18'h000aa; 
        10'b0110100100: data <= 18'h0013e; 
        10'b0110100101: data <= 18'h00034; 
        10'b0110100110: data <= 18'h000cc; 
        10'b0110100111: data <= 18'h00081; 
        10'b0110101000: data <= 18'h00049; 
        10'b0110101001: data <= 18'h000b9; 
        10'b0110101010: data <= 18'h3ff4c; 
        10'b0110101011: data <= 18'h3ff33; 
        10'b0110101100: data <= 18'h3febb; 
        10'b0110101101: data <= 18'h3fc38; 
        10'b0110101110: data <= 18'h3fbc3; 
        10'b0110101111: data <= 18'h3feef; 
        10'b0110110000: data <= 18'h0018e; 
        10'b0110110001: data <= 18'h004e8; 
        10'b0110110010: data <= 18'h00834; 
        10'b0110110011: data <= 18'h002e7; 
        10'b0110110100: data <= 18'h00088; 
        10'b0110110101: data <= 18'h3fad6; 
        10'b0110110110: data <= 18'h3fb6d; 
        10'b0110110111: data <= 18'h3fd33; 
        10'b0110111000: data <= 18'h3fe50; 
        10'b0110111001: data <= 18'h3feca; 
        10'b0110111010: data <= 18'h3ffb2; 
        10'b0110111011: data <= 18'h00018; 
        10'b0110111100: data <= 18'h00070; 
        10'b0110111101: data <= 18'h0008f; 
        10'b0110111110: data <= 18'h00128; 
        10'b0110111111: data <= 18'h00031; 
        10'b0111000000: data <= 18'h00133; 
        10'b0111000001: data <= 18'h00096; 
        10'b0111000010: data <= 18'h00119; 
        10'b0111000011: data <= 18'h000ab; 
        10'b0111000100: data <= 18'h0005b; 
        10'b0111000101: data <= 18'h3ff83; 
        10'b0111000110: data <= 18'h3fee3; 
        10'b0111000111: data <= 18'h3fecd; 
        10'b0111001000: data <= 18'h3fd12; 
        10'b0111001001: data <= 18'h3fe3f; 
        10'b0111001010: data <= 18'h3fe9a; 
        10'b0111001011: data <= 18'h3ff3a; 
        10'b0111001100: data <= 18'h3ffce; 
        10'b0111001101: data <= 18'h00674; 
        10'b0111001110: data <= 18'h007bf; 
        10'b0111001111: data <= 18'h00072; 
        10'b0111010000: data <= 18'h3fd9a; 
        10'b0111010001: data <= 18'h3fa6a; 
        10'b0111010010: data <= 18'h3fb61; 
        10'b0111010011: data <= 18'h3fd06; 
        10'b0111010100: data <= 18'h3fdbd; 
        10'b0111010101: data <= 18'h3ff09; 
        10'b0111010110: data <= 18'h3ff05; 
        10'b0111010111: data <= 18'h00003; 
        10'b0111011000: data <= 18'h3ff91; 
        10'b0111011001: data <= 18'h00011; 
        10'b0111011010: data <= 18'h0004b; 
        10'b0111011011: data <= 18'h0009f; 
        10'b0111011100: data <= 18'h0007f; 
        10'b0111011101: data <= 18'h00130; 
        10'b0111011110: data <= 18'h00043; 
        10'b0111011111: data <= 18'h0012b; 
        10'b0111100000: data <= 18'h000dd; 
        10'b0111100001: data <= 18'h3ff52; 
        10'b0111100010: data <= 18'h3fd8c; 
        10'b0111100011: data <= 18'h3fd58; 
        10'b0111100100: data <= 18'h3fe19; 
        10'b0111100101: data <= 18'h3fec9; 
        10'b0111100110: data <= 18'h000e0; 
        10'b0111100111: data <= 18'h00003; 
        10'b0111101000: data <= 18'h0021c; 
        10'b0111101001: data <= 18'h00765; 
        10'b0111101010: data <= 18'h00657; 
        10'b0111101011: data <= 18'h3feb6; 
        10'b0111101100: data <= 18'h3fb98; 
        10'b0111101101: data <= 18'h3fa65; 
        10'b0111101110: data <= 18'h3fb68; 
        10'b0111101111: data <= 18'h3fd19; 
        10'b0111110000: data <= 18'h3fee9; 
        10'b0111110001: data <= 18'h3ff74; 
        10'b0111110010: data <= 18'h3ff9b; 
        10'b0111110011: data <= 18'h3ff79; 
        10'b0111110100: data <= 18'h3ff18; 
        10'b0111110101: data <= 18'h00042; 
        10'b0111110110: data <= 18'h000b1; 
        10'b0111110111: data <= 18'h000cf; 
        10'b0111111000: data <= 18'h000bc; 
        10'b0111111001: data <= 18'h000ad; 
        10'b0111111010: data <= 18'h0006a; 
        10'b0111111011: data <= 18'h000fa; 
        10'b0111111100: data <= 18'h0008b; 
        10'b0111111101: data <= 18'h3ff08; 
        10'b0111111110: data <= 18'h3fd62; 
        10'b0111111111: data <= 18'h3fd67; 
        10'b1000000000: data <= 18'h3ff07; 
        10'b1000000001: data <= 18'h000ff; 
        10'b1000000010: data <= 18'h000d2; 
        10'b1000000011: data <= 18'h00151; 
        10'b1000000100: data <= 18'h0036e; 
        10'b1000000101: data <= 18'h00586; 
        10'b1000000110: data <= 18'h003d2; 
        10'b1000000111: data <= 18'h3fd7d; 
        10'b1000001000: data <= 18'h3fbe0; 
        10'b1000001001: data <= 18'h3fc77; 
        10'b1000001010: data <= 18'h3fcfb; 
        10'b1000001011: data <= 18'h3fdfa; 
        10'b1000001100: data <= 18'h3ff02; 
        10'b1000001101: data <= 18'h3fe52; 
        10'b1000001110: data <= 18'h3ff41; 
        10'b1000001111: data <= 18'h3fedb; 
        10'b1000010000: data <= 18'h3ff4d; 
        10'b1000010001: data <= 18'h000a2; 
        10'b1000010010: data <= 18'h00119; 
        10'b1000010011: data <= 18'h0011f; 
        10'b1000010100: data <= 18'h00128; 
        10'b1000010101: data <= 18'h000d0; 
        10'b1000010110: data <= 18'h000d9; 
        10'b1000010111: data <= 18'h000f0; 
        10'b1000011000: data <= 18'h0001c; 
        10'b1000011001: data <= 18'h3fe8c; 
        10'b1000011010: data <= 18'h3fcc1; 
        10'b1000011011: data <= 18'h3fdcf; 
        10'b1000011100: data <= 18'h3ff1b; 
        10'b1000011101: data <= 18'h00084; 
        10'b1000011110: data <= 18'h00042; 
        10'b1000011111: data <= 18'h0002e; 
        10'b1000100000: data <= 18'h00074; 
        10'b1000100001: data <= 18'h0028b; 
        10'b1000100010: data <= 18'h0008f; 
        10'b1000100011: data <= 18'h3fded; 
        10'b1000100100: data <= 18'h3fe45; 
        10'b1000100101: data <= 18'h3fe7f; 
        10'b1000100110: data <= 18'h3fe1c; 
        10'b1000100111: data <= 18'h3fe89; 
        10'b1000101000: data <= 18'h3fddb; 
        10'b1000101001: data <= 18'h3fe36; 
        10'b1000101010: data <= 18'h3feec; 
        10'b1000101011: data <= 18'h3ff0d; 
        10'b1000101100: data <= 18'h0000d; 
        10'b1000101101: data <= 18'h0005d; 
        10'b1000101110: data <= 18'h00066; 
        10'b1000101111: data <= 18'h00029; 
        10'b1000110000: data <= 18'h0002f; 
        10'b1000110001: data <= 18'h00137; 
        10'b1000110010: data <= 18'h000a7; 
        10'b1000110011: data <= 18'h0006b; 
        10'b1000110100: data <= 18'h3ffad; 
        10'b1000110101: data <= 18'h3fef7; 
        10'b1000110110: data <= 18'h3ffce; 
        10'b1000110111: data <= 18'h3ff4a; 
        10'b1000111000: data <= 18'h3fffc; 
        10'b1000111001: data <= 18'h0004e; 
        10'b1000111010: data <= 18'h3ff34; 
        10'b1000111011: data <= 18'h3ffb6; 
        10'b1000111100: data <= 18'h3feb2; 
        10'b1000111101: data <= 18'h3ff8e; 
        10'b1000111110: data <= 18'h3ffad; 
        10'b1000111111: data <= 18'h00015; 
        10'b1001000000: data <= 18'h0013d; 
        10'b1001000001: data <= 18'h00072; 
        10'b1001000010: data <= 18'h3ff88; 
        10'b1001000011: data <= 18'h3fe43; 
        10'b1001000100: data <= 18'h3fdde; 
        10'b1001000101: data <= 18'h3fe06; 
        10'b1001000110: data <= 18'h3fe73; 
        10'b1001000111: data <= 18'h3ffa7; 
        10'b1001001000: data <= 18'h0002a; 
        10'b1001001001: data <= 18'h000fe; 
        10'b1001001010: data <= 18'h00065; 
        10'b1001001011: data <= 18'h00138; 
        10'b1001001100: data <= 18'h000de; 
        10'b1001001101: data <= 18'h00075; 
        10'b1001001110: data <= 18'h000b6; 
        10'b1001001111: data <= 18'h000d9; 
        10'b1001010000: data <= 18'h000ad; 
        10'b1001010001: data <= 18'h001d2; 
        10'b1001010010: data <= 18'h0017f; 
        10'b1001010011: data <= 18'h000b4; 
        10'b1001010100: data <= 18'h0001e; 
        10'b1001010101: data <= 18'h3ff7b; 
        10'b1001010110: data <= 18'h00006; 
        10'b1001010111: data <= 18'h3fef3; 
        10'b1001011000: data <= 18'h3fd9e; 
        10'b1001011001: data <= 18'h3fd47; 
        10'b1001011010: data <= 18'h3ffc1; 
        10'b1001011011: data <= 18'h000d1; 
        10'b1001011100: data <= 18'h0014e; 
        10'b1001011101: data <= 18'h0017d; 
        10'b1001011110: data <= 18'h00107; 
        10'b1001011111: data <= 18'h3fe46; 
        10'b1001100000: data <= 18'h3fe4d; 
        10'b1001100001: data <= 18'h3fe0f; 
        10'b1001100010: data <= 18'h3feaa; 
        10'b1001100011: data <= 18'h3ff3b; 
        10'b1001100100: data <= 18'h0002c; 
        10'b1001100101: data <= 18'h00087; 
        10'b1001100110: data <= 18'h0001b; 
        10'b1001100111: data <= 18'h00026; 
        10'b1001101000: data <= 18'h000ac; 
        10'b1001101001: data <= 18'h000b0; 
        10'b1001101010: data <= 18'h000c6; 
        10'b1001101011: data <= 18'h00029; 
        10'b1001101100: data <= 18'h00194; 
        10'b1001101101: data <= 18'h00385; 
        10'b1001101110: data <= 18'h003a5; 
        10'b1001101111: data <= 18'h00233; 
        10'b1001110000: data <= 18'h0004d; 
        10'b1001110001: data <= 18'h3ffc1; 
        10'b1001110010: data <= 18'h3ff2a; 
        10'b1001110011: data <= 18'h3fc87; 
        10'b1001110100: data <= 18'h3fa5c; 
        10'b1001110101: data <= 18'h3fbb0; 
        10'b1001110110: data <= 18'h00003; 
        10'b1001110111: data <= 18'h000d8; 
        10'b1001111000: data <= 18'h0033b; 
        10'b1001111001: data <= 18'h0054d; 
        10'b1001111010: data <= 18'h00252; 
        10'b1001111011: data <= 18'h0007c; 
        10'b1001111100: data <= 18'h3fece; 
        10'b1001111101: data <= 18'h3ff12; 
        10'b1001111110: data <= 18'h3ffeb; 
        10'b1001111111: data <= 18'h00028; 
        10'b1010000000: data <= 18'h00013; 
        10'b1010000001: data <= 18'h00084; 
        10'b1010000010: data <= 18'h0012c; 
        10'b1010000011: data <= 18'h00091; 
        10'b1010000100: data <= 18'h00117; 
        10'b1010000101: data <= 18'h000af; 
        10'b1010000110: data <= 18'h000e0; 
        10'b1010000111: data <= 18'h0007c; 
        10'b1010001000: data <= 18'h00168; 
        10'b1010001001: data <= 18'h00307; 
        10'b1010001010: data <= 18'h00339; 
        10'b1010001011: data <= 18'h0017b; 
        10'b1010001100: data <= 18'h00068; 
        10'b1010001101: data <= 18'h3ff40; 
        10'b1010001110: data <= 18'h3ff7d; 
        10'b1010001111: data <= 18'h3fe09; 
        10'b1010010000: data <= 18'h3fea1; 
        10'b1010010001: data <= 18'h3fec6; 
        10'b1010010010: data <= 18'h3fe5d; 
        10'b1010010011: data <= 18'h000a4; 
        10'b1010010100: data <= 18'h003c2; 
        10'b1010010101: data <= 18'h00489; 
        10'b1010010110: data <= 18'h00209; 
        10'b1010010111: data <= 18'h3ffa3; 
        10'b1010011000: data <= 18'h3ff22; 
        10'b1010011001: data <= 18'h3fea9; 
        10'b1010011010: data <= 18'h3ff8a; 
        10'b1010011011: data <= 18'h3ff93; 
        10'b1010011100: data <= 18'h00044; 
        10'b1010011101: data <= 18'h00022; 
        10'b1010011110: data <= 18'h00040; 
        10'b1010011111: data <= 18'h00020; 
        10'b1010100000: data <= 18'h00044; 
        10'b1010100001: data <= 18'h0002b; 
        10'b1010100010: data <= 18'h00071; 
        10'b1010100011: data <= 18'h00024; 
        10'b1010100100: data <= 18'h000b0; 
        10'b1010100101: data <= 18'h00157; 
        10'b1010100110: data <= 18'h00162; 
        10'b1010100111: data <= 18'h3ff8e; 
        10'b1010101000: data <= 18'h3fdff; 
        10'b1010101001: data <= 18'h3fdfc; 
        10'b1010101010: data <= 18'h3fc75; 
        10'b1010101011: data <= 18'h3fc9c; 
        10'b1010101100: data <= 18'h3fcf5; 
        10'b1010101101: data <= 18'h3fd65; 
        10'b1010101110: data <= 18'h3fd68; 
        10'b1010101111: data <= 18'h3fd66; 
        10'b1010110000: data <= 18'h3ff3f; 
        10'b1010110001: data <= 18'h00051; 
        10'b1010110010: data <= 18'h00093; 
        10'b1010110011: data <= 18'h000d5; 
        10'b1010110100: data <= 18'h000b2; 
        10'b1010110101: data <= 18'h0002b; 
        10'b1010110110: data <= 18'h0005d; 
        10'b1010110111: data <= 18'h000f7; 
        10'b1010111000: data <= 18'h0004b; 
        10'b1010111001: data <= 18'h0007a; 
        10'b1010111010: data <= 18'h000ea; 
        10'b1010111011: data <= 18'h0004d; 
        10'b1010111100: data <= 18'h0012f; 
        10'b1010111101: data <= 18'h00061; 
        10'b1010111110: data <= 18'h00074; 
        10'b1010111111: data <= 18'h000a4; 
        10'b1011000000: data <= 18'h000ea; 
        10'b1011000001: data <= 18'h000d6; 
        10'b1011000010: data <= 18'h00003; 
        10'b1011000011: data <= 18'h3ff7c; 
        10'b1011000100: data <= 18'h3ffcc; 
        10'b1011000101: data <= 18'h3ff86; 
        10'b1011000110: data <= 18'h3fe05; 
        10'b1011000111: data <= 18'h3fd97; 
        10'b1011001000: data <= 18'h3fe38; 
        10'b1011001001: data <= 18'h3fd80; 
        10'b1011001010: data <= 18'h3fe79; 
        10'b1011001011: data <= 18'h3fe11; 
        10'b1011001100: data <= 18'h3fee3; 
        10'b1011001101: data <= 18'h3ffcd; 
        10'b1011001110: data <= 18'h00063; 
        10'b1011001111: data <= 18'h000cd; 
        10'b1011010000: data <= 18'h00014; 
        10'b1011010001: data <= 18'h000ba; 
        10'b1011010010: data <= 18'h0006e; 
        10'b1011010011: data <= 18'h00109; 
        10'b1011010100: data <= 18'h00043; 
        10'b1011010101: data <= 18'h0004f; 
        10'b1011010110: data <= 18'h00071; 
        10'b1011010111: data <= 18'h00062; 
        10'b1011011000: data <= 18'h00070; 
        10'b1011011001: data <= 18'h000d7; 
        10'b1011011010: data <= 18'h000bf; 
        10'b1011011011: data <= 18'h0003a; 
        10'b1011011100: data <= 18'h000cf; 
        10'b1011011101: data <= 18'h00113; 
        10'b1011011110: data <= 18'h000ba; 
        10'b1011011111: data <= 18'h000ac; 
        10'b1011100000: data <= 18'h000f6; 
        10'b1011100001: data <= 18'h000d0; 
        10'b1011100010: data <= 18'h0001d; 
        10'b1011100011: data <= 18'h000a9; 
        10'b1011100100: data <= 18'h0009a; 
        10'b1011100101: data <= 18'h00059; 
        10'b1011100110: data <= 18'h3fffb; 
        10'b1011100111: data <= 18'h00050; 
        10'b1011101000: data <= 18'h000b4; 
        10'b1011101001: data <= 18'h00117; 
        10'b1011101010: data <= 18'h000ce; 
        10'b1011101011: data <= 18'h00021; 
        10'b1011101100: data <= 18'h000bf; 
        10'b1011101101: data <= 18'h000b4; 
        10'b1011101110: data <= 18'h000ab; 
        10'b1011101111: data <= 18'h00052; 
        10'b1011110000: data <= 18'h00048; 
        10'b1011110001: data <= 18'h000cf; 
        10'b1011110010: data <= 18'h0011c; 
        10'b1011110011: data <= 18'h000e6; 
        10'b1011110100: data <= 18'h000e7; 
        10'b1011110101: data <= 18'h00125; 
        10'b1011110110: data <= 18'h0002e; 
        10'b1011110111: data <= 18'h000a2; 
        10'b1011111000: data <= 18'h00133; 
        10'b1011111001: data <= 18'h000f4; 
        10'b1011111010: data <= 18'h00115; 
        10'b1011111011: data <= 18'h000ff; 
        10'b1011111100: data <= 18'h00115; 
        10'b1011111101: data <= 18'h00083; 
        10'b1011111110: data <= 18'h000f3; 
        10'b1011111111: data <= 18'h000fc; 
        10'b1100000000: data <= 18'h00019; 
        10'b1100000001: data <= 18'h00035; 
        10'b1100000010: data <= 18'h0012d; 
        10'b1100000011: data <= 18'h000c5; 
        10'b1100000100: data <= 18'h000b5; 
        10'b1100000101: data <= 18'h0001a; 
        10'b1100000110: data <= 18'h00083; 
        10'b1100000111: data <= 18'h0003a; 
        10'b1100001000: data <= 18'h00036; 
        10'b1100001001: data <= 18'h00063; 
        10'b1100001010: data <= 18'h000b2; 
        10'b1100001011: data <= 18'h00100; 
        10'b1100001100: data <= 18'h0011c; 
        10'b1100001101: data <= 18'h00115; 
        10'b1100001110: data <= 18'h00111; 
        10'b1100001111: data <= 18'h0005b; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 13) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 19'h001ff; 
        10'b0000000001: data <= 19'h000f4; 
        10'b0000000010: data <= 19'h00110; 
        10'b0000000011: data <= 19'h00070; 
        10'b0000000100: data <= 19'h001b1; 
        10'b0000000101: data <= 19'h001a5; 
        10'b0000000110: data <= 19'h001d1; 
        10'b0000000111: data <= 19'h00074; 
        10'b0000001000: data <= 19'h00196; 
        10'b0000001001: data <= 19'h0007c; 
        10'b0000001010: data <= 19'h00182; 
        10'b0000001011: data <= 19'h00137; 
        10'b0000001100: data <= 19'h001b2; 
        10'b0000001101: data <= 19'h00243; 
        10'b0000001110: data <= 19'h001fd; 
        10'b0000001111: data <= 19'h0015d; 
        10'b0000010000: data <= 19'h00162; 
        10'b0000010001: data <= 19'h0007d; 
        10'b0000010010: data <= 19'h00252; 
        10'b0000010011: data <= 19'h0024f; 
        10'b0000010100: data <= 19'h00152; 
        10'b0000010101: data <= 19'h001b1; 
        10'b0000010110: data <= 19'h0014f; 
        10'b0000010111: data <= 19'h00207; 
        10'b0000011000: data <= 19'h000c5; 
        10'b0000011001: data <= 19'h00224; 
        10'b0000011010: data <= 19'h0014f; 
        10'b0000011011: data <= 19'h001e3; 
        10'b0000011100: data <= 19'h0003f; 
        10'b0000011101: data <= 19'h00201; 
        10'b0000011110: data <= 19'h00097; 
        10'b0000011111: data <= 19'h0016d; 
        10'b0000100000: data <= 19'h00146; 
        10'b0000100001: data <= 19'h00081; 
        10'b0000100010: data <= 19'h000b6; 
        10'b0000100011: data <= 19'h001e2; 
        10'b0000100100: data <= 19'h001cf; 
        10'b0000100101: data <= 19'h00178; 
        10'b0000100110: data <= 19'h00174; 
        10'b0000100111: data <= 19'h00112; 
        10'b0000101000: data <= 19'h001bb; 
        10'b0000101001: data <= 19'h001f4; 
        10'b0000101010: data <= 19'h00286; 
        10'b0000101011: data <= 19'h00142; 
        10'b0000101100: data <= 19'h00104; 
        10'b0000101101: data <= 19'h00207; 
        10'b0000101110: data <= 19'h0015d; 
        10'b0000101111: data <= 19'h000ed; 
        10'b0000110000: data <= 19'h00233; 
        10'b0000110001: data <= 19'h0021d; 
        10'b0000110010: data <= 19'h000de; 
        10'b0000110011: data <= 19'h00245; 
        10'b0000110100: data <= 19'h0026e; 
        10'b0000110101: data <= 19'h00149; 
        10'b0000110110: data <= 19'h00212; 
        10'b0000110111: data <= 19'h001aa; 
        10'b0000111000: data <= 19'h0020b; 
        10'b0000111001: data <= 19'h00189; 
        10'b0000111010: data <= 19'h00272; 
        10'b0000111011: data <= 19'h00079; 
        10'b0000111100: data <= 19'h00075; 
        10'b0000111101: data <= 19'h0019c; 
        10'b0000111110: data <= 19'h00131; 
        10'b0000111111: data <= 19'h00125; 
        10'b0001000000: data <= 19'h000c5; 
        10'b0001000001: data <= 19'h00159; 
        10'b0001000010: data <= 19'h00009; 
        10'b0001000011: data <= 19'h000ad; 
        10'b0001000100: data <= 19'h00016; 
        10'b0001000101: data <= 19'h00098; 
        10'b0001000110: data <= 19'h0013e; 
        10'b0001000111: data <= 19'h001fe; 
        10'b0001001000: data <= 19'h00182; 
        10'b0001001001: data <= 19'h00000; 
        10'b0001001010: data <= 19'h0017d; 
        10'b0001001011: data <= 19'h000e5; 
        10'b0001001100: data <= 19'h001f5; 
        10'b0001001101: data <= 19'h000da; 
        10'b0001001110: data <= 19'h00228; 
        10'b0001001111: data <= 19'h00192; 
        10'b0001010000: data <= 19'h001b0; 
        10'b0001010001: data <= 19'h0004a; 
        10'b0001010010: data <= 19'h001d6; 
        10'b0001010011: data <= 19'h001e1; 
        10'b0001010100: data <= 19'h000ba; 
        10'b0001010101: data <= 19'h000d1; 
        10'b0001010110: data <= 19'h00160; 
        10'b0001010111: data <= 19'h00121; 
        10'b0001011000: data <= 19'h0024c; 
        10'b0001011001: data <= 19'h00136; 
        10'b0001011010: data <= 19'h00044; 
        10'b0001011011: data <= 19'h00240; 
        10'b0001011100: data <= 19'h7ffc1; 
        10'b0001011101: data <= 19'h7ff8c; 
        10'b0001011110: data <= 19'h7ff90; 
        10'b0001011111: data <= 19'h7fec0; 
        10'b0001100000: data <= 19'h7ff8f; 
        10'b0001100001: data <= 19'h0002b; 
        10'b0001100010: data <= 19'h000f0; 
        10'b0001100011: data <= 19'h001e0; 
        10'b0001100100: data <= 19'h7ff12; 
        10'b0001100101: data <= 19'h7ffa9; 
        10'b0001100110: data <= 19'h7fff4; 
        10'b0001100111: data <= 19'h7fe8e; 
        10'b0001101000: data <= 19'h7ffda; 
        10'b0001101001: data <= 19'h00098; 
        10'b0001101010: data <= 19'h0017f; 
        10'b0001101011: data <= 19'h00176; 
        10'b0001101100: data <= 19'h7ffbb; 
        10'b0001101101: data <= 19'h00213; 
        10'b0001101110: data <= 19'h000c8; 
        10'b0001101111: data <= 19'h00231; 
        10'b0001110000: data <= 19'h001b0; 
        10'b0001110001: data <= 19'h00106; 
        10'b0001110010: data <= 19'h00253; 
        10'b0001110011: data <= 19'h0024e; 
        10'b0001110100: data <= 19'h00042; 
        10'b0001110101: data <= 19'h00075; 
        10'b0001110110: data <= 19'h00207; 
        10'b0001110111: data <= 19'h0014b; 
        10'b0001111000: data <= 19'h0007d; 
        10'b0001111001: data <= 19'h7fde1; 
        10'b0001111010: data <= 19'h00032; 
        10'b0001111011: data <= 19'h000be; 
        10'b0001111100: data <= 19'h00128; 
        10'b0001111101: data <= 19'h00210; 
        10'b0001111110: data <= 19'h0026c; 
        10'b0001111111: data <= 19'h004f3; 
        10'b0010000000: data <= 19'h0015a; 
        10'b0010000001: data <= 19'h7fef6; 
        10'b0010000010: data <= 19'h7fede; 
        10'b0010000011: data <= 19'h000c5; 
        10'b0010000100: data <= 19'h002bd; 
        10'b0010000101: data <= 19'h00312; 
        10'b0010000110: data <= 19'h0030e; 
        10'b0010000111: data <= 19'h00394; 
        10'b0010001000: data <= 19'h001df; 
        10'b0010001001: data <= 19'h000e3; 
        10'b0010001010: data <= 19'h000c6; 
        10'b0010001011: data <= 19'h000da; 
        10'b0010001100: data <= 19'h0004e; 
        10'b0010001101: data <= 19'h001ff; 
        10'b0010001110: data <= 19'h00064; 
        10'b0010001111: data <= 19'h00168; 
        10'b0010010000: data <= 19'h0005a; 
        10'b0010010001: data <= 19'h00159; 
        10'b0010010010: data <= 19'h00068; 
        10'b0010010011: data <= 19'h7ff7a; 
        10'b0010010100: data <= 19'h7fb8b; 
        10'b0010010101: data <= 19'h7fb82; 
        10'b0010010110: data <= 19'h7fdf1; 
        10'b0010010111: data <= 19'h00007; 
        10'b0010011000: data <= 19'h001b0; 
        10'b0010011001: data <= 19'h001e6; 
        10'b0010011010: data <= 19'h0034d; 
        10'b0010011011: data <= 19'h00291; 
        10'b0010011100: data <= 19'h00184; 
        10'b0010011101: data <= 19'h7fd81; 
        10'b0010011110: data <= 19'h7ffc0; 
        10'b0010011111: data <= 19'h00086; 
        10'b0010100000: data <= 19'h00270; 
        10'b0010100001: data <= 19'h003ed; 
        10'b0010100010: data <= 19'h00689; 
        10'b0010100011: data <= 19'h00414; 
        10'b0010100100: data <= 19'h00357; 
        10'b0010100101: data <= 19'h7ff24; 
        10'b0010100110: data <= 19'h000ec; 
        10'b0010100111: data <= 19'h00083; 
        10'b0010101000: data <= 19'h0006d; 
        10'b0010101001: data <= 19'h00173; 
        10'b0010101010: data <= 19'h00044; 
        10'b0010101011: data <= 19'h00121; 
        10'b0010101100: data <= 19'h00044; 
        10'b0010101101: data <= 19'h7ff56; 
        10'b0010101110: data <= 19'h7fd8c; 
        10'b0010101111: data <= 19'h7fd94; 
        10'b0010110000: data <= 19'h7fa6e; 
        10'b0010110001: data <= 19'h7f945; 
        10'b0010110010: data <= 19'h7fbc9; 
        10'b0010110011: data <= 19'h7ff03; 
        10'b0010110100: data <= 19'h7fef8; 
        10'b0010110101: data <= 19'h7fde2; 
        10'b0010110110: data <= 19'h7ff07; 
        10'b0010110111: data <= 19'h7fb2b; 
        10'b0010111000: data <= 19'h7face; 
        10'b0010111001: data <= 19'h7fac3; 
        10'b0010111010: data <= 19'h7fdcf; 
        10'b0010111011: data <= 19'h7fe61; 
        10'b0010111100: data <= 19'h00273; 
        10'b0010111101: data <= 19'h00409; 
        10'b0010111110: data <= 19'h003be; 
        10'b0010111111: data <= 19'h00326; 
        10'b0011000000: data <= 19'h000d2; 
        10'b0011000001: data <= 19'h7ff55; 
        10'b0011000010: data <= 19'h0000e; 
        10'b0011000011: data <= 19'h0012e; 
        10'b0011000100: data <= 19'h000f4; 
        10'b0011000101: data <= 19'h0008a; 
        10'b0011000110: data <= 19'h000ab; 
        10'b0011000111: data <= 19'h00026; 
        10'b0011001000: data <= 19'h00195; 
        10'b0011001001: data <= 19'h7ffa9; 
        10'b0011001010: data <= 19'h7fda6; 
        10'b0011001011: data <= 19'h7fb31; 
        10'b0011001100: data <= 19'h7f87c; 
        10'b0011001101: data <= 19'h7f66d; 
        10'b0011001110: data <= 19'h7f980; 
        10'b0011001111: data <= 19'h7fd29; 
        10'b0011010000: data <= 19'h7fd66; 
        10'b0011010001: data <= 19'h7fc42; 
        10'b0011010010: data <= 19'h7fb60; 
        10'b0011010011: data <= 19'h7f8cf; 
        10'b0011010100: data <= 19'h7f9b8; 
        10'b0011010101: data <= 19'h7fa1b; 
        10'b0011010110: data <= 19'h7fab0; 
        10'b0011010111: data <= 19'h7ffd2; 
        10'b0011011000: data <= 19'h0011d; 
        10'b0011011001: data <= 19'h000b1; 
        10'b0011011010: data <= 19'h000a9; 
        10'b0011011011: data <= 19'h7fdfa; 
        10'b0011011100: data <= 19'h7fd3e; 
        10'b0011011101: data <= 19'h7fee6; 
        10'b0011011110: data <= 19'h000e6; 
        10'b0011011111: data <= 19'h0010c; 
        10'b0011100000: data <= 19'h00129; 
        10'b0011100001: data <= 19'h000fb; 
        10'b0011100010: data <= 19'h000f7; 
        10'b0011100011: data <= 19'h0020c; 
        10'b0011100100: data <= 19'h000a7; 
        10'b0011100101: data <= 19'h7ffef; 
        10'b0011100110: data <= 19'h7fd34; 
        10'b0011100111: data <= 19'h7fbc3; 
        10'b0011101000: data <= 19'h7f73d; 
        10'b0011101001: data <= 19'h7f67d; 
        10'b0011101010: data <= 19'h7f6f2; 
        10'b0011101011: data <= 19'h7fb21; 
        10'b0011101100: data <= 19'h7fdc3; 
        10'b0011101101: data <= 19'h7fd40; 
        10'b0011101110: data <= 19'h7fdc1; 
        10'b0011101111: data <= 19'h000fc; 
        10'b0011110000: data <= 19'h7fc04; 
        10'b0011110001: data <= 19'h7fea6; 
        10'b0011110010: data <= 19'h7ffc6; 
        10'b0011110011: data <= 19'h00084; 
        10'b0011110100: data <= 19'h7fd01; 
        10'b0011110101: data <= 19'h7fd1a; 
        10'b0011110110: data <= 19'h7fb5c; 
        10'b0011110111: data <= 19'h7f9e9; 
        10'b0011111000: data <= 19'h7fb28; 
        10'b0011111001: data <= 19'h7fed0; 
        10'b0011111010: data <= 19'h001ce; 
        10'b0011111011: data <= 19'h00260; 
        10'b0011111100: data <= 19'h00266; 
        10'b0011111101: data <= 19'h0008e; 
        10'b0011111110: data <= 19'h000fc; 
        10'b0011111111: data <= 19'h000d7; 
        10'b0100000000: data <= 19'h7ffd9; 
        10'b0100000001: data <= 19'h7ffbc; 
        10'b0100000010: data <= 19'h7fc71; 
        10'b0100000011: data <= 19'h7fca1; 
        10'b0100000100: data <= 19'h7f9f8; 
        10'b0100000101: data <= 19'h7f6cf; 
        10'b0100000110: data <= 19'h7f794; 
        10'b0100000111: data <= 19'h7fcac; 
        10'b0100001000: data <= 19'h7fd84; 
        10'b0100001001: data <= 19'h001e4; 
        10'b0100001010: data <= 19'h005f3; 
        10'b0100001011: data <= 19'h00885; 
        10'b0100001100: data <= 19'h00328; 
        10'b0100001101: data <= 19'h7ffc8; 
        10'b0100001110: data <= 19'h7fe94; 
        10'b0100001111: data <= 19'h7fa39; 
        10'b0100010000: data <= 19'h7f8e5; 
        10'b0100010001: data <= 19'h7f8fd; 
        10'b0100010010: data <= 19'h7f72b; 
        10'b0100010011: data <= 19'h7f859; 
        10'b0100010100: data <= 19'h7fbe5; 
        10'b0100010101: data <= 19'h0007a; 
        10'b0100010110: data <= 19'h001fb; 
        10'b0100010111: data <= 19'h00170; 
        10'b0100011000: data <= 19'h00230; 
        10'b0100011001: data <= 19'h0026c; 
        10'b0100011010: data <= 19'h00201; 
        10'b0100011011: data <= 19'h00043; 
        10'b0100011100: data <= 19'h001a3; 
        10'b0100011101: data <= 19'h7fe1b; 
        10'b0100011110: data <= 19'h7fca2; 
        10'b0100011111: data <= 19'h7fe70; 
        10'b0100100000: data <= 19'h7fb53; 
        10'b0100100001: data <= 19'h7fb42; 
        10'b0100100010: data <= 19'h7fc89; 
        10'b0100100011: data <= 19'h7fdaf; 
        10'b0100100100: data <= 19'h7fe71; 
        10'b0100100101: data <= 19'h004c0; 
        10'b0100100110: data <= 19'h00f60; 
        10'b0100100111: data <= 19'h0103b; 
        10'b0100101000: data <= 19'h007b5; 
        10'b0100101001: data <= 19'h7ffd5; 
        10'b0100101010: data <= 19'h7fb63; 
        10'b0100101011: data <= 19'h7fa70; 
        10'b0100101100: data <= 19'h7f945; 
        10'b0100101101: data <= 19'h7f9ee; 
        10'b0100101110: data <= 19'h7fa48; 
        10'b0100101111: data <= 19'h7fc73; 
        10'b0100110000: data <= 19'h7fecf; 
        10'b0100110001: data <= 19'h7ffcb; 
        10'b0100110010: data <= 19'h0020f; 
        10'b0100110011: data <= 19'h000d8; 
        10'b0100110100: data <= 19'h0006a; 
        10'b0100110101: data <= 19'h0005f; 
        10'b0100110110: data <= 19'h001aa; 
        10'b0100110111: data <= 19'h001c6; 
        10'b0100111000: data <= 19'h00002; 
        10'b0100111001: data <= 19'h7ff77; 
        10'b0100111010: data <= 19'h7ffb8; 
        10'b0100111011: data <= 19'h7fd13; 
        10'b0100111100: data <= 19'h7fe1c; 
        10'b0100111101: data <= 19'h7fd15; 
        10'b0100111110: data <= 19'h7fbb5; 
        10'b0100111111: data <= 19'h7f984; 
        10'b0101000000: data <= 19'h7ff42; 
        10'b0101000001: data <= 19'h00820; 
        10'b0101000010: data <= 19'h01289; 
        10'b0101000011: data <= 19'h013a3; 
        10'b0101000100: data <= 19'h00746; 
        10'b0101000101: data <= 19'h7fe69; 
        10'b0101000110: data <= 19'h7fe89; 
        10'b0101000111: data <= 19'h7fc21; 
        10'b0101001000: data <= 19'h7fbe8; 
        10'b0101001001: data <= 19'h7fc32; 
        10'b0101001010: data <= 19'h7fc7b; 
        10'b0101001011: data <= 19'h7fe5a; 
        10'b0101001100: data <= 19'h7ff4d; 
        10'b0101001101: data <= 19'h001a1; 
        10'b0101001110: data <= 19'h00249; 
        10'b0101001111: data <= 19'h0019c; 
        10'b0101010000: data <= 19'h00041; 
        10'b0101010001: data <= 19'h00230; 
        10'b0101010010: data <= 19'h0010d; 
        10'b0101010011: data <= 19'h000b6; 
        10'b0101010100: data <= 19'h0023d; 
        10'b0101010101: data <= 19'h7ff92; 
        10'b0101010110: data <= 19'h7ff51; 
        10'b0101010111: data <= 19'h7ff08; 
        10'b0101011000: data <= 19'h7fd37; 
        10'b0101011001: data <= 19'h7fc59; 
        10'b0101011010: data <= 19'h7f843; 
        10'b0101011011: data <= 19'h7f525; 
        10'b0101011100: data <= 19'h7ffa7; 
        10'b0101011101: data <= 19'h0083f; 
        10'b0101011110: data <= 19'h015d1; 
        10'b0101011111: data <= 19'h00f22; 
        10'b0101100000: data <= 19'h002ff; 
        10'b0101100001: data <= 19'h00196; 
        10'b0101100010: data <= 19'h7ff11; 
        10'b0101100011: data <= 19'h7fb94; 
        10'b0101100100: data <= 19'h7fd36; 
        10'b0101100101: data <= 19'h7fea5; 
        10'b0101100110: data <= 19'h7ff3d; 
        10'b0101100111: data <= 19'h7ff10; 
        10'b0101101000: data <= 19'h00024; 
        10'b0101101001: data <= 19'h00239; 
        10'b0101101010: data <= 19'h00055; 
        10'b0101101011: data <= 19'h00190; 
        10'b0101101100: data <= 19'h00039; 
        10'b0101101101: data <= 19'h0017c; 
        10'b0101101110: data <= 19'h00163; 
        10'b0101101111: data <= 19'h0017b; 
        10'b0101110000: data <= 19'h00277; 
        10'b0101110001: data <= 19'h00004; 
        10'b0101110010: data <= 19'h00035; 
        10'b0101110011: data <= 19'h7fee5; 
        10'b0101110100: data <= 19'h7fe83; 
        10'b0101110101: data <= 19'h7f9ea; 
        10'b0101110110: data <= 19'h7f316; 
        10'b0101110111: data <= 19'h7f2e7; 
        10'b0101111000: data <= 19'h00005; 
        10'b0101111001: data <= 19'h006e1; 
        10'b0101111010: data <= 19'h011fa; 
        10'b0101111011: data <= 19'h00a29; 
        10'b0101111100: data <= 19'h002b0; 
        10'b0101111101: data <= 19'h0014e; 
        10'b0101111110: data <= 19'h7fbe6; 
        10'b0101111111: data <= 19'h7fa0a; 
        10'b0110000000: data <= 19'h7fdd6; 
        10'b0110000001: data <= 19'h7ff3d; 
        10'b0110000010: data <= 19'h7ff35; 
        10'b0110000011: data <= 19'h7ffb7; 
        10'b0110000100: data <= 19'h00101; 
        10'b0110000101: data <= 19'h00181; 
        10'b0110000110: data <= 19'h0022b; 
        10'b0110000111: data <= 19'h00167; 
        10'b0110001000: data <= 19'h00118; 
        10'b0110001001: data <= 19'h00257; 
        10'b0110001010: data <= 19'h00151; 
        10'b0110001011: data <= 19'h001e0; 
        10'b0110001100: data <= 19'h001e2; 
        10'b0110001101: data <= 19'h7fffe; 
        10'b0110001110: data <= 19'h00052; 
        10'b0110001111: data <= 19'h7ff48; 
        10'b0110010000: data <= 19'h7fbf9; 
        10'b0110010001: data <= 19'h7f916; 
        10'b0110010010: data <= 19'h7f322; 
        10'b0110010011: data <= 19'h7f63c; 
        10'b0110010100: data <= 19'h7ffc8; 
        10'b0110010101: data <= 19'h006fb; 
        10'b0110010110: data <= 19'h00f55; 
        10'b0110010111: data <= 19'h009e0; 
        10'b0110011000: data <= 19'h002f4; 
        10'b0110011001: data <= 19'h7fa85; 
        10'b0110011010: data <= 19'h7f894; 
        10'b0110011011: data <= 19'h7fa5d; 
        10'b0110011100: data <= 19'h7fcaa; 
        10'b0110011101: data <= 19'h7ff09; 
        10'b0110011110: data <= 19'h7fef4; 
        10'b0110011111: data <= 19'h7ff49; 
        10'b0110100000: data <= 19'h001ac; 
        10'b0110100001: data <= 19'h00042; 
        10'b0110100010: data <= 19'h00076; 
        10'b0110100011: data <= 19'h00155; 
        10'b0110100100: data <= 19'h0027b; 
        10'b0110100101: data <= 19'h00068; 
        10'b0110100110: data <= 19'h00197; 
        10'b0110100111: data <= 19'h00102; 
        10'b0110101000: data <= 19'h00092; 
        10'b0110101001: data <= 19'h00172; 
        10'b0110101010: data <= 19'h7fe98; 
        10'b0110101011: data <= 19'h7fe66; 
        10'b0110101100: data <= 19'h7fd76; 
        10'b0110101101: data <= 19'h7f870; 
        10'b0110101110: data <= 19'h7f785; 
        10'b0110101111: data <= 19'h7fddd; 
        10'b0110110000: data <= 19'h0031c; 
        10'b0110110001: data <= 19'h009d1; 
        10'b0110110010: data <= 19'h01069; 
        10'b0110110011: data <= 19'h005ce; 
        10'b0110110100: data <= 19'h00110; 
        10'b0110110101: data <= 19'h7f5ac; 
        10'b0110110110: data <= 19'h7f6d9; 
        10'b0110110111: data <= 19'h7fa66; 
        10'b0110111000: data <= 19'h7fca1; 
        10'b0110111001: data <= 19'h7fd94; 
        10'b0110111010: data <= 19'h7ff64; 
        10'b0110111011: data <= 19'h0002f; 
        10'b0110111100: data <= 19'h000e0; 
        10'b0110111101: data <= 19'h0011f; 
        10'b0110111110: data <= 19'h0024f; 
        10'b0110111111: data <= 19'h00063; 
        10'b0111000000: data <= 19'h00267; 
        10'b0111000001: data <= 19'h0012d; 
        10'b0111000010: data <= 19'h00232; 
        10'b0111000011: data <= 19'h00156; 
        10'b0111000100: data <= 19'h000b6; 
        10'b0111000101: data <= 19'h7ff06; 
        10'b0111000110: data <= 19'h7fdc5; 
        10'b0111000111: data <= 19'h7fd9b; 
        10'b0111001000: data <= 19'h7fa24; 
        10'b0111001001: data <= 19'h7fc7e; 
        10'b0111001010: data <= 19'h7fd35; 
        10'b0111001011: data <= 19'h7fe73; 
        10'b0111001100: data <= 19'h7ff9b; 
        10'b0111001101: data <= 19'h00ce9; 
        10'b0111001110: data <= 19'h00f7d; 
        10'b0111001111: data <= 19'h000e3; 
        10'b0111010000: data <= 19'h7fb34; 
        10'b0111010001: data <= 19'h7f4d3; 
        10'b0111010010: data <= 19'h7f6c1; 
        10'b0111010011: data <= 19'h7fa0c; 
        10'b0111010100: data <= 19'h7fb7b; 
        10'b0111010101: data <= 19'h7fe12; 
        10'b0111010110: data <= 19'h7fe0b; 
        10'b0111010111: data <= 19'h00006; 
        10'b0111011000: data <= 19'h7ff23; 
        10'b0111011001: data <= 19'h00022; 
        10'b0111011010: data <= 19'h00097; 
        10'b0111011011: data <= 19'h0013f; 
        10'b0111011100: data <= 19'h000ff; 
        10'b0111011101: data <= 19'h0025f; 
        10'b0111011110: data <= 19'h00087; 
        10'b0111011111: data <= 19'h00257; 
        10'b0111100000: data <= 19'h001bb; 
        10'b0111100001: data <= 19'h7fea4; 
        10'b0111100010: data <= 19'h7fb18; 
        10'b0111100011: data <= 19'h7fab0; 
        10'b0111100100: data <= 19'h7fc32; 
        10'b0111100101: data <= 19'h7fd91; 
        10'b0111100110: data <= 19'h001bf; 
        10'b0111100111: data <= 19'h00005; 
        10'b0111101000: data <= 19'h00438; 
        10'b0111101001: data <= 19'h00ec9; 
        10'b0111101010: data <= 19'h00cae; 
        10'b0111101011: data <= 19'h7fd6d; 
        10'b0111101100: data <= 19'h7f730; 
        10'b0111101101: data <= 19'h7f4c9; 
        10'b0111101110: data <= 19'h7f6d0; 
        10'b0111101111: data <= 19'h7fa31; 
        10'b0111110000: data <= 19'h7fdd1; 
        10'b0111110001: data <= 19'h7fee7; 
        10'b0111110010: data <= 19'h7ff36; 
        10'b0111110011: data <= 19'h7fef2; 
        10'b0111110100: data <= 19'h7fe31; 
        10'b0111110101: data <= 19'h00085; 
        10'b0111110110: data <= 19'h00162; 
        10'b0111110111: data <= 19'h0019e; 
        10'b0111111000: data <= 19'h00177; 
        10'b0111111001: data <= 19'h0015a; 
        10'b0111111010: data <= 19'h000d5; 
        10'b0111111011: data <= 19'h001f4; 
        10'b0111111100: data <= 19'h00115; 
        10'b0111111101: data <= 19'h7fe10; 
        10'b0111111110: data <= 19'h7fac4; 
        10'b0111111111: data <= 19'h7facf; 
        10'b1000000000: data <= 19'h7fe0e; 
        10'b1000000001: data <= 19'h001fd; 
        10'b1000000010: data <= 19'h001a4; 
        10'b1000000011: data <= 19'h002a1; 
        10'b1000000100: data <= 19'h006dc; 
        10'b1000000101: data <= 19'h00b0c; 
        10'b1000000110: data <= 19'h007a3; 
        10'b1000000111: data <= 19'h7fafb; 
        10'b1000001000: data <= 19'h7f7c0; 
        10'b1000001001: data <= 19'h7f8ef; 
        10'b1000001010: data <= 19'h7f9f7; 
        10'b1000001011: data <= 19'h7fbf5; 
        10'b1000001100: data <= 19'h7fe03; 
        10'b1000001101: data <= 19'h7fca3; 
        10'b1000001110: data <= 19'h7fe82; 
        10'b1000001111: data <= 19'h7fdb6; 
        10'b1000010000: data <= 19'h7fe9a; 
        10'b1000010001: data <= 19'h00144; 
        10'b1000010010: data <= 19'h00233; 
        10'b1000010011: data <= 19'h0023f; 
        10'b1000010100: data <= 19'h0024f; 
        10'b1000010101: data <= 19'h001a0; 
        10'b1000010110: data <= 19'h001b1; 
        10'b1000010111: data <= 19'h001e0; 
        10'b1000011000: data <= 19'h00038; 
        10'b1000011001: data <= 19'h7fd18; 
        10'b1000011010: data <= 19'h7f982; 
        10'b1000011011: data <= 19'h7fb9e; 
        10'b1000011100: data <= 19'h7fe36; 
        10'b1000011101: data <= 19'h00108; 
        10'b1000011110: data <= 19'h00084; 
        10'b1000011111: data <= 19'h0005c; 
        10'b1000100000: data <= 19'h000e9; 
        10'b1000100001: data <= 19'h00516; 
        10'b1000100010: data <= 19'h0011f; 
        10'b1000100011: data <= 19'h7fbd9; 
        10'b1000100100: data <= 19'h7fc8b; 
        10'b1000100101: data <= 19'h7fcfd; 
        10'b1000100110: data <= 19'h7fc38; 
        10'b1000100111: data <= 19'h7fd11; 
        10'b1000101000: data <= 19'h7fbb5; 
        10'b1000101001: data <= 19'h7fc6d; 
        10'b1000101010: data <= 19'h7fdd8; 
        10'b1000101011: data <= 19'h7fe19; 
        10'b1000101100: data <= 19'h0001b; 
        10'b1000101101: data <= 19'h000ba; 
        10'b1000101110: data <= 19'h000cd; 
        10'b1000101111: data <= 19'h00052; 
        10'b1000110000: data <= 19'h0005e; 
        10'b1000110001: data <= 19'h0026d; 
        10'b1000110010: data <= 19'h0014f; 
        10'b1000110011: data <= 19'h000d7; 
        10'b1000110100: data <= 19'h7ff59; 
        10'b1000110101: data <= 19'h7fdee; 
        10'b1000110110: data <= 19'h7ff9d; 
        10'b1000110111: data <= 19'h7fe94; 
        10'b1000111000: data <= 19'h7fff7; 
        10'b1000111001: data <= 19'h0009c; 
        10'b1000111010: data <= 19'h7fe67; 
        10'b1000111011: data <= 19'h7ff6d; 
        10'b1000111100: data <= 19'h7fd65; 
        10'b1000111101: data <= 19'h7ff1c; 
        10'b1000111110: data <= 19'h7ff5a; 
        10'b1000111111: data <= 19'h0002a; 
        10'b1001000000: data <= 19'h00279; 
        10'b1001000001: data <= 19'h000e4; 
        10'b1001000010: data <= 19'h7ff11; 
        10'b1001000011: data <= 19'h7fc87; 
        10'b1001000100: data <= 19'h7fbbb; 
        10'b1001000101: data <= 19'h7fc0c; 
        10'b1001000110: data <= 19'h7fce5; 
        10'b1001000111: data <= 19'h7ff4d; 
        10'b1001001000: data <= 19'h00054; 
        10'b1001001001: data <= 19'h001fb; 
        10'b1001001010: data <= 19'h000cb; 
        10'b1001001011: data <= 19'h00271; 
        10'b1001001100: data <= 19'h001bc; 
        10'b1001001101: data <= 19'h000ea; 
        10'b1001001110: data <= 19'h0016b; 
        10'b1001001111: data <= 19'h001b3; 
        10'b1001010000: data <= 19'h00159; 
        10'b1001010001: data <= 19'h003a4; 
        10'b1001010010: data <= 19'h002fe; 
        10'b1001010011: data <= 19'h00168; 
        10'b1001010100: data <= 19'h0003c; 
        10'b1001010101: data <= 19'h7fef7; 
        10'b1001010110: data <= 19'h0000b; 
        10'b1001010111: data <= 19'h7fde7; 
        10'b1001011000: data <= 19'h7fb3b; 
        10'b1001011001: data <= 19'h7fa8f; 
        10'b1001011010: data <= 19'h7ff83; 
        10'b1001011011: data <= 19'h001a3; 
        10'b1001011100: data <= 19'h0029d; 
        10'b1001011101: data <= 19'h002f9; 
        10'b1001011110: data <= 19'h0020d; 
        10'b1001011111: data <= 19'h7fc8b; 
        10'b1001100000: data <= 19'h7fc9a; 
        10'b1001100001: data <= 19'h7fc1f; 
        10'b1001100010: data <= 19'h7fd55; 
        10'b1001100011: data <= 19'h7fe76; 
        10'b1001100100: data <= 19'h00058; 
        10'b1001100101: data <= 19'h0010e; 
        10'b1001100110: data <= 19'h00035; 
        10'b1001100111: data <= 19'h0004d; 
        10'b1001101000: data <= 19'h00159; 
        10'b1001101001: data <= 19'h00160; 
        10'b1001101010: data <= 19'h0018d; 
        10'b1001101011: data <= 19'h00051; 
        10'b1001101100: data <= 19'h00327; 
        10'b1001101101: data <= 19'h0070a; 
        10'b1001101110: data <= 19'h0074a; 
        10'b1001101111: data <= 19'h00466; 
        10'b1001110000: data <= 19'h00099; 
        10'b1001110001: data <= 19'h7ff83; 
        10'b1001110010: data <= 19'h7fe54; 
        10'b1001110011: data <= 19'h7f90d; 
        10'b1001110100: data <= 19'h7f4b9; 
        10'b1001110101: data <= 19'h7f760; 
        10'b1001110110: data <= 19'h00007; 
        10'b1001110111: data <= 19'h001b1; 
        10'b1001111000: data <= 19'h00677; 
        10'b1001111001: data <= 19'h00a99; 
        10'b1001111010: data <= 19'h004a3; 
        10'b1001111011: data <= 19'h000f7; 
        10'b1001111100: data <= 19'h7fd9d; 
        10'b1001111101: data <= 19'h7fe24; 
        10'b1001111110: data <= 19'h7ffd6; 
        10'b1001111111: data <= 19'h00050; 
        10'b1010000000: data <= 19'h00026; 
        10'b1010000001: data <= 19'h00107; 
        10'b1010000010: data <= 19'h00258; 
        10'b1010000011: data <= 19'h00121; 
        10'b1010000100: data <= 19'h0022f; 
        10'b1010000101: data <= 19'h0015d; 
        10'b1010000110: data <= 19'h001bf; 
        10'b1010000111: data <= 19'h000f9; 
        10'b1010001000: data <= 19'h002d1; 
        10'b1010001001: data <= 19'h0060d; 
        10'b1010001010: data <= 19'h00673; 
        10'b1010001011: data <= 19'h002f6; 
        10'b1010001100: data <= 19'h000d1; 
        10'b1010001101: data <= 19'h7fe80; 
        10'b1010001110: data <= 19'h7fefa; 
        10'b1010001111: data <= 19'h7fc12; 
        10'b1010010000: data <= 19'h7fd42; 
        10'b1010010001: data <= 19'h7fd8d; 
        10'b1010010010: data <= 19'h7fcba; 
        10'b1010010011: data <= 19'h00148; 
        10'b1010010100: data <= 19'h00785; 
        10'b1010010101: data <= 19'h00911; 
        10'b1010010110: data <= 19'h00413; 
        10'b1010010111: data <= 19'h7ff47; 
        10'b1010011000: data <= 19'h7fe45; 
        10'b1010011001: data <= 19'h7fd52; 
        10'b1010011010: data <= 19'h7ff14; 
        10'b1010011011: data <= 19'h7ff26; 
        10'b1010011100: data <= 19'h00088; 
        10'b1010011101: data <= 19'h00045; 
        10'b1010011110: data <= 19'h00080; 
        10'b1010011111: data <= 19'h0003f; 
        10'b1010100000: data <= 19'h00088; 
        10'b1010100001: data <= 19'h00056; 
        10'b1010100010: data <= 19'h000e2; 
        10'b1010100011: data <= 19'h00047; 
        10'b1010100100: data <= 19'h00160; 
        10'b1010100101: data <= 19'h002ad; 
        10'b1010100110: data <= 19'h002c3; 
        10'b1010100111: data <= 19'h7ff1c; 
        10'b1010101000: data <= 19'h7fbfd; 
        10'b1010101001: data <= 19'h7fbf8; 
        10'b1010101010: data <= 19'h7f8ea; 
        10'b1010101011: data <= 19'h7f938; 
        10'b1010101100: data <= 19'h7f9ea; 
        10'b1010101101: data <= 19'h7fac9; 
        10'b1010101110: data <= 19'h7facf; 
        10'b1010101111: data <= 19'h7facc; 
        10'b1010110000: data <= 19'h7fe7f; 
        10'b1010110001: data <= 19'h000a1; 
        10'b1010110010: data <= 19'h00126; 
        10'b1010110011: data <= 19'h001aa; 
        10'b1010110100: data <= 19'h00165; 
        10'b1010110101: data <= 19'h00056; 
        10'b1010110110: data <= 19'h000b9; 
        10'b1010110111: data <= 19'h001ee; 
        10'b1010111000: data <= 19'h00096; 
        10'b1010111001: data <= 19'h000f3; 
        10'b1010111010: data <= 19'h001d5; 
        10'b1010111011: data <= 19'h0009b; 
        10'b1010111100: data <= 19'h0025f; 
        10'b1010111101: data <= 19'h000c1; 
        10'b1010111110: data <= 19'h000e7; 
        10'b1010111111: data <= 19'h00147; 
        10'b1011000000: data <= 19'h001d4; 
        10'b1011000001: data <= 19'h001ab; 
        10'b1011000010: data <= 19'h00007; 
        10'b1011000011: data <= 19'h7fef7; 
        10'b1011000100: data <= 19'h7ff97; 
        10'b1011000101: data <= 19'h7ff0c; 
        10'b1011000110: data <= 19'h7fc0a; 
        10'b1011000111: data <= 19'h7fb2e; 
        10'b1011001000: data <= 19'h7fc70; 
        10'b1011001001: data <= 19'h7fb00; 
        10'b1011001010: data <= 19'h7fcf2; 
        10'b1011001011: data <= 19'h7fc22; 
        10'b1011001100: data <= 19'h7fdc6; 
        10'b1011001101: data <= 19'h7ff99; 
        10'b1011001110: data <= 19'h000c5; 
        10'b1011001111: data <= 19'h00199; 
        10'b1011010000: data <= 19'h00027; 
        10'b1011010001: data <= 19'h00174; 
        10'b1011010010: data <= 19'h000dd; 
        10'b1011010011: data <= 19'h00213; 
        10'b1011010100: data <= 19'h00085; 
        10'b1011010101: data <= 19'h0009e; 
        10'b1011010110: data <= 19'h000e3; 
        10'b1011010111: data <= 19'h000c4; 
        10'b1011011000: data <= 19'h000df; 
        10'b1011011001: data <= 19'h001ae; 
        10'b1011011010: data <= 19'h0017e; 
        10'b1011011011: data <= 19'h00075; 
        10'b1011011100: data <= 19'h0019e; 
        10'b1011011101: data <= 19'h00226; 
        10'b1011011110: data <= 19'h00175; 
        10'b1011011111: data <= 19'h00158; 
        10'b1011100000: data <= 19'h001eb; 
        10'b1011100001: data <= 19'h001a0; 
        10'b1011100010: data <= 19'h0003a; 
        10'b1011100011: data <= 19'h00152; 
        10'b1011100100: data <= 19'h00134; 
        10'b1011100101: data <= 19'h000b2; 
        10'b1011100110: data <= 19'h7fff5; 
        10'b1011100111: data <= 19'h000a0; 
        10'b1011101000: data <= 19'h00168; 
        10'b1011101001: data <= 19'h0022e; 
        10'b1011101010: data <= 19'h0019b; 
        10'b1011101011: data <= 19'h00042; 
        10'b1011101100: data <= 19'h0017f; 
        10'b1011101101: data <= 19'h00167; 
        10'b1011101110: data <= 19'h00156; 
        10'b1011101111: data <= 19'h000a3; 
        10'b1011110000: data <= 19'h00090; 
        10'b1011110001: data <= 19'h0019f; 
        10'b1011110010: data <= 19'h00237; 
        10'b1011110011: data <= 19'h001cc; 
        10'b1011110100: data <= 19'h001cf; 
        10'b1011110101: data <= 19'h0024a; 
        10'b1011110110: data <= 19'h0005c; 
        10'b1011110111: data <= 19'h00144; 
        10'b1011111000: data <= 19'h00266; 
        10'b1011111001: data <= 19'h001e8; 
        10'b1011111010: data <= 19'h00229; 
        10'b1011111011: data <= 19'h001ff; 
        10'b1011111100: data <= 19'h0022a; 
        10'b1011111101: data <= 19'h00106; 
        10'b1011111110: data <= 19'h001e5; 
        10'b1011111111: data <= 19'h001f8; 
        10'b1100000000: data <= 19'h00032; 
        10'b1100000001: data <= 19'h00069; 
        10'b1100000010: data <= 19'h0025b; 
        10'b1100000011: data <= 19'h00189; 
        10'b1100000100: data <= 19'h0016a; 
        10'b1100000101: data <= 19'h00035; 
        10'b1100000110: data <= 19'h00107; 
        10'b1100000111: data <= 19'h00074; 
        10'b1100001000: data <= 19'h0006c; 
        10'b1100001001: data <= 19'h000c5; 
        10'b1100001010: data <= 19'h00163; 
        10'b1100001011: data <= 19'h00200; 
        10'b1100001100: data <= 19'h00238; 
        10'b1100001101: data <= 19'h0022a; 
        10'b1100001110: data <= 19'h00222; 
        10'b1100001111: data <= 19'h000b6; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 14) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 20'h003fe; 
        10'b0000000001: data <= 20'h001e7; 
        10'b0000000010: data <= 20'h00220; 
        10'b0000000011: data <= 20'h000e0; 
        10'b0000000100: data <= 20'h00362; 
        10'b0000000101: data <= 20'h0034b; 
        10'b0000000110: data <= 20'h003a2; 
        10'b0000000111: data <= 20'h000e7; 
        10'b0000001000: data <= 20'h0032b; 
        10'b0000001001: data <= 20'h000f8; 
        10'b0000001010: data <= 20'h00303; 
        10'b0000001011: data <= 20'h0026e; 
        10'b0000001100: data <= 20'h00364; 
        10'b0000001101: data <= 20'h00486; 
        10'b0000001110: data <= 20'h003fb; 
        10'b0000001111: data <= 20'h002ba; 
        10'b0000010000: data <= 20'h002c5; 
        10'b0000010001: data <= 20'h000fa; 
        10'b0000010010: data <= 20'h004a5; 
        10'b0000010011: data <= 20'h0049f; 
        10'b0000010100: data <= 20'h002a3; 
        10'b0000010101: data <= 20'h00362; 
        10'b0000010110: data <= 20'h0029d; 
        10'b0000010111: data <= 20'h0040e; 
        10'b0000011000: data <= 20'h0018b; 
        10'b0000011001: data <= 20'h00449; 
        10'b0000011010: data <= 20'h0029d; 
        10'b0000011011: data <= 20'h003c7; 
        10'b0000011100: data <= 20'h0007d; 
        10'b0000011101: data <= 20'h00403; 
        10'b0000011110: data <= 20'h0012f; 
        10'b0000011111: data <= 20'h002db; 
        10'b0000100000: data <= 20'h0028d; 
        10'b0000100001: data <= 20'h00102; 
        10'b0000100010: data <= 20'h0016c; 
        10'b0000100011: data <= 20'h003c4; 
        10'b0000100100: data <= 20'h0039e; 
        10'b0000100101: data <= 20'h002f0; 
        10'b0000100110: data <= 20'h002e9; 
        10'b0000100111: data <= 20'h00224; 
        10'b0000101000: data <= 20'h00377; 
        10'b0000101001: data <= 20'h003e7; 
        10'b0000101010: data <= 20'h0050c; 
        10'b0000101011: data <= 20'h00283; 
        10'b0000101100: data <= 20'h00208; 
        10'b0000101101: data <= 20'h0040e; 
        10'b0000101110: data <= 20'h002bb; 
        10'b0000101111: data <= 20'h001da; 
        10'b0000110000: data <= 20'h00465; 
        10'b0000110001: data <= 20'h0043b; 
        10'b0000110010: data <= 20'h001bc; 
        10'b0000110011: data <= 20'h00489; 
        10'b0000110100: data <= 20'h004dc; 
        10'b0000110101: data <= 20'h00293; 
        10'b0000110110: data <= 20'h00423; 
        10'b0000110111: data <= 20'h00354; 
        10'b0000111000: data <= 20'h00415; 
        10'b0000111001: data <= 20'h00312; 
        10'b0000111010: data <= 20'h004e4; 
        10'b0000111011: data <= 20'h000f3; 
        10'b0000111100: data <= 20'h000e9; 
        10'b0000111101: data <= 20'h00338; 
        10'b0000111110: data <= 20'h00261; 
        10'b0000111111: data <= 20'h0024a; 
        10'b0001000000: data <= 20'h0018a; 
        10'b0001000001: data <= 20'h002b2; 
        10'b0001000010: data <= 20'h00011; 
        10'b0001000011: data <= 20'h0015b; 
        10'b0001000100: data <= 20'h0002d; 
        10'b0001000101: data <= 20'h0012f; 
        10'b0001000110: data <= 20'h0027b; 
        10'b0001000111: data <= 20'h003fc; 
        10'b0001001000: data <= 20'h00304; 
        10'b0001001001: data <= 20'h00001; 
        10'b0001001010: data <= 20'h002fb; 
        10'b0001001011: data <= 20'h001c9; 
        10'b0001001100: data <= 20'h003eb; 
        10'b0001001101: data <= 20'h001b3; 
        10'b0001001110: data <= 20'h00450; 
        10'b0001001111: data <= 20'h00323; 
        10'b0001010000: data <= 20'h00361; 
        10'b0001010001: data <= 20'h00094; 
        10'b0001010010: data <= 20'h003ac; 
        10'b0001010011: data <= 20'h003c2; 
        10'b0001010100: data <= 20'h00174; 
        10'b0001010101: data <= 20'h001a1; 
        10'b0001010110: data <= 20'h002c0; 
        10'b0001010111: data <= 20'h00242; 
        10'b0001011000: data <= 20'h00498; 
        10'b0001011001: data <= 20'h0026c; 
        10'b0001011010: data <= 20'h00088; 
        10'b0001011011: data <= 20'h00480; 
        10'b0001011100: data <= 20'hfff81; 
        10'b0001011101: data <= 20'hfff18; 
        10'b0001011110: data <= 20'hfff20; 
        10'b0001011111: data <= 20'hffd80; 
        10'b0001100000: data <= 20'hfff1d; 
        10'b0001100001: data <= 20'h00055; 
        10'b0001100010: data <= 20'h001e0; 
        10'b0001100011: data <= 20'h003bf; 
        10'b0001100100: data <= 20'hffe24; 
        10'b0001100101: data <= 20'hfff52; 
        10'b0001100110: data <= 20'hfffe8; 
        10'b0001100111: data <= 20'hffd1d; 
        10'b0001101000: data <= 20'hfffb3; 
        10'b0001101001: data <= 20'h00130; 
        10'b0001101010: data <= 20'h002fe; 
        10'b0001101011: data <= 20'h002ed; 
        10'b0001101100: data <= 20'hfff77; 
        10'b0001101101: data <= 20'h00426; 
        10'b0001101110: data <= 20'h0018f; 
        10'b0001101111: data <= 20'h00462; 
        10'b0001110000: data <= 20'h00360; 
        10'b0001110001: data <= 20'h0020c; 
        10'b0001110010: data <= 20'h004a6; 
        10'b0001110011: data <= 20'h0049c; 
        10'b0001110100: data <= 20'h00084; 
        10'b0001110101: data <= 20'h000eb; 
        10'b0001110110: data <= 20'h0040f; 
        10'b0001110111: data <= 20'h00295; 
        10'b0001111000: data <= 20'h000fb; 
        10'b0001111001: data <= 20'hffbc2; 
        10'b0001111010: data <= 20'h00064; 
        10'b0001111011: data <= 20'h0017c; 
        10'b0001111100: data <= 20'h0024f; 
        10'b0001111101: data <= 20'h00421; 
        10'b0001111110: data <= 20'h004d7; 
        10'b0001111111: data <= 20'h009e7; 
        10'b0010000000: data <= 20'h002b5; 
        10'b0010000001: data <= 20'hffdeb; 
        10'b0010000010: data <= 20'hffdbc; 
        10'b0010000011: data <= 20'h0018a; 
        10'b0010000100: data <= 20'h0057a; 
        10'b0010000101: data <= 20'h00623; 
        10'b0010000110: data <= 20'h0061c; 
        10'b0010000111: data <= 20'h00727; 
        10'b0010001000: data <= 20'h003be; 
        10'b0010001001: data <= 20'h001c6; 
        10'b0010001010: data <= 20'h0018d; 
        10'b0010001011: data <= 20'h001b5; 
        10'b0010001100: data <= 20'h0009d; 
        10'b0010001101: data <= 20'h003ff; 
        10'b0010001110: data <= 20'h000c8; 
        10'b0010001111: data <= 20'h002d0; 
        10'b0010010000: data <= 20'h000b4; 
        10'b0010010001: data <= 20'h002b2; 
        10'b0010010010: data <= 20'h000cf; 
        10'b0010010011: data <= 20'hffef5; 
        10'b0010010100: data <= 20'hff717; 
        10'b0010010101: data <= 20'hff704; 
        10'b0010010110: data <= 20'hffbe2; 
        10'b0010010111: data <= 20'h0000e; 
        10'b0010011000: data <= 20'h00360; 
        10'b0010011001: data <= 20'h003cd; 
        10'b0010011010: data <= 20'h0069a; 
        10'b0010011011: data <= 20'h00521; 
        10'b0010011100: data <= 20'h00309; 
        10'b0010011101: data <= 20'hffb03; 
        10'b0010011110: data <= 20'hfff80; 
        10'b0010011111: data <= 20'h0010b; 
        10'b0010100000: data <= 20'h004e1; 
        10'b0010100001: data <= 20'h007da; 
        10'b0010100010: data <= 20'h00d11; 
        10'b0010100011: data <= 20'h00828; 
        10'b0010100100: data <= 20'h006ae; 
        10'b0010100101: data <= 20'hffe48; 
        10'b0010100110: data <= 20'h001d8; 
        10'b0010100111: data <= 20'h00105; 
        10'b0010101000: data <= 20'h000da; 
        10'b0010101001: data <= 20'h002e6; 
        10'b0010101010: data <= 20'h00088; 
        10'b0010101011: data <= 20'h00242; 
        10'b0010101100: data <= 20'h00087; 
        10'b0010101101: data <= 20'hffeab; 
        10'b0010101110: data <= 20'hffb19; 
        10'b0010101111: data <= 20'hffb28; 
        10'b0010110000: data <= 20'hff4dc; 
        10'b0010110001: data <= 20'hff289; 
        10'b0010110010: data <= 20'hff791; 
        10'b0010110011: data <= 20'hffe05; 
        10'b0010110100: data <= 20'hffdf0; 
        10'b0010110101: data <= 20'hffbc4; 
        10'b0010110110: data <= 20'hffe0d; 
        10'b0010110111: data <= 20'hff656; 
        10'b0010111000: data <= 20'hff59b; 
        10'b0010111001: data <= 20'hff587; 
        10'b0010111010: data <= 20'hffb9f; 
        10'b0010111011: data <= 20'hffcc3; 
        10'b0010111100: data <= 20'h004e6; 
        10'b0010111101: data <= 20'h00812; 
        10'b0010111110: data <= 20'h0077c; 
        10'b0010111111: data <= 20'h0064c; 
        10'b0011000000: data <= 20'h001a4; 
        10'b0011000001: data <= 20'hffea9; 
        10'b0011000010: data <= 20'h0001c; 
        10'b0011000011: data <= 20'h0025c; 
        10'b0011000100: data <= 20'h001e9; 
        10'b0011000101: data <= 20'h00114; 
        10'b0011000110: data <= 20'h00156; 
        10'b0011000111: data <= 20'h0004d; 
        10'b0011001000: data <= 20'h0032a; 
        10'b0011001001: data <= 20'hfff53; 
        10'b0011001010: data <= 20'hffb4c; 
        10'b0011001011: data <= 20'hff661; 
        10'b0011001100: data <= 20'hff0f7; 
        10'b0011001101: data <= 20'hfecdb; 
        10'b0011001110: data <= 20'hff300; 
        10'b0011001111: data <= 20'hffa52; 
        10'b0011010000: data <= 20'hffacc; 
        10'b0011010001: data <= 20'hff884; 
        10'b0011010010: data <= 20'hff6c0; 
        10'b0011010011: data <= 20'hff19f; 
        10'b0011010100: data <= 20'hff371; 
        10'b0011010101: data <= 20'hff437; 
        10'b0011010110: data <= 20'hff561; 
        10'b0011010111: data <= 20'hfffa3; 
        10'b0011011000: data <= 20'h0023a; 
        10'b0011011001: data <= 20'h00162; 
        10'b0011011010: data <= 20'h00152; 
        10'b0011011011: data <= 20'hffbf4; 
        10'b0011011100: data <= 20'hffa7b; 
        10'b0011011101: data <= 20'hffdcc; 
        10'b0011011110: data <= 20'h001cb; 
        10'b0011011111: data <= 20'h00218; 
        10'b0011100000: data <= 20'h00252; 
        10'b0011100001: data <= 20'h001f7; 
        10'b0011100010: data <= 20'h001ed; 
        10'b0011100011: data <= 20'h00418; 
        10'b0011100100: data <= 20'h0014f; 
        10'b0011100101: data <= 20'hfffde; 
        10'b0011100110: data <= 20'hffa69; 
        10'b0011100111: data <= 20'hff786; 
        10'b0011101000: data <= 20'hfee7a; 
        10'b0011101001: data <= 20'hfecfa; 
        10'b0011101010: data <= 20'hfede4; 
        10'b0011101011: data <= 20'hff641; 
        10'b0011101100: data <= 20'hffb87; 
        10'b0011101101: data <= 20'hffa7f; 
        10'b0011101110: data <= 20'hffb82; 
        10'b0011101111: data <= 20'h001f7; 
        10'b0011110000: data <= 20'hff808; 
        10'b0011110001: data <= 20'hffd4c; 
        10'b0011110010: data <= 20'hfff8d; 
        10'b0011110011: data <= 20'h00108; 
        10'b0011110100: data <= 20'hffa02; 
        10'b0011110101: data <= 20'hffa35; 
        10'b0011110110: data <= 20'hff6b9; 
        10'b0011110111: data <= 20'hff3d3; 
        10'b0011111000: data <= 20'hff650; 
        10'b0011111001: data <= 20'hffd9f; 
        10'b0011111010: data <= 20'h0039c; 
        10'b0011111011: data <= 20'h004c0; 
        10'b0011111100: data <= 20'h004cc; 
        10'b0011111101: data <= 20'h0011c; 
        10'b0011111110: data <= 20'h001f8; 
        10'b0011111111: data <= 20'h001ae; 
        10'b0100000000: data <= 20'hfffb2; 
        10'b0100000001: data <= 20'hfff78; 
        10'b0100000010: data <= 20'hff8e1; 
        10'b0100000011: data <= 20'hff942; 
        10'b0100000100: data <= 20'hff3f1; 
        10'b0100000101: data <= 20'hfed9e; 
        10'b0100000110: data <= 20'hfef28; 
        10'b0100000111: data <= 20'hff958; 
        10'b0100001000: data <= 20'hffb07; 
        10'b0100001001: data <= 20'h003c7; 
        10'b0100001010: data <= 20'h00be5; 
        10'b0100001011: data <= 20'h01109; 
        10'b0100001100: data <= 20'h00650; 
        10'b0100001101: data <= 20'hfff8f; 
        10'b0100001110: data <= 20'hffd27; 
        10'b0100001111: data <= 20'hff472; 
        10'b0100010000: data <= 20'hff1c9; 
        10'b0100010001: data <= 20'hff1fa; 
        10'b0100010010: data <= 20'hfee56; 
        10'b0100010011: data <= 20'hff0b1; 
        10'b0100010100: data <= 20'hff7ca; 
        10'b0100010101: data <= 20'h000f4; 
        10'b0100010110: data <= 20'h003f6; 
        10'b0100010111: data <= 20'h002df; 
        10'b0100011000: data <= 20'h0045f; 
        10'b0100011001: data <= 20'h004d8; 
        10'b0100011010: data <= 20'h00402; 
        10'b0100011011: data <= 20'h00086; 
        10'b0100011100: data <= 20'h00345; 
        10'b0100011101: data <= 20'hffc36; 
        10'b0100011110: data <= 20'hff944; 
        10'b0100011111: data <= 20'hffce1; 
        10'b0100100000: data <= 20'hff6a5; 
        10'b0100100001: data <= 20'hff683; 
        10'b0100100010: data <= 20'hff912; 
        10'b0100100011: data <= 20'hffb5e; 
        10'b0100100100: data <= 20'hffce1; 
        10'b0100100101: data <= 20'h00980; 
        10'b0100100110: data <= 20'h01ebf; 
        10'b0100100111: data <= 20'h02076; 
        10'b0100101000: data <= 20'h00f6a; 
        10'b0100101001: data <= 20'hfffab; 
        10'b0100101010: data <= 20'hff6c6; 
        10'b0100101011: data <= 20'hff4e0; 
        10'b0100101100: data <= 20'hff289; 
        10'b0100101101: data <= 20'hff3db; 
        10'b0100101110: data <= 20'hff48f; 
        10'b0100101111: data <= 20'hff8e5; 
        10'b0100110000: data <= 20'hffd9f; 
        10'b0100110001: data <= 20'hfff96; 
        10'b0100110010: data <= 20'h0041e; 
        10'b0100110011: data <= 20'h001b1; 
        10'b0100110100: data <= 20'h000d3; 
        10'b0100110101: data <= 20'h000be; 
        10'b0100110110: data <= 20'h00355; 
        10'b0100110111: data <= 20'h0038c; 
        10'b0100111000: data <= 20'h00003; 
        10'b0100111001: data <= 20'hffeee; 
        10'b0100111010: data <= 20'hfff71; 
        10'b0100111011: data <= 20'hffa27; 
        10'b0100111100: data <= 20'hffc38; 
        10'b0100111101: data <= 20'hffa2a; 
        10'b0100111110: data <= 20'hff76a; 
        10'b0100111111: data <= 20'hff308; 
        10'b0101000000: data <= 20'hffe84; 
        10'b0101000001: data <= 20'h0103f; 
        10'b0101000010: data <= 20'h02511; 
        10'b0101000011: data <= 20'h02746; 
        10'b0101000100: data <= 20'h00e8c; 
        10'b0101000101: data <= 20'hffcd2; 
        10'b0101000110: data <= 20'hffd13; 
        10'b0101000111: data <= 20'hff843; 
        10'b0101001000: data <= 20'hff7cf; 
        10'b0101001001: data <= 20'hff865; 
        10'b0101001010: data <= 20'hff8f6; 
        10'b0101001011: data <= 20'hffcb5; 
        10'b0101001100: data <= 20'hffe9b; 
        10'b0101001101: data <= 20'h00343; 
        10'b0101001110: data <= 20'h00493; 
        10'b0101001111: data <= 20'h00337; 
        10'b0101010000: data <= 20'h00081; 
        10'b0101010001: data <= 20'h00460; 
        10'b0101010010: data <= 20'h00219; 
        10'b0101010011: data <= 20'h0016c; 
        10'b0101010100: data <= 20'h00479; 
        10'b0101010101: data <= 20'hfff25; 
        10'b0101010110: data <= 20'hffea2; 
        10'b0101010111: data <= 20'hffe0f; 
        10'b0101011000: data <= 20'hffa6d; 
        10'b0101011001: data <= 20'hff8b2; 
        10'b0101011010: data <= 20'hff086; 
        10'b0101011011: data <= 20'hfea4a; 
        10'b0101011100: data <= 20'hfff4d; 
        10'b0101011101: data <= 20'h0107e; 
        10'b0101011110: data <= 20'h02ba2; 
        10'b0101011111: data <= 20'h01e43; 
        10'b0101100000: data <= 20'h005fe; 
        10'b0101100001: data <= 20'h0032c; 
        10'b0101100010: data <= 20'hffe23; 
        10'b0101100011: data <= 20'hff728; 
        10'b0101100100: data <= 20'hffa6b; 
        10'b0101100101: data <= 20'hffd4a; 
        10'b0101100110: data <= 20'hffe7a; 
        10'b0101100111: data <= 20'hffe1f; 
        10'b0101101000: data <= 20'h00049; 
        10'b0101101001: data <= 20'h00472; 
        10'b0101101010: data <= 20'h000ab; 
        10'b0101101011: data <= 20'h00320; 
        10'b0101101100: data <= 20'h00072; 
        10'b0101101101: data <= 20'h002f8; 
        10'b0101101110: data <= 20'h002c5; 
        10'b0101101111: data <= 20'h002f5; 
        10'b0101110000: data <= 20'h004ee; 
        10'b0101110001: data <= 20'h00008; 
        10'b0101110010: data <= 20'h0006a; 
        10'b0101110011: data <= 20'hffdcb; 
        10'b0101110100: data <= 20'hffd06; 
        10'b0101110101: data <= 20'hff3d3; 
        10'b0101110110: data <= 20'hfe62d; 
        10'b0101110111: data <= 20'hfe5cd; 
        10'b0101111000: data <= 20'h00009; 
        10'b0101111001: data <= 20'h00dc2; 
        10'b0101111010: data <= 20'h023f5; 
        10'b0101111011: data <= 20'h01452; 
        10'b0101111100: data <= 20'h0055f; 
        10'b0101111101: data <= 20'h0029c; 
        10'b0101111110: data <= 20'hff7cb; 
        10'b0101111111: data <= 20'hff414; 
        10'b0110000000: data <= 20'hffbac; 
        10'b0110000001: data <= 20'hffe7a; 
        10'b0110000010: data <= 20'hffe69; 
        10'b0110000011: data <= 20'hfff6d; 
        10'b0110000100: data <= 20'h00203; 
        10'b0110000101: data <= 20'h00301; 
        10'b0110000110: data <= 20'h00456; 
        10'b0110000111: data <= 20'h002ce; 
        10'b0110001000: data <= 20'h00230; 
        10'b0110001001: data <= 20'h004ae; 
        10'b0110001010: data <= 20'h002a2; 
        10'b0110001011: data <= 20'h003bf; 
        10'b0110001100: data <= 20'h003c3; 
        10'b0110001101: data <= 20'hffffc; 
        10'b0110001110: data <= 20'h000a5; 
        10'b0110001111: data <= 20'hffe90; 
        10'b0110010000: data <= 20'hff7f2; 
        10'b0110010001: data <= 20'hff22c; 
        10'b0110010010: data <= 20'hfe645; 
        10'b0110010011: data <= 20'hfec79; 
        10'b0110010100: data <= 20'hfff91; 
        10'b0110010101: data <= 20'h00df7; 
        10'b0110010110: data <= 20'h01eab; 
        10'b0110010111: data <= 20'h013c0; 
        10'b0110011000: data <= 20'h005e7; 
        10'b0110011001: data <= 20'hff50b; 
        10'b0110011010: data <= 20'hff128; 
        10'b0110011011: data <= 20'hff4ba; 
        10'b0110011100: data <= 20'hff955; 
        10'b0110011101: data <= 20'hffe12; 
        10'b0110011110: data <= 20'hffde7; 
        10'b0110011111: data <= 20'hffe91; 
        10'b0110100000: data <= 20'h00357; 
        10'b0110100001: data <= 20'h00083; 
        10'b0110100010: data <= 20'h000ed; 
        10'b0110100011: data <= 20'h002aa; 
        10'b0110100100: data <= 20'h004f6; 
        10'b0110100101: data <= 20'h000d0; 
        10'b0110100110: data <= 20'h0032f; 
        10'b0110100111: data <= 20'h00204; 
        10'b0110101000: data <= 20'h00123; 
        10'b0110101001: data <= 20'h002e3; 
        10'b0110101010: data <= 20'hffd30; 
        10'b0110101011: data <= 20'hffccc; 
        10'b0110101100: data <= 20'hffaec; 
        10'b0110101101: data <= 20'hff0e0; 
        10'b0110101110: data <= 20'hfef0b; 
        10'b0110101111: data <= 20'hffbba; 
        10'b0110110000: data <= 20'h00639; 
        10'b0110110001: data <= 20'h013a2; 
        10'b0110110010: data <= 20'h020d1; 
        10'b0110110011: data <= 20'h00b9b; 
        10'b0110110100: data <= 20'h00220; 
        10'b0110110101: data <= 20'hfeb58; 
        10'b0110110110: data <= 20'hfedb2; 
        10'b0110110111: data <= 20'hff4cc; 
        10'b0110111000: data <= 20'hff942; 
        10'b0110111001: data <= 20'hffb28; 
        10'b0110111010: data <= 20'hffec7; 
        10'b0110111011: data <= 20'h0005e; 
        10'b0110111100: data <= 20'h001c0; 
        10'b0110111101: data <= 20'h0023d; 
        10'b0110111110: data <= 20'h0049e; 
        10'b0110111111: data <= 20'h000c5; 
        10'b0111000000: data <= 20'h004ce; 
        10'b0111000001: data <= 20'h00259; 
        10'b0111000010: data <= 20'h00464; 
        10'b0111000011: data <= 20'h002ad; 
        10'b0111000100: data <= 20'h0016b; 
        10'b0111000101: data <= 20'hffe0d; 
        10'b0111000110: data <= 20'hffb8b; 
        10'b0111000111: data <= 20'hffb35; 
        10'b0111001000: data <= 20'hff449; 
        10'b0111001001: data <= 20'hff8fc; 
        10'b0111001010: data <= 20'hffa6a; 
        10'b0111001011: data <= 20'hffce6; 
        10'b0111001100: data <= 20'hfff37; 
        10'b0111001101: data <= 20'h019d2; 
        10'b0111001110: data <= 20'h01efb; 
        10'b0111001111: data <= 20'h001c7; 
        10'b0111010000: data <= 20'hff669; 
        10'b0111010001: data <= 20'hfe9a7; 
        10'b0111010010: data <= 20'hfed83; 
        10'b0111010011: data <= 20'hff419; 
        10'b0111010100: data <= 20'hff6f5; 
        10'b0111010101: data <= 20'hffc25; 
        10'b0111010110: data <= 20'hffc16; 
        10'b0111010111: data <= 20'h0000c; 
        10'b0111011000: data <= 20'hffe46; 
        10'b0111011001: data <= 20'h00045; 
        10'b0111011010: data <= 20'h0012d; 
        10'b0111011011: data <= 20'h0027e; 
        10'b0111011100: data <= 20'h001fe; 
        10'b0111011101: data <= 20'h004be; 
        10'b0111011110: data <= 20'h0010e; 
        10'b0111011111: data <= 20'h004ae; 
        10'b0111100000: data <= 20'h00375; 
        10'b0111100001: data <= 20'hffd48; 
        10'b0111100010: data <= 20'hff630; 
        10'b0111100011: data <= 20'hff560; 
        10'b0111100100: data <= 20'hff865; 
        10'b0111100101: data <= 20'hffb22; 
        10'b0111100110: data <= 20'h0037e; 
        10'b0111100111: data <= 20'h0000a; 
        10'b0111101000: data <= 20'h00870; 
        10'b0111101001: data <= 20'h01d93; 
        10'b0111101010: data <= 20'h0195d; 
        10'b0111101011: data <= 20'hffada; 
        10'b0111101100: data <= 20'hfee60; 
        10'b0111101101: data <= 20'hfe992; 
        10'b0111101110: data <= 20'hfeda0; 
        10'b0111101111: data <= 20'hff463; 
        10'b0111110000: data <= 20'hffba2; 
        10'b0111110001: data <= 20'hffdce; 
        10'b0111110010: data <= 20'hffe6d; 
        10'b0111110011: data <= 20'hffde4; 
        10'b0111110100: data <= 20'hffc62; 
        10'b0111110101: data <= 20'h0010a; 
        10'b0111110110: data <= 20'h002c4; 
        10'b0111110111: data <= 20'h0033c; 
        10'b0111111000: data <= 20'h002ef; 
        10'b0111111001: data <= 20'h002b4; 
        10'b0111111010: data <= 20'h001a9; 
        10'b0111111011: data <= 20'h003e8; 
        10'b0111111100: data <= 20'h0022b; 
        10'b0111111101: data <= 20'hffc20; 
        10'b0111111110: data <= 20'hff589; 
        10'b0111111111: data <= 20'hff59e; 
        10'b1000000000: data <= 20'hffc1b; 
        10'b1000000001: data <= 20'h003fb; 
        10'b1000000010: data <= 20'h00349; 
        10'b1000000011: data <= 20'h00543; 
        10'b1000000100: data <= 20'h00db9; 
        10'b1000000101: data <= 20'h01617; 
        10'b1000000110: data <= 20'h00f46; 
        10'b1000000111: data <= 20'hff5f5; 
        10'b1000001000: data <= 20'hfef80; 
        10'b1000001001: data <= 20'hff1dd; 
        10'b1000001010: data <= 20'hff3ee; 
        10'b1000001011: data <= 20'hff7e9; 
        10'b1000001100: data <= 20'hffc06; 
        10'b1000001101: data <= 20'hff947; 
        10'b1000001110: data <= 20'hffd04; 
        10'b1000001111: data <= 20'hffb6b; 
        10'b1000010000: data <= 20'hffd33; 
        10'b1000010001: data <= 20'h00289; 
        10'b1000010010: data <= 20'h00466; 
        10'b1000010011: data <= 20'h0047e; 
        10'b1000010100: data <= 20'h0049e; 
        10'b1000010101: data <= 20'h00341; 
        10'b1000010110: data <= 20'h00363; 
        10'b1000010111: data <= 20'h003c0; 
        10'b1000011000: data <= 20'h00070; 
        10'b1000011001: data <= 20'hffa30; 
        10'b1000011010: data <= 20'hff304; 
        10'b1000011011: data <= 20'hff73d; 
        10'b1000011100: data <= 20'hffc6c; 
        10'b1000011101: data <= 20'h00210; 
        10'b1000011110: data <= 20'h00109; 
        10'b1000011111: data <= 20'h000b8; 
        10'b1000100000: data <= 20'h001d2; 
        10'b1000100001: data <= 20'h00a2c; 
        10'b1000100010: data <= 20'h0023e; 
        10'b1000100011: data <= 20'hff7b2; 
        10'b1000100100: data <= 20'hff916; 
        10'b1000100101: data <= 20'hff9fb; 
        10'b1000100110: data <= 20'hff870; 
        10'b1000100111: data <= 20'hffa23; 
        10'b1000101000: data <= 20'hff76b; 
        10'b1000101001: data <= 20'hff8d9; 
        10'b1000101010: data <= 20'hffbaf; 
        10'b1000101011: data <= 20'hffc33; 
        10'b1000101100: data <= 20'h00035; 
        10'b1000101101: data <= 20'h00175; 
        10'b1000101110: data <= 20'h0019a; 
        10'b1000101111: data <= 20'h000a3; 
        10'b1000110000: data <= 20'h000bc; 
        10'b1000110001: data <= 20'h004db; 
        10'b1000110010: data <= 20'h0029e; 
        10'b1000110011: data <= 20'h001ad; 
        10'b1000110100: data <= 20'hffeb3; 
        10'b1000110101: data <= 20'hffbdd; 
        10'b1000110110: data <= 20'hfff39; 
        10'b1000110111: data <= 20'hffd27; 
        10'b1000111000: data <= 20'hfffee; 
        10'b1000111001: data <= 20'h00137; 
        10'b1000111010: data <= 20'hffccf; 
        10'b1000111011: data <= 20'hffeda; 
        10'b1000111100: data <= 20'hffaca; 
        10'b1000111101: data <= 20'hffe38; 
        10'b1000111110: data <= 20'hffeb4; 
        10'b1000111111: data <= 20'h00055; 
        10'b1001000000: data <= 20'h004f2; 
        10'b1001000001: data <= 20'h001c7; 
        10'b1001000010: data <= 20'hffe22; 
        10'b1001000011: data <= 20'hff90d; 
        10'b1001000100: data <= 20'hff777; 
        10'b1001000101: data <= 20'hff819; 
        10'b1001000110: data <= 20'hff9cb; 
        10'b1001000111: data <= 20'hffe9a; 
        10'b1001001000: data <= 20'h000a8; 
        10'b1001001001: data <= 20'h003f7; 
        10'b1001001010: data <= 20'h00195; 
        10'b1001001011: data <= 20'h004e1; 
        10'b1001001100: data <= 20'h00378; 
        10'b1001001101: data <= 20'h001d3; 
        10'b1001001110: data <= 20'h002d6; 
        10'b1001001111: data <= 20'h00365; 
        10'b1001010000: data <= 20'h002b2; 
        10'b1001010001: data <= 20'h00747; 
        10'b1001010010: data <= 20'h005fc; 
        10'b1001010011: data <= 20'h002d1; 
        10'b1001010100: data <= 20'h00078; 
        10'b1001010101: data <= 20'hffdee; 
        10'b1001010110: data <= 20'h00016; 
        10'b1001010111: data <= 20'hffbcd; 
        10'b1001011000: data <= 20'hff676; 
        10'b1001011001: data <= 20'hff51d; 
        10'b1001011010: data <= 20'hfff05; 
        10'b1001011011: data <= 20'h00345; 
        10'b1001011100: data <= 20'h00539; 
        10'b1001011101: data <= 20'h005f3; 
        10'b1001011110: data <= 20'h0041a; 
        10'b1001011111: data <= 20'hff917; 
        10'b1001100000: data <= 20'hff934; 
        10'b1001100001: data <= 20'hff83e; 
        10'b1001100010: data <= 20'hffaaa; 
        10'b1001100011: data <= 20'hffcec; 
        10'b1001100100: data <= 20'h000b1; 
        10'b1001100101: data <= 20'h0021c; 
        10'b1001100110: data <= 20'h0006a; 
        10'b1001100111: data <= 20'h00099; 
        10'b1001101000: data <= 20'h002b2; 
        10'b1001101001: data <= 20'h002c0; 
        10'b1001101010: data <= 20'h00319; 
        10'b1001101011: data <= 20'h000a2; 
        10'b1001101100: data <= 20'h0064e; 
        10'b1001101101: data <= 20'h00e14; 
        10'b1001101110: data <= 20'h00e94; 
        10'b1001101111: data <= 20'h008cd; 
        10'b1001110000: data <= 20'h00132; 
        10'b1001110001: data <= 20'hfff06; 
        10'b1001110010: data <= 20'hffca9; 
        10'b1001110011: data <= 20'hff21b; 
        10'b1001110100: data <= 20'hfe971; 
        10'b1001110101: data <= 20'hfeec1; 
        10'b1001110110: data <= 20'h0000d; 
        10'b1001110111: data <= 20'h00361; 
        10'b1001111000: data <= 20'h00ced; 
        10'b1001111001: data <= 20'h01532; 
        10'b1001111010: data <= 20'h00946; 
        10'b1001111011: data <= 20'h001ef; 
        10'b1001111100: data <= 20'hffb3a; 
        10'b1001111101: data <= 20'hffc48; 
        10'b1001111110: data <= 20'hfffab; 
        10'b1001111111: data <= 20'h000a1; 
        10'b1010000000: data <= 20'h0004c; 
        10'b1010000001: data <= 20'h0020e; 
        10'b1010000010: data <= 20'h004b1; 
        10'b1010000011: data <= 20'h00242; 
        10'b1010000100: data <= 20'h0045d; 
        10'b1010000101: data <= 20'h002bb; 
        10'b1010000110: data <= 20'h0037e; 
        10'b1010000111: data <= 20'h001f1; 
        10'b1010001000: data <= 20'h005a1; 
        10'b1010001001: data <= 20'h00c1b; 
        10'b1010001010: data <= 20'h00ce6; 
        10'b1010001011: data <= 20'h005eb; 
        10'b1010001100: data <= 20'h001a1; 
        10'b1010001101: data <= 20'hffcff; 
        10'b1010001110: data <= 20'hffdf4; 
        10'b1010001111: data <= 20'hff824; 
        10'b1010010000: data <= 20'hffa84; 
        10'b1010010001: data <= 20'hffb1a; 
        10'b1010010010: data <= 20'hff973; 
        10'b1010010011: data <= 20'h00290; 
        10'b1010010100: data <= 20'h00f09; 
        10'b1010010101: data <= 20'h01223; 
        10'b1010010110: data <= 20'h00826; 
        10'b1010010111: data <= 20'hffe8d; 
        10'b1010011000: data <= 20'hffc89; 
        10'b1010011001: data <= 20'hffaa4; 
        10'b1010011010: data <= 20'hffe27; 
        10'b1010011011: data <= 20'hffe4c; 
        10'b1010011100: data <= 20'h00111; 
        10'b1010011101: data <= 20'h0008a; 
        10'b1010011110: data <= 20'h00101; 
        10'b1010011111: data <= 20'h0007f; 
        10'b1010100000: data <= 20'h00110; 
        10'b1010100001: data <= 20'h000ac; 
        10'b1010100010: data <= 20'h001c5; 
        10'b1010100011: data <= 20'h0008e; 
        10'b1010100100: data <= 20'h002bf; 
        10'b1010100101: data <= 20'h0055a; 
        10'b1010100110: data <= 20'h00587; 
        10'b1010100111: data <= 20'hffe38; 
        10'b1010101000: data <= 20'hff7fb; 
        10'b1010101001: data <= 20'hff7f1; 
        10'b1010101010: data <= 20'hff1d5; 
        10'b1010101011: data <= 20'hff26f; 
        10'b1010101100: data <= 20'hff3d4; 
        10'b1010101101: data <= 20'hff593; 
        10'b1010101110: data <= 20'hff59f; 
        10'b1010101111: data <= 20'hff599; 
        10'b1010110000: data <= 20'hffcfe; 
        10'b1010110001: data <= 20'h00142; 
        10'b1010110010: data <= 20'h0024c; 
        10'b1010110011: data <= 20'h00354; 
        10'b1010110100: data <= 20'h002ca; 
        10'b1010110101: data <= 20'h000ac; 
        10'b1010110110: data <= 20'h00172; 
        10'b1010110111: data <= 20'h003dd; 
        10'b1010111000: data <= 20'h0012c; 
        10'b1010111001: data <= 20'h001e7; 
        10'b1010111010: data <= 20'h003aa; 
        10'b1010111011: data <= 20'h00136; 
        10'b1010111100: data <= 20'h004bd; 
        10'b1010111101: data <= 20'h00182; 
        10'b1010111110: data <= 20'h001cf; 
        10'b1010111111: data <= 20'h0028f; 
        10'b1011000000: data <= 20'h003a8; 
        10'b1011000001: data <= 20'h00356; 
        10'b1011000010: data <= 20'h0000d; 
        10'b1011000011: data <= 20'hffdee; 
        10'b1011000100: data <= 20'hfff2e; 
        10'b1011000101: data <= 20'hffe18; 
        10'b1011000110: data <= 20'hff814; 
        10'b1011000111: data <= 20'hff65b; 
        10'b1011001000: data <= 20'hff8df; 
        10'b1011001001: data <= 20'hff601; 
        10'b1011001010: data <= 20'hff9e4; 
        10'b1011001011: data <= 20'hff843; 
        10'b1011001100: data <= 20'hffb8c; 
        10'b1011001101: data <= 20'hfff32; 
        10'b1011001110: data <= 20'h0018a; 
        10'b1011001111: data <= 20'h00332; 
        10'b1011010000: data <= 20'h0004e; 
        10'b1011010001: data <= 20'h002e8; 
        10'b1011010010: data <= 20'h001ba; 
        10'b1011010011: data <= 20'h00425; 
        10'b1011010100: data <= 20'h0010b; 
        10'b1011010101: data <= 20'h0013c; 
        10'b1011010110: data <= 20'h001c6; 
        10'b1011010111: data <= 20'h00187; 
        10'b1011011000: data <= 20'h001be; 
        10'b1011011001: data <= 20'h0035b; 
        10'b1011011010: data <= 20'h002fc; 
        10'b1011011011: data <= 20'h000ea; 
        10'b1011011100: data <= 20'h0033b; 
        10'b1011011101: data <= 20'h0044c; 
        10'b1011011110: data <= 20'h002ea; 
        10'b1011011111: data <= 20'h002b0; 
        10'b1011100000: data <= 20'h003d6; 
        10'b1011100001: data <= 20'h00340; 
        10'b1011100010: data <= 20'h00074; 
        10'b1011100011: data <= 20'h002a5; 
        10'b1011100100: data <= 20'h00268; 
        10'b1011100101: data <= 20'h00164; 
        10'b1011100110: data <= 20'hfffeb; 
        10'b1011100111: data <= 20'h00140; 
        10'b1011101000: data <= 20'h002d1; 
        10'b1011101001: data <= 20'h0045c; 
        10'b1011101010: data <= 20'h00337; 
        10'b1011101011: data <= 20'h00083; 
        10'b1011101100: data <= 20'h002fd; 
        10'b1011101101: data <= 20'h002ce; 
        10'b1011101110: data <= 20'h002ad; 
        10'b1011101111: data <= 20'h00146; 
        10'b1011110000: data <= 20'h00120; 
        10'b1011110001: data <= 20'h0033e; 
        10'b1011110010: data <= 20'h0046e; 
        10'b1011110011: data <= 20'h00399; 
        10'b1011110100: data <= 20'h0039e; 
        10'b1011110101: data <= 20'h00493; 
        10'b1011110110: data <= 20'h000b9; 
        10'b1011110111: data <= 20'h00288; 
        10'b1011111000: data <= 20'h004cd; 
        10'b1011111001: data <= 20'h003d1; 
        10'b1011111010: data <= 20'h00453; 
        10'b1011111011: data <= 20'h003fe; 
        10'b1011111100: data <= 20'h00454; 
        10'b1011111101: data <= 20'h0020b; 
        10'b1011111110: data <= 20'h003ca; 
        10'b1011111111: data <= 20'h003f0; 
        10'b1100000000: data <= 20'h00065; 
        10'b1100000001: data <= 20'h000d3; 
        10'b1100000010: data <= 20'h004b6; 
        10'b1100000011: data <= 20'h00312; 
        10'b1100000100: data <= 20'h002d4; 
        10'b1100000101: data <= 20'h00069; 
        10'b1100000110: data <= 20'h0020e; 
        10'b1100000111: data <= 20'h000e7; 
        10'b1100001000: data <= 20'h000d7; 
        10'b1100001001: data <= 20'h0018a; 
        10'b1100001010: data <= 20'h002c7; 
        10'b1100001011: data <= 20'h003ff; 
        10'b1100001100: data <= 20'h0046f; 
        10'b1100001101: data <= 20'h00454; 
        10'b1100001110: data <= 20'h00443; 
        10'b1100001111: data <= 20'h0016c; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 15) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 21'h0007fb; 
        10'b0000000001: data <= 21'h0003ce; 
        10'b0000000010: data <= 21'h000440; 
        10'b0000000011: data <= 21'h0001bf; 
        10'b0000000100: data <= 21'h0006c4; 
        10'b0000000101: data <= 21'h000696; 
        10'b0000000110: data <= 21'h000745; 
        10'b0000000111: data <= 21'h0001ce; 
        10'b0000001000: data <= 21'h000656; 
        10'b0000001001: data <= 21'h0001f1; 
        10'b0000001010: data <= 21'h000606; 
        10'b0000001011: data <= 21'h0004dc; 
        10'b0000001100: data <= 21'h0006c8; 
        10'b0000001101: data <= 21'h00090d; 
        10'b0000001110: data <= 21'h0007f5; 
        10'b0000001111: data <= 21'h000575; 
        10'b0000010000: data <= 21'h00058a; 
        10'b0000010001: data <= 21'h0001f3; 
        10'b0000010010: data <= 21'h00094a; 
        10'b0000010011: data <= 21'h00093d; 
        10'b0000010100: data <= 21'h000546; 
        10'b0000010101: data <= 21'h0006c4; 
        10'b0000010110: data <= 21'h00053a; 
        10'b0000010111: data <= 21'h00081b; 
        10'b0000011000: data <= 21'h000315; 
        10'b0000011001: data <= 21'h000891; 
        10'b0000011010: data <= 21'h00053a; 
        10'b0000011011: data <= 21'h00078e; 
        10'b0000011100: data <= 21'h0000fa; 
        10'b0000011101: data <= 21'h000806; 
        10'b0000011110: data <= 21'h00025e; 
        10'b0000011111: data <= 21'h0005b6; 
        10'b0000100000: data <= 21'h000519; 
        10'b0000100001: data <= 21'h000205; 
        10'b0000100010: data <= 21'h0002d8; 
        10'b0000100011: data <= 21'h000789; 
        10'b0000100100: data <= 21'h00073c; 
        10'b0000100101: data <= 21'h0005e1; 
        10'b0000100110: data <= 21'h0005d2; 
        10'b0000100111: data <= 21'h000449; 
        10'b0000101000: data <= 21'h0006ed; 
        10'b0000101001: data <= 21'h0007cf; 
        10'b0000101010: data <= 21'h000a19; 
        10'b0000101011: data <= 21'h000506; 
        10'b0000101100: data <= 21'h000410; 
        10'b0000101101: data <= 21'h00081d; 
        10'b0000101110: data <= 21'h000576; 
        10'b0000101111: data <= 21'h0003b4; 
        10'b0000110000: data <= 21'h0008ca; 
        10'b0000110001: data <= 21'h000875; 
        10'b0000110010: data <= 21'h000377; 
        10'b0000110011: data <= 21'h000912; 
        10'b0000110100: data <= 21'h0009b7; 
        10'b0000110101: data <= 21'h000525; 
        10'b0000110110: data <= 21'h000847; 
        10'b0000110111: data <= 21'h0006a7; 
        10'b0000111000: data <= 21'h00082b; 
        10'b0000111001: data <= 21'h000623; 
        10'b0000111010: data <= 21'h0009c9; 
        10'b0000111011: data <= 21'h0001e5; 
        10'b0000111100: data <= 21'h0001d3; 
        10'b0000111101: data <= 21'h000670; 
        10'b0000111110: data <= 21'h0004c2; 
        10'b0000111111: data <= 21'h000495; 
        10'b0001000000: data <= 21'h000314; 
        10'b0001000001: data <= 21'h000564; 
        10'b0001000010: data <= 21'h000023; 
        10'b0001000011: data <= 21'h0002b5; 
        10'b0001000100: data <= 21'h000059; 
        10'b0001000101: data <= 21'h00025e; 
        10'b0001000110: data <= 21'h0004f6; 
        10'b0001000111: data <= 21'h0007f8; 
        10'b0001001000: data <= 21'h000609; 
        10'b0001001001: data <= 21'h000001; 
        10'b0001001010: data <= 21'h0005f5; 
        10'b0001001011: data <= 21'h000393; 
        10'b0001001100: data <= 21'h0007d6; 
        10'b0001001101: data <= 21'h000367; 
        10'b0001001110: data <= 21'h0008a0; 
        10'b0001001111: data <= 21'h000646; 
        10'b0001010000: data <= 21'h0006c1; 
        10'b0001010001: data <= 21'h000127; 
        10'b0001010010: data <= 21'h000757; 
        10'b0001010011: data <= 21'h000784; 
        10'b0001010100: data <= 21'h0002e8; 
        10'b0001010101: data <= 21'h000343; 
        10'b0001010110: data <= 21'h000580; 
        10'b0001010111: data <= 21'h000484; 
        10'b0001011000: data <= 21'h000930; 
        10'b0001011001: data <= 21'h0004d7; 
        10'b0001011010: data <= 21'h00010f; 
        10'b0001011011: data <= 21'h0008ff; 
        10'b0001011100: data <= 21'h1fff02; 
        10'b0001011101: data <= 21'h1ffe2f; 
        10'b0001011110: data <= 21'h1ffe41; 
        10'b0001011111: data <= 21'h1ffaff; 
        10'b0001100000: data <= 21'h1ffe3b; 
        10'b0001100001: data <= 21'h0000ab; 
        10'b0001100010: data <= 21'h0003bf; 
        10'b0001100011: data <= 21'h00077e; 
        10'b0001100100: data <= 21'h1ffc49; 
        10'b0001100101: data <= 21'h1ffea5; 
        10'b0001100110: data <= 21'h1fffcf; 
        10'b0001100111: data <= 21'h1ffa3a; 
        10'b0001101000: data <= 21'h1fff67; 
        10'b0001101001: data <= 21'h000260; 
        10'b0001101010: data <= 21'h0005fc; 
        10'b0001101011: data <= 21'h0005da; 
        10'b0001101100: data <= 21'h1ffeed; 
        10'b0001101101: data <= 21'h00084d; 
        10'b0001101110: data <= 21'h00031f; 
        10'b0001101111: data <= 21'h0008c4; 
        10'b0001110000: data <= 21'h0006c0; 
        10'b0001110001: data <= 21'h000418; 
        10'b0001110010: data <= 21'h00094c; 
        10'b0001110011: data <= 21'h000937; 
        10'b0001110100: data <= 21'h000107; 
        10'b0001110101: data <= 21'h0001d5; 
        10'b0001110110: data <= 21'h00081e; 
        10'b0001110111: data <= 21'h00052a; 
        10'b0001111000: data <= 21'h0001f5; 
        10'b0001111001: data <= 21'h1ff784; 
        10'b0001111010: data <= 21'h0000c8; 
        10'b0001111011: data <= 21'h0002f8; 
        10'b0001111100: data <= 21'h00049e; 
        10'b0001111101: data <= 21'h000842; 
        10'b0001111110: data <= 21'h0009af; 
        10'b0001111111: data <= 21'h0013cd; 
        10'b0010000000: data <= 21'h000569; 
        10'b0010000001: data <= 21'h1ffbd7; 
        10'b0010000010: data <= 21'h1ffb77; 
        10'b0010000011: data <= 21'h000313; 
        10'b0010000100: data <= 21'h000af4; 
        10'b0010000101: data <= 21'h000c46; 
        10'b0010000110: data <= 21'h000c37; 
        10'b0010000111: data <= 21'h000e4f; 
        10'b0010001000: data <= 21'h00077b; 
        10'b0010001001: data <= 21'h00038b; 
        10'b0010001010: data <= 21'h00031a; 
        10'b0010001011: data <= 21'h00036a; 
        10'b0010001100: data <= 21'h000139; 
        10'b0010001101: data <= 21'h0007fd; 
        10'b0010001110: data <= 21'h000190; 
        10'b0010001111: data <= 21'h00059f; 
        10'b0010010000: data <= 21'h000168; 
        10'b0010010001: data <= 21'h000563; 
        10'b0010010010: data <= 21'h00019e; 
        10'b0010010011: data <= 21'h1ffde9; 
        10'b0010010100: data <= 21'h1fee2e; 
        10'b0010010101: data <= 21'h1fee07; 
        10'b0010010110: data <= 21'h1ff7c4; 
        10'b0010010111: data <= 21'h00001c; 
        10'b0010011000: data <= 21'h0006c0; 
        10'b0010011001: data <= 21'h000799; 
        10'b0010011010: data <= 21'h000d34; 
        10'b0010011011: data <= 21'h000a42; 
        10'b0010011100: data <= 21'h000611; 
        10'b0010011101: data <= 21'h1ff605; 
        10'b0010011110: data <= 21'h1ffeff; 
        10'b0010011111: data <= 21'h000217; 
        10'b0010100000: data <= 21'h0009c1; 
        10'b0010100001: data <= 21'h000fb5; 
        10'b0010100010: data <= 21'h001a23; 
        10'b0010100011: data <= 21'h00104f; 
        10'b0010100100: data <= 21'h000d5b; 
        10'b0010100101: data <= 21'h1ffc90; 
        10'b0010100110: data <= 21'h0003b1; 
        10'b0010100111: data <= 21'h00020a; 
        10'b0010101000: data <= 21'h0001b4; 
        10'b0010101001: data <= 21'h0005cc; 
        10'b0010101010: data <= 21'h000110; 
        10'b0010101011: data <= 21'h000484; 
        10'b0010101100: data <= 21'h00010e; 
        10'b0010101101: data <= 21'h1ffd57; 
        10'b0010101110: data <= 21'h1ff631; 
        10'b0010101111: data <= 21'h1ff64f; 
        10'b0010110000: data <= 21'h1fe9b8; 
        10'b0010110001: data <= 21'h1fe513; 
        10'b0010110010: data <= 21'h1fef22; 
        10'b0010110011: data <= 21'h1ffc0b; 
        10'b0010110100: data <= 21'h1ffbe1; 
        10'b0010110101: data <= 21'h1ff788; 
        10'b0010110110: data <= 21'h1ffc1a; 
        10'b0010110111: data <= 21'h1fecab; 
        10'b0010111000: data <= 21'h1feb36; 
        10'b0010111001: data <= 21'h1feb0d; 
        10'b0010111010: data <= 21'h1ff73d; 
        10'b0010111011: data <= 21'h1ff986; 
        10'b0010111100: data <= 21'h0009cd; 
        10'b0010111101: data <= 21'h001024; 
        10'b0010111110: data <= 21'h000ef7; 
        10'b0010111111: data <= 21'h000c98; 
        10'b0011000000: data <= 21'h000348; 
        10'b0011000001: data <= 21'h1ffd53; 
        10'b0011000010: data <= 21'h000038; 
        10'b0011000011: data <= 21'h0004b9; 
        10'b0011000100: data <= 21'h0003d2; 
        10'b0011000101: data <= 21'h000227; 
        10'b0011000110: data <= 21'h0002ac; 
        10'b0011000111: data <= 21'h000099; 
        10'b0011001000: data <= 21'h000653; 
        10'b0011001001: data <= 21'h1ffea6; 
        10'b0011001010: data <= 21'h1ff699; 
        10'b0011001011: data <= 21'h1fecc3; 
        10'b0011001100: data <= 21'h1fe1ee; 
        10'b0011001101: data <= 21'h1fd9b6; 
        10'b0011001110: data <= 21'h1fe601; 
        10'b0011001111: data <= 21'h1ff4a3; 
        10'b0011010000: data <= 21'h1ff599; 
        10'b0011010001: data <= 21'h1ff109; 
        10'b0011010010: data <= 21'h1fed81; 
        10'b0011010011: data <= 21'h1fe33d; 
        10'b0011010100: data <= 21'h1fe6e2; 
        10'b0011010101: data <= 21'h1fe86d; 
        10'b0011010110: data <= 21'h1feac1; 
        10'b0011010111: data <= 21'h1fff47; 
        10'b0011011000: data <= 21'h000475; 
        10'b0011011001: data <= 21'h0002c4; 
        10'b0011011010: data <= 21'h0002a3; 
        10'b0011011011: data <= 21'h1ff7e9; 
        10'b0011011100: data <= 21'h1ff4f7; 
        10'b0011011101: data <= 21'h1ffb97; 
        10'b0011011110: data <= 21'h000396; 
        10'b0011011111: data <= 21'h000430; 
        10'b0011100000: data <= 21'h0004a4; 
        10'b0011100001: data <= 21'h0003ed; 
        10'b0011100010: data <= 21'h0003da; 
        10'b0011100011: data <= 21'h000830; 
        10'b0011100100: data <= 21'h00029e; 
        10'b0011100101: data <= 21'h1fffbc; 
        10'b0011100110: data <= 21'h1ff4d1; 
        10'b0011100111: data <= 21'h1fef0c; 
        10'b0011101000: data <= 21'h1fdcf4; 
        10'b0011101001: data <= 21'h1fd9f3; 
        10'b0011101010: data <= 21'h1fdbc7; 
        10'b0011101011: data <= 21'h1fec82; 
        10'b0011101100: data <= 21'h1ff70d; 
        10'b0011101101: data <= 21'h1ff4fe; 
        10'b0011101110: data <= 21'h1ff704; 
        10'b0011101111: data <= 21'h0003ee; 
        10'b0011110000: data <= 21'h1ff011; 
        10'b0011110001: data <= 21'h1ffa99; 
        10'b0011110010: data <= 21'h1fff19; 
        10'b0011110011: data <= 21'h000210; 
        10'b0011110100: data <= 21'h1ff403; 
        10'b0011110101: data <= 21'h1ff469; 
        10'b0011110110: data <= 21'h1fed72; 
        10'b0011110111: data <= 21'h1fe7a5; 
        10'b0011111000: data <= 21'h1feca0; 
        10'b0011111001: data <= 21'h1ffb3e; 
        10'b0011111010: data <= 21'h000737; 
        10'b0011111011: data <= 21'h000980; 
        10'b0011111100: data <= 21'h000998; 
        10'b0011111101: data <= 21'h000237; 
        10'b0011111110: data <= 21'h0003ef; 
        10'b0011111111: data <= 21'h00035c; 
        10'b0100000000: data <= 21'h1fff65; 
        10'b0100000001: data <= 21'h1ffef0; 
        10'b0100000010: data <= 21'h1ff1c2; 
        10'b0100000011: data <= 21'h1ff283; 
        10'b0100000100: data <= 21'h1fe7e2; 
        10'b0100000101: data <= 21'h1fdb3c; 
        10'b0100000110: data <= 21'h1fde50; 
        10'b0100000111: data <= 21'h1ff2b0; 
        10'b0100001000: data <= 21'h1ff60f; 
        10'b0100001001: data <= 21'h00078e; 
        10'b0100001010: data <= 21'h0017ca; 
        10'b0100001011: data <= 21'h002213; 
        10'b0100001100: data <= 21'h000ca0; 
        10'b0100001101: data <= 21'h1fff1e; 
        10'b0100001110: data <= 21'h1ffa4f; 
        10'b0100001111: data <= 21'h1fe8e4; 
        10'b0100010000: data <= 21'h1fe393; 
        10'b0100010001: data <= 21'h1fe3f5; 
        10'b0100010010: data <= 21'h1fdcab; 
        10'b0100010011: data <= 21'h1fe163; 
        10'b0100010100: data <= 21'h1fef93; 
        10'b0100010101: data <= 21'h0001e8; 
        10'b0100010110: data <= 21'h0007ed; 
        10'b0100010111: data <= 21'h0005bf; 
        10'b0100011000: data <= 21'h0008be; 
        10'b0100011001: data <= 21'h0009af; 
        10'b0100011010: data <= 21'h000804; 
        10'b0100011011: data <= 21'h00010c; 
        10'b0100011100: data <= 21'h00068a; 
        10'b0100011101: data <= 21'h1ff86b; 
        10'b0100011110: data <= 21'h1ff288; 
        10'b0100011111: data <= 21'h1ff9c1; 
        10'b0100100000: data <= 21'h1fed4b; 
        10'b0100100001: data <= 21'h1fed06; 
        10'b0100100010: data <= 21'h1ff224; 
        10'b0100100011: data <= 21'h1ff6bc; 
        10'b0100100100: data <= 21'h1ff9c3; 
        10'b0100100101: data <= 21'h001300; 
        10'b0100100110: data <= 21'h003d7e; 
        10'b0100100111: data <= 21'h0040ec; 
        10'b0100101000: data <= 21'h001ed4; 
        10'b0100101001: data <= 21'h1fff55; 
        10'b0100101010: data <= 21'h1fed8c; 
        10'b0100101011: data <= 21'h1fe9c1; 
        10'b0100101100: data <= 21'h1fe512; 
        10'b0100101101: data <= 21'h1fe7b6; 
        10'b0100101110: data <= 21'h1fe91f; 
        10'b0100101111: data <= 21'h1ff1cb; 
        10'b0100110000: data <= 21'h1ffb3d; 
        10'b0100110001: data <= 21'h1fff2d; 
        10'b0100110010: data <= 21'h00083c; 
        10'b0100110011: data <= 21'h000361; 
        10'b0100110100: data <= 21'h0001a6; 
        10'b0100110101: data <= 21'h00017c; 
        10'b0100110110: data <= 21'h0006aa; 
        10'b0100110111: data <= 21'h000718; 
        10'b0100111000: data <= 21'h000007; 
        10'b0100111001: data <= 21'h1ffddb; 
        10'b0100111010: data <= 21'h1ffee2; 
        10'b0100111011: data <= 21'h1ff44e; 
        10'b0100111100: data <= 21'h1ff871; 
        10'b0100111101: data <= 21'h1ff454; 
        10'b0100111110: data <= 21'h1feed4; 
        10'b0100111111: data <= 21'h1fe610; 
        10'b0101000000: data <= 21'h1ffd07; 
        10'b0101000001: data <= 21'h00207f; 
        10'b0101000010: data <= 21'h004a23; 
        10'b0101000011: data <= 21'h004e8c; 
        10'b0101000100: data <= 21'h001d18; 
        10'b0101000101: data <= 21'h1ff9a3; 
        10'b0101000110: data <= 21'h1ffa26; 
        10'b0101000111: data <= 21'h1ff085; 
        10'b0101001000: data <= 21'h1fef9f; 
        10'b0101001001: data <= 21'h1ff0c9; 
        10'b0101001010: data <= 21'h1ff1ec; 
        10'b0101001011: data <= 21'h1ff969; 
        10'b0101001100: data <= 21'h1ffd36; 
        10'b0101001101: data <= 21'h000686; 
        10'b0101001110: data <= 21'h000926; 
        10'b0101001111: data <= 21'h00066e; 
        10'b0101010000: data <= 21'h000103; 
        10'b0101010001: data <= 21'h0008c1; 
        10'b0101010010: data <= 21'h000432; 
        10'b0101010011: data <= 21'h0002d7; 
        10'b0101010100: data <= 21'h0008f3; 
        10'b0101010101: data <= 21'h1ffe49; 
        10'b0101010110: data <= 21'h1ffd44; 
        10'b0101010111: data <= 21'h1ffc1f; 
        10'b0101011000: data <= 21'h1ff4db; 
        10'b0101011001: data <= 21'h1ff163; 
        10'b0101011010: data <= 21'h1fe10c; 
        10'b0101011011: data <= 21'h1fd495; 
        10'b0101011100: data <= 21'h1ffe9a; 
        10'b0101011101: data <= 21'h0020fc; 
        10'b0101011110: data <= 21'h005743; 
        10'b0101011111: data <= 21'h003c87; 
        10'b0101100000: data <= 21'h000bfc; 
        10'b0101100001: data <= 21'h000658; 
        10'b0101100010: data <= 21'h1ffc46; 
        10'b0101100011: data <= 21'h1fee51; 
        10'b0101100100: data <= 21'h1ff4d6; 
        10'b0101100101: data <= 21'h1ffa94; 
        10'b0101100110: data <= 21'h1ffcf3; 
        10'b0101100111: data <= 21'h1ffc3e; 
        10'b0101101000: data <= 21'h000092; 
        10'b0101101001: data <= 21'h0008e4; 
        10'b0101101010: data <= 21'h000156; 
        10'b0101101011: data <= 21'h000640; 
        10'b0101101100: data <= 21'h0000e5; 
        10'b0101101101: data <= 21'h0005f0; 
        10'b0101101110: data <= 21'h00058b; 
        10'b0101101111: data <= 21'h0005ea; 
        10'b0101110000: data <= 21'h0009dc; 
        10'b0101110001: data <= 21'h00000f; 
        10'b0101110010: data <= 21'h0000d5; 
        10'b0101110011: data <= 21'h1ffb96; 
        10'b0101110100: data <= 21'h1ffa0c; 
        10'b0101110101: data <= 21'h1fe7a6; 
        10'b0101110110: data <= 21'h1fcc59; 
        10'b0101110111: data <= 21'h1fcb9b; 
        10'b0101111000: data <= 21'h000012; 
        10'b0101111001: data <= 21'h001b84; 
        10'b0101111010: data <= 21'h0047e9; 
        10'b0101111011: data <= 21'h0028a3; 
        10'b0101111100: data <= 21'h000abe; 
        10'b0101111101: data <= 21'h000538; 
        10'b0101111110: data <= 21'h1fef97; 
        10'b0101111111: data <= 21'h1fe828; 
        10'b0110000000: data <= 21'h1ff758; 
        10'b0110000001: data <= 21'h1ffcf4; 
        10'b0110000010: data <= 21'h1ffcd3; 
        10'b0110000011: data <= 21'h1ffeda; 
        10'b0110000100: data <= 21'h000405; 
        10'b0110000101: data <= 21'h000602; 
        10'b0110000110: data <= 21'h0008ac; 
        10'b0110000111: data <= 21'h00059c; 
        10'b0110001000: data <= 21'h000461; 
        10'b0110001001: data <= 21'h00095c; 
        10'b0110001010: data <= 21'h000545; 
        10'b0110001011: data <= 21'h00077f; 
        10'b0110001100: data <= 21'h000787; 
        10'b0110001101: data <= 21'h1ffff8; 
        10'b0110001110: data <= 21'h00014a; 
        10'b0110001111: data <= 21'h1ffd1f; 
        10'b0110010000: data <= 21'h1fefe4; 
        10'b0110010001: data <= 21'h1fe458; 
        10'b0110010010: data <= 21'h1fcc89; 
        10'b0110010011: data <= 21'h1fd8f1; 
        10'b0110010100: data <= 21'h1fff21; 
        10'b0110010101: data <= 21'h001bee; 
        10'b0110010110: data <= 21'h003d55; 
        10'b0110010111: data <= 21'h00277f; 
        10'b0110011000: data <= 21'h000bce; 
        10'b0110011001: data <= 21'h1fea16; 
        10'b0110011010: data <= 21'h1fe250; 
        10'b0110011011: data <= 21'h1fe974; 
        10'b0110011100: data <= 21'h1ff2a9; 
        10'b0110011101: data <= 21'h1ffc24; 
        10'b0110011110: data <= 21'h1ffbce; 
        10'b0110011111: data <= 21'h1ffd22; 
        10'b0110100000: data <= 21'h0006af; 
        10'b0110100001: data <= 21'h000106; 
        10'b0110100010: data <= 21'h0001da; 
        10'b0110100011: data <= 21'h000554; 
        10'b0110100100: data <= 21'h0009ed; 
        10'b0110100101: data <= 21'h0001a1; 
        10'b0110100110: data <= 21'h00065d; 
        10'b0110100111: data <= 21'h000409; 
        10'b0110101000: data <= 21'h000247; 
        10'b0110101001: data <= 21'h0005c6; 
        10'b0110101010: data <= 21'h1ffa5f; 
        10'b0110101011: data <= 21'h1ff998; 
        10'b0110101100: data <= 21'h1ff5d9; 
        10'b0110101101: data <= 21'h1fe1c0; 
        10'b0110101110: data <= 21'h1fde15; 
        10'b0110101111: data <= 21'h1ff775; 
        10'b0110110000: data <= 21'h000c71; 
        10'b0110110001: data <= 21'h002743; 
        10'b0110110010: data <= 21'h0041a3; 
        10'b0110110011: data <= 21'h001736; 
        10'b0110110100: data <= 21'h000440; 
        10'b0110110101: data <= 21'h1fd6af; 
        10'b0110110110: data <= 21'h1fdb64; 
        10'b0110110111: data <= 21'h1fe998; 
        10'b0110111000: data <= 21'h1ff283; 
        10'b0110111001: data <= 21'h1ff651; 
        10'b0110111010: data <= 21'h1ffd8e; 
        10'b0110111011: data <= 21'h0000bd; 
        10'b0110111100: data <= 21'h00037f; 
        10'b0110111101: data <= 21'h00047b; 
        10'b0110111110: data <= 21'h00093d; 
        10'b0110111111: data <= 21'h00018a; 
        10'b0111000000: data <= 21'h00099c; 
        10'b0111000001: data <= 21'h0004b3; 
        10'b0111000010: data <= 21'h0008c8; 
        10'b0111000011: data <= 21'h00055a; 
        10'b0111000100: data <= 21'h0002d6; 
        10'b0111000101: data <= 21'h1ffc19; 
        10'b0111000110: data <= 21'h1ff715; 
        10'b0111000111: data <= 21'h1ff66b; 
        10'b0111001000: data <= 21'h1fe892; 
        10'b0111001001: data <= 21'h1ff1f9; 
        10'b0111001010: data <= 21'h1ff4d3; 
        10'b0111001011: data <= 21'h1ff9cd; 
        10'b0111001100: data <= 21'h1ffe6d; 
        10'b0111001101: data <= 21'h0033a4; 
        10'b0111001110: data <= 21'h003df6; 
        10'b0111001111: data <= 21'h00038d; 
        10'b0111010000: data <= 21'h1fecd2; 
        10'b0111010001: data <= 21'h1fd34e; 
        10'b0111010010: data <= 21'h1fdb06; 
        10'b0111010011: data <= 21'h1fe832; 
        10'b0111010100: data <= 21'h1fedeb; 
        10'b0111010101: data <= 21'h1ff84a; 
        10'b0111010110: data <= 21'h1ff82b; 
        10'b0111010111: data <= 21'h000018; 
        10'b0111011000: data <= 21'h1ffc8b; 
        10'b0111011001: data <= 21'h000089; 
        10'b0111011010: data <= 21'h00025b; 
        10'b0111011011: data <= 21'h0004fb; 
        10'b0111011100: data <= 21'h0003fc; 
        10'b0111011101: data <= 21'h00097c; 
        10'b0111011110: data <= 21'h00021b; 
        10'b0111011111: data <= 21'h00095b; 
        10'b0111100000: data <= 21'h0006eb; 
        10'b0111100001: data <= 21'h1ffa90; 
        10'b0111100010: data <= 21'h1fec60; 
        10'b0111100011: data <= 21'h1feabf; 
        10'b0111100100: data <= 21'h1ff0ca; 
        10'b0111100101: data <= 21'h1ff645; 
        10'b0111100110: data <= 21'h0006fc; 
        10'b0111100111: data <= 21'h000014; 
        10'b0111101000: data <= 21'h0010e0; 
        10'b0111101001: data <= 21'h003b25; 
        10'b0111101010: data <= 21'h0032ba; 
        10'b0111101011: data <= 21'h1ff5b3; 
        10'b0111101100: data <= 21'h1fdcc1; 
        10'b0111101101: data <= 21'h1fd324; 
        10'b0111101110: data <= 21'h1fdb41; 
        10'b0111101111: data <= 21'h1fe8c6; 
        10'b0111110000: data <= 21'h1ff744; 
        10'b0111110001: data <= 21'h1ffb9c; 
        10'b0111110010: data <= 21'h1ffcd9; 
        10'b0111110011: data <= 21'h1ffbc8; 
        10'b0111110100: data <= 21'h1ff8c3; 
        10'b0111110101: data <= 21'h000213; 
        10'b0111110110: data <= 21'h000587; 
        10'b0111110111: data <= 21'h000677; 
        10'b0111111000: data <= 21'h0005dd; 
        10'b0111111001: data <= 21'h000568; 
        10'b0111111010: data <= 21'h000353; 
        10'b0111111011: data <= 21'h0007d0; 
        10'b0111111100: data <= 21'h000455; 
        10'b0111111101: data <= 21'h1ff840; 
        10'b0111111110: data <= 21'h1feb12; 
        10'b0111111111: data <= 21'h1feb3c; 
        10'b1000000000: data <= 21'h1ff837; 
        10'b1000000001: data <= 21'h0007f6; 
        10'b1000000010: data <= 21'h000692; 
        10'b1000000011: data <= 21'h000a86; 
        10'b1000000100: data <= 21'h001b72; 
        10'b1000000101: data <= 21'h002c2e; 
        10'b1000000110: data <= 21'h001e8d; 
        10'b1000000111: data <= 21'h1febea; 
        10'b1000001000: data <= 21'h1fdf01; 
        10'b1000001001: data <= 21'h1fe3bb; 
        10'b1000001010: data <= 21'h1fe7dc; 
        10'b1000001011: data <= 21'h1fefd2; 
        10'b1000001100: data <= 21'h1ff80c; 
        10'b1000001101: data <= 21'h1ff28d; 
        10'b1000001110: data <= 21'h1ffa08; 
        10'b1000001111: data <= 21'h1ff6d6; 
        10'b1000010000: data <= 21'h1ffa66; 
        10'b1000010001: data <= 21'h000512; 
        10'b1000010010: data <= 21'h0008cb; 
        10'b1000010011: data <= 21'h0008fc; 
        10'b1000010100: data <= 21'h00093c; 
        10'b1000010101: data <= 21'h000682; 
        10'b1000010110: data <= 21'h0006c6; 
        10'b1000010111: data <= 21'h000780; 
        10'b1000011000: data <= 21'h0000e0; 
        10'b1000011001: data <= 21'h1ff45f; 
        10'b1000011010: data <= 21'h1fe608; 
        10'b1000011011: data <= 21'h1fee7a; 
        10'b1000011100: data <= 21'h1ff8d9; 
        10'b1000011101: data <= 21'h00041f; 
        10'b1000011110: data <= 21'h000211; 
        10'b1000011111: data <= 21'h000170; 
        10'b1000100000: data <= 21'h0003a3; 
        10'b1000100001: data <= 21'h001459; 
        10'b1000100010: data <= 21'h00047c; 
        10'b1000100011: data <= 21'h1fef64; 
        10'b1000100100: data <= 21'h1ff22b; 
        10'b1000100101: data <= 21'h1ff3f5; 
        10'b1000100110: data <= 21'h1ff0e0; 
        10'b1000100111: data <= 21'h1ff446; 
        10'b1000101000: data <= 21'h1feed5; 
        10'b1000101001: data <= 21'h1ff1b2; 
        10'b1000101010: data <= 21'h1ff75f; 
        10'b1000101011: data <= 21'h1ff865; 
        10'b1000101100: data <= 21'h00006a; 
        10'b1000101101: data <= 21'h0002ea; 
        10'b1000101110: data <= 21'h000333; 
        10'b1000101111: data <= 21'h000146; 
        10'b1000110000: data <= 21'h000179; 
        10'b1000110001: data <= 21'h0009b5; 
        10'b1000110010: data <= 21'h00053b; 
        10'b1000110011: data <= 21'h00035a; 
        10'b1000110100: data <= 21'h1ffd66; 
        10'b1000110101: data <= 21'h1ff7b9; 
        10'b1000110110: data <= 21'h1ffe72; 
        10'b1000110111: data <= 21'h1ffa4f; 
        10'b1000111000: data <= 21'h1fffdc; 
        10'b1000111001: data <= 21'h00026e; 
        10'b1000111010: data <= 21'h1ff99d; 
        10'b1000111011: data <= 21'h1ffdb3; 
        10'b1000111100: data <= 21'h1ff594; 
        10'b1000111101: data <= 21'h1ffc70; 
        10'b1000111110: data <= 21'h1ffd67; 
        10'b1000111111: data <= 21'h0000aa; 
        10'b1001000000: data <= 21'h0009e5; 
        10'b1001000001: data <= 21'h00038f; 
        10'b1001000010: data <= 21'h1ffc43; 
        10'b1001000011: data <= 21'h1ff21a; 
        10'b1001000100: data <= 21'h1feeed; 
        10'b1001000101: data <= 21'h1ff031; 
        10'b1001000110: data <= 21'h1ff396; 
        10'b1001000111: data <= 21'h1ffd34; 
        10'b1001001000: data <= 21'h000150; 
        10'b1001001001: data <= 21'h0007ee; 
        10'b1001001010: data <= 21'h00032a; 
        10'b1001001011: data <= 21'h0009c2; 
        10'b1001001100: data <= 21'h0006f0; 
        10'b1001001101: data <= 21'h0003a7; 
        10'b1001001110: data <= 21'h0005ac; 
        10'b1001001111: data <= 21'h0006ca; 
        10'b1001010000: data <= 21'h000565; 
        10'b1001010001: data <= 21'h000e8e; 
        10'b1001010010: data <= 21'h000bf7; 
        10'b1001010011: data <= 21'h0005a1; 
        10'b1001010100: data <= 21'h0000f0; 
        10'b1001010101: data <= 21'h1ffbdb; 
        10'b1001010110: data <= 21'h00002c; 
        10'b1001010111: data <= 21'h1ff79a; 
        10'b1001011000: data <= 21'h1fecec; 
        10'b1001011001: data <= 21'h1fea3a; 
        10'b1001011010: data <= 21'h1ffe0b; 
        10'b1001011011: data <= 21'h00068b; 
        10'b1001011100: data <= 21'h000a72; 
        10'b1001011101: data <= 21'h000be6; 
        10'b1001011110: data <= 21'h000835; 
        10'b1001011111: data <= 21'h1ff22e; 
        10'b1001100000: data <= 21'h1ff268; 
        10'b1001100001: data <= 21'h1ff07c; 
        10'b1001100010: data <= 21'h1ff553; 
        10'b1001100011: data <= 21'h1ff9d7; 
        10'b1001100100: data <= 21'h000161; 
        10'b1001100101: data <= 21'h000438; 
        10'b1001100110: data <= 21'h0000d4; 
        10'b1001100111: data <= 21'h000132; 
        10'b1001101000: data <= 21'h000564; 
        10'b1001101001: data <= 21'h000580; 
        10'b1001101010: data <= 21'h000633; 
        10'b1001101011: data <= 21'h000145; 
        10'b1001101100: data <= 21'h000c9d; 
        10'b1001101101: data <= 21'h001c27; 
        10'b1001101110: data <= 21'h001d29; 
        10'b1001101111: data <= 21'h001199; 
        10'b1001110000: data <= 21'h000265; 
        10'b1001110001: data <= 21'h1ffe0b; 
        10'b1001110010: data <= 21'h1ff951; 
        10'b1001110011: data <= 21'h1fe436; 
        10'b1001110100: data <= 21'h1fd2e2; 
        10'b1001110101: data <= 21'h1fdd82; 
        10'b1001110110: data <= 21'h00001b; 
        10'b1001110111: data <= 21'h0006c3; 
        10'b1001111000: data <= 21'h0019db; 
        10'b1001111001: data <= 21'h002a65; 
        10'b1001111010: data <= 21'h00128c; 
        10'b1001111011: data <= 21'h0003de; 
        10'b1001111100: data <= 21'h1ff673; 
        10'b1001111101: data <= 21'h1ff890; 
        10'b1001111110: data <= 21'h1fff56; 
        10'b1001111111: data <= 21'h000141; 
        10'b1010000000: data <= 21'h000099; 
        10'b1010000001: data <= 21'h00041c; 
        10'b1010000010: data <= 21'h000961; 
        10'b1010000011: data <= 21'h000484; 
        10'b1010000100: data <= 21'h0008ba; 
        10'b1010000101: data <= 21'h000575; 
        10'b1010000110: data <= 21'h0006fc; 
        10'b1010000111: data <= 21'h0003e3; 
        10'b1010001000: data <= 21'h000b43; 
        10'b1010001001: data <= 21'h001836; 
        10'b1010001010: data <= 21'h0019cc; 
        10'b1010001011: data <= 21'h000bd7; 
        10'b1010001100: data <= 21'h000343; 
        10'b1010001101: data <= 21'h1ff9ff; 
        10'b1010001110: data <= 21'h1ffbe9; 
        10'b1010001111: data <= 21'h1ff049; 
        10'b1010010000: data <= 21'h1ff508; 
        10'b1010010001: data <= 21'h1ff633; 
        10'b1010010010: data <= 21'h1ff2e7; 
        10'b1010010011: data <= 21'h000520; 
        10'b1010010100: data <= 21'h001e13; 
        10'b1010010101: data <= 21'h002446; 
        10'b1010010110: data <= 21'h00104c; 
        10'b1010010111: data <= 21'h1ffd1a; 
        10'b1010011000: data <= 21'h1ff912; 
        10'b1010011001: data <= 21'h1ff547; 
        10'b1010011010: data <= 21'h1ffc4e; 
        10'b1010011011: data <= 21'h1ffc98; 
        10'b1010011100: data <= 21'h000222; 
        10'b1010011101: data <= 21'h000113; 
        10'b1010011110: data <= 21'h000201; 
        10'b1010011111: data <= 21'h0000fd; 
        10'b1010100000: data <= 21'h000220; 
        10'b1010100001: data <= 21'h000159; 
        10'b1010100010: data <= 21'h00038a; 
        10'b1010100011: data <= 21'h00011c; 
        10'b1010100100: data <= 21'h00057f; 
        10'b1010100101: data <= 21'h000ab4; 
        10'b1010100110: data <= 21'h000b0e; 
        10'b1010100111: data <= 21'h1ffc6f; 
        10'b1010101000: data <= 21'h1feff6; 
        10'b1010101001: data <= 21'h1fefe2; 
        10'b1010101010: data <= 21'h1fe3a9; 
        10'b1010101011: data <= 21'h1fe4de; 
        10'b1010101100: data <= 21'h1fe7a8; 
        10'b1010101101: data <= 21'h1feb26; 
        10'b1010101110: data <= 21'h1feb3d; 
        10'b1010101111: data <= 21'h1feb31; 
        10'b1010110000: data <= 21'h1ff9fb; 
        10'b1010110001: data <= 21'h000285; 
        10'b1010110010: data <= 21'h000497; 
        10'b1010110011: data <= 21'h0006a7; 
        10'b1010110100: data <= 21'h000593; 
        10'b1010110101: data <= 21'h000158; 
        10'b1010110110: data <= 21'h0002e4; 
        10'b1010110111: data <= 21'h0007b9; 
        10'b1010111000: data <= 21'h000257; 
        10'b1010111001: data <= 21'h0003ce; 
        10'b1010111010: data <= 21'h000754; 
        10'b1010111011: data <= 21'h00026b; 
        10'b1010111100: data <= 21'h00097a; 
        10'b1010111101: data <= 21'h000305; 
        10'b1010111110: data <= 21'h00039d; 
        10'b1010111111: data <= 21'h00051e; 
        10'b1011000000: data <= 21'h000751; 
        10'b1011000001: data <= 21'h0006ac; 
        10'b1011000010: data <= 21'h00001a; 
        10'b1011000011: data <= 21'h1ffbdd; 
        10'b1011000100: data <= 21'h1ffe5c; 
        10'b1011000101: data <= 21'h1ffc30; 
        10'b1011000110: data <= 21'h1ff029; 
        10'b1011000111: data <= 21'h1fecb7; 
        10'b1011001000: data <= 21'h1ff1be; 
        10'b1011001001: data <= 21'h1fec01; 
        10'b1011001010: data <= 21'h1ff3c7; 
        10'b1011001011: data <= 21'h1ff086; 
        10'b1011001100: data <= 21'h1ff717; 
        10'b1011001101: data <= 21'h1ffe65; 
        10'b1011001110: data <= 21'h000315; 
        10'b1011001111: data <= 21'h000665; 
        10'b1011010000: data <= 21'h00009c; 
        10'b1011010001: data <= 21'h0005cf; 
        10'b1011010010: data <= 21'h000373; 
        10'b1011010011: data <= 21'h00084a; 
        10'b1011010100: data <= 21'h000216; 
        10'b1011010101: data <= 21'h000279; 
        10'b1011010110: data <= 21'h00038b; 
        10'b1011010111: data <= 21'h00030f; 
        10'b1011011000: data <= 21'h00037c; 
        10'b1011011001: data <= 21'h0006b6; 
        10'b1011011010: data <= 21'h0005f9; 
        10'b1011011011: data <= 21'h0001d3; 
        10'b1011011100: data <= 21'h000676; 
        10'b1011011101: data <= 21'h000898; 
        10'b1011011110: data <= 21'h0005d4; 
        10'b1011011111: data <= 21'h00055f; 
        10'b1011100000: data <= 21'h0007ad; 
        10'b1011100001: data <= 21'h00067f; 
        10'b1011100010: data <= 21'h0000e7; 
        10'b1011100011: data <= 21'h000549; 
        10'b1011100100: data <= 21'h0004d0; 
        10'b1011100101: data <= 21'h0002c9; 
        10'b1011100110: data <= 21'h1fffd6; 
        10'b1011100111: data <= 21'h000280; 
        10'b1011101000: data <= 21'h0005a2; 
        10'b1011101001: data <= 21'h0008b7; 
        10'b1011101010: data <= 21'h00066e; 
        10'b1011101011: data <= 21'h000107; 
        10'b1011101100: data <= 21'h0005fa; 
        10'b1011101101: data <= 21'h00059c; 
        10'b1011101110: data <= 21'h00055a; 
        10'b1011101111: data <= 21'h00028d; 
        10'b1011110000: data <= 21'h000240; 
        10'b1011110001: data <= 21'h00067b; 
        10'b1011110010: data <= 21'h0008dd; 
        10'b1011110011: data <= 21'h000732; 
        10'b1011110100: data <= 21'h00073b; 
        10'b1011110101: data <= 21'h000926; 
        10'b1011110110: data <= 21'h000172; 
        10'b1011110111: data <= 21'h000510; 
        10'b1011111000: data <= 21'h00099a; 
        10'b1011111001: data <= 21'h0007a1; 
        10'b1011111010: data <= 21'h0008a6; 
        10'b1011111011: data <= 21'h0007fb; 
        10'b1011111100: data <= 21'h0008a7; 
        10'b1011111101: data <= 21'h000416; 
        10'b1011111110: data <= 21'h000795; 
        10'b1011111111: data <= 21'h0007e0; 
        10'b1100000000: data <= 21'h0000ca; 
        10'b1100000001: data <= 21'h0001a5; 
        10'b1100000010: data <= 21'h00096b; 
        10'b1100000011: data <= 21'h000625; 
        10'b1100000100: data <= 21'h0005a9; 
        10'b1100000101: data <= 21'h0000d2; 
        10'b1100000110: data <= 21'h00041b; 
        10'b1100000111: data <= 21'h0001cf; 
        10'b1100001000: data <= 21'h0001af; 
        10'b1100001001: data <= 21'h000314; 
        10'b1100001010: data <= 21'h00058d; 
        10'b1100001011: data <= 21'h0007fe; 
        10'b1100001100: data <= 21'h0008de; 
        10'b1100001101: data <= 21'h0008a7; 
        10'b1100001110: data <= 21'h000887; 
        10'b1100001111: data <= 21'h0002d9; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 16) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 22'h000ff7; 
        10'b0000000001: data <= 22'h00079c; 
        10'b0000000010: data <= 22'h00087f; 
        10'b0000000011: data <= 22'h00037f; 
        10'b0000000100: data <= 22'h000d88; 
        10'b0000000101: data <= 22'h000d2c; 
        10'b0000000110: data <= 22'h000e8a; 
        10'b0000000111: data <= 22'h00039d; 
        10'b0000001000: data <= 22'h000cac; 
        10'b0000001001: data <= 22'h0003e1; 
        10'b0000001010: data <= 22'h000c0c; 
        10'b0000001011: data <= 22'h0009b9; 
        10'b0000001100: data <= 22'h000d91; 
        10'b0000001101: data <= 22'h00121a; 
        10'b0000001110: data <= 22'h000fea; 
        10'b0000001111: data <= 22'h000aea; 
        10'b0000010000: data <= 22'h000b14; 
        10'b0000010001: data <= 22'h0003e6; 
        10'b0000010010: data <= 22'h001294; 
        10'b0000010011: data <= 22'h00127a; 
        10'b0000010100: data <= 22'h000a8d; 
        10'b0000010101: data <= 22'h000d88; 
        10'b0000010110: data <= 22'h000a74; 
        10'b0000010111: data <= 22'h001037; 
        10'b0000011000: data <= 22'h00062b; 
        10'b0000011001: data <= 22'h001122; 
        10'b0000011010: data <= 22'h000a74; 
        10'b0000011011: data <= 22'h000f1b; 
        10'b0000011100: data <= 22'h0001f4; 
        10'b0000011101: data <= 22'h00100b; 
        10'b0000011110: data <= 22'h0004bb; 
        10'b0000011111: data <= 22'h000b6b; 
        10'b0000100000: data <= 22'h000a32; 
        10'b0000100001: data <= 22'h00040a; 
        10'b0000100010: data <= 22'h0005b1; 
        10'b0000100011: data <= 22'h000f12; 
        10'b0000100100: data <= 22'h000e79; 
        10'b0000100101: data <= 22'h000bc2; 
        10'b0000100110: data <= 22'h000ba3; 
        10'b0000100111: data <= 22'h000891; 
        10'b0000101000: data <= 22'h000dda; 
        10'b0000101001: data <= 22'h000f9e; 
        10'b0000101010: data <= 22'h001431; 
        10'b0000101011: data <= 22'h000a0c; 
        10'b0000101100: data <= 22'h000820; 
        10'b0000101101: data <= 22'h001039; 
        10'b0000101110: data <= 22'h000aeb; 
        10'b0000101111: data <= 22'h000769; 
        10'b0000110000: data <= 22'h001194; 
        10'b0000110001: data <= 22'h0010eb; 
        10'b0000110010: data <= 22'h0006ef; 
        10'b0000110011: data <= 22'h001224; 
        10'b0000110100: data <= 22'h00136f; 
        10'b0000110101: data <= 22'h000a4a; 
        10'b0000110110: data <= 22'h00108e; 
        10'b0000110111: data <= 22'h000d4f; 
        10'b0000111000: data <= 22'h001056; 
        10'b0000111001: data <= 22'h000c47; 
        10'b0000111010: data <= 22'h001391; 
        10'b0000111011: data <= 22'h0003cb; 
        10'b0000111100: data <= 22'h0003a6; 
        10'b0000111101: data <= 22'h000ce0; 
        10'b0000111110: data <= 22'h000985; 
        10'b0000111111: data <= 22'h000929; 
        10'b0001000000: data <= 22'h000629; 
        10'b0001000001: data <= 22'h000ac8; 
        10'b0001000010: data <= 22'h000045; 
        10'b0001000011: data <= 22'h00056a; 
        10'b0001000100: data <= 22'h0000b3; 
        10'b0001000101: data <= 22'h0004bd; 
        10'b0001000110: data <= 22'h0009ed; 
        10'b0001000111: data <= 22'h000ff1; 
        10'b0001001000: data <= 22'h000c11; 
        10'b0001001001: data <= 22'h000003; 
        10'b0001001010: data <= 22'h000beb; 
        10'b0001001011: data <= 22'h000725; 
        10'b0001001100: data <= 22'h000fac; 
        10'b0001001101: data <= 22'h0006cd; 
        10'b0001001110: data <= 22'h001140; 
        10'b0001001111: data <= 22'h000c8c; 
        10'b0001010000: data <= 22'h000d82; 
        10'b0001010001: data <= 22'h00024f; 
        10'b0001010010: data <= 22'h000eaf; 
        10'b0001010011: data <= 22'h000f08; 
        10'b0001010100: data <= 22'h0005d0; 
        10'b0001010101: data <= 22'h000685; 
        10'b0001010110: data <= 22'h000b01; 
        10'b0001010111: data <= 22'h000908; 
        10'b0001011000: data <= 22'h001260; 
        10'b0001011001: data <= 22'h0009ae; 
        10'b0001011010: data <= 22'h00021f; 
        10'b0001011011: data <= 22'h0011fe; 
        10'b0001011100: data <= 22'h3ffe04; 
        10'b0001011101: data <= 22'h3ffc5f; 
        10'b0001011110: data <= 22'h3ffc82; 
        10'b0001011111: data <= 22'h3ff5fe; 
        10'b0001100000: data <= 22'h3ffc75; 
        10'b0001100001: data <= 22'h000155; 
        10'b0001100010: data <= 22'h00077f; 
        10'b0001100011: data <= 22'h000efd; 
        10'b0001100100: data <= 22'h3ff891; 
        10'b0001100101: data <= 22'h3ffd49; 
        10'b0001100110: data <= 22'h3fff9f; 
        10'b0001100111: data <= 22'h3ff473; 
        10'b0001101000: data <= 22'h3ffece; 
        10'b0001101001: data <= 22'h0004c1; 
        10'b0001101010: data <= 22'h000bf9; 
        10'b0001101011: data <= 22'h000bb4; 
        10'b0001101100: data <= 22'h3ffdda; 
        10'b0001101101: data <= 22'h00109a; 
        10'b0001101110: data <= 22'h00063d; 
        10'b0001101111: data <= 22'h001187; 
        10'b0001110000: data <= 22'h000d7f; 
        10'b0001110001: data <= 22'h000830; 
        10'b0001110010: data <= 22'h001298; 
        10'b0001110011: data <= 22'h00126e; 
        10'b0001110100: data <= 22'h00020f; 
        10'b0001110101: data <= 22'h0003aa; 
        10'b0001110110: data <= 22'h00103c; 
        10'b0001110111: data <= 22'h000a55; 
        10'b0001111000: data <= 22'h0003ea; 
        10'b0001111001: data <= 22'h3fef07; 
        10'b0001111010: data <= 22'h00018f; 
        10'b0001111011: data <= 22'h0005f1; 
        10'b0001111100: data <= 22'h00093c; 
        10'b0001111101: data <= 22'h001084; 
        10'b0001111110: data <= 22'h00135d; 
        10'b0001111111: data <= 22'h00279a; 
        10'b0010000000: data <= 22'h000ad2; 
        10'b0010000001: data <= 22'h3ff7ad; 
        10'b0010000010: data <= 22'h3ff6ef; 
        10'b0010000011: data <= 22'h000627; 
        10'b0010000100: data <= 22'h0015e9; 
        10'b0010000101: data <= 22'h00188c; 
        10'b0010000110: data <= 22'h00186f; 
        10'b0010000111: data <= 22'h001c9e; 
        10'b0010001000: data <= 22'h000ef6; 
        10'b0010001001: data <= 22'h000716; 
        10'b0010001010: data <= 22'h000633; 
        10'b0010001011: data <= 22'h0006d3; 
        10'b0010001100: data <= 22'h000272; 
        10'b0010001101: data <= 22'h000ffb; 
        10'b0010001110: data <= 22'h000320; 
        10'b0010001111: data <= 22'h000b3e; 
        10'b0010010000: data <= 22'h0002d0; 
        10'b0010010001: data <= 22'h000ac7; 
        10'b0010010010: data <= 22'h00033c; 
        10'b0010010011: data <= 22'h3ffbd2; 
        10'b0010010100: data <= 22'h3fdc5b; 
        10'b0010010101: data <= 22'h3fdc0f; 
        10'b0010010110: data <= 22'h3fef88; 
        10'b0010010111: data <= 22'h000038; 
        10'b0010011000: data <= 22'h000d80; 
        10'b0010011001: data <= 22'h000f32; 
        10'b0010011010: data <= 22'h001a68; 
        10'b0010011011: data <= 22'h001484; 
        10'b0010011100: data <= 22'h000c23; 
        10'b0010011101: data <= 22'h3fec0b; 
        10'b0010011110: data <= 22'h3ffdff; 
        10'b0010011111: data <= 22'h00042e; 
        10'b0010100000: data <= 22'h001383; 
        10'b0010100001: data <= 22'h001f69; 
        10'b0010100010: data <= 22'h003445; 
        10'b0010100011: data <= 22'h00209e; 
        10'b0010100100: data <= 22'h001ab6; 
        10'b0010100101: data <= 22'h3ff920; 
        10'b0010100110: data <= 22'h000761; 
        10'b0010100111: data <= 22'h000414; 
        10'b0010101000: data <= 22'h000368; 
        10'b0010101001: data <= 22'h000b97; 
        10'b0010101010: data <= 22'h000220; 
        10'b0010101011: data <= 22'h000908; 
        10'b0010101100: data <= 22'h00021d; 
        10'b0010101101: data <= 22'h3ffaae; 
        10'b0010101110: data <= 22'h3fec62; 
        10'b0010101111: data <= 22'h3fec9f; 
        10'b0010110000: data <= 22'h3fd36f; 
        10'b0010110001: data <= 22'h3fca26; 
        10'b0010110010: data <= 22'h3fde45; 
        10'b0010110011: data <= 22'h3ff816; 
        10'b0010110100: data <= 22'h3ff7c1; 
        10'b0010110101: data <= 22'h3fef10; 
        10'b0010110110: data <= 22'h3ff835; 
        10'b0010110111: data <= 22'h3fd956; 
        10'b0010111000: data <= 22'h3fd66c; 
        10'b0010111001: data <= 22'h3fd61b; 
        10'b0010111010: data <= 22'h3fee7b; 
        10'b0010111011: data <= 22'h3ff30b; 
        10'b0010111100: data <= 22'h00139a; 
        10'b0010111101: data <= 22'h002047; 
        10'b0010111110: data <= 22'h001def; 
        10'b0010111111: data <= 22'h001930; 
        10'b0011000000: data <= 22'h000690; 
        10'b0011000001: data <= 22'h3ffaa5; 
        10'b0011000010: data <= 22'h000071; 
        10'b0011000011: data <= 22'h000971; 
        10'b0011000100: data <= 22'h0007a3; 
        10'b0011000101: data <= 22'h00044e; 
        10'b0011000110: data <= 22'h000558; 
        10'b0011000111: data <= 22'h000133; 
        10'b0011001000: data <= 22'h000ca7; 
        10'b0011001001: data <= 22'h3ffd4b; 
        10'b0011001010: data <= 22'h3fed31; 
        10'b0011001011: data <= 22'h3fd986; 
        10'b0011001100: data <= 22'h3fc3dc; 
        10'b0011001101: data <= 22'h3fb36b; 
        10'b0011001110: data <= 22'h3fcc01; 
        10'b0011001111: data <= 22'h3fe946; 
        10'b0011010000: data <= 22'h3feb31; 
        10'b0011010001: data <= 22'h3fe212; 
        10'b0011010010: data <= 22'h3fdb01; 
        10'b0011010011: data <= 22'h3fc67b; 
        10'b0011010100: data <= 22'h3fcdc3; 
        10'b0011010101: data <= 22'h3fd0da; 
        10'b0011010110: data <= 22'h3fd582; 
        10'b0011010111: data <= 22'h3ffe8e; 
        10'b0011011000: data <= 22'h0008ea; 
        10'b0011011001: data <= 22'h000589; 
        10'b0011011010: data <= 22'h000547; 
        10'b0011011011: data <= 22'h3fefd2; 
        10'b0011011100: data <= 22'h3fe9ee; 
        10'b0011011101: data <= 22'h3ff72e; 
        10'b0011011110: data <= 22'h00072c; 
        10'b0011011111: data <= 22'h00085f; 
        10'b0011100000: data <= 22'h000949; 
        10'b0011100001: data <= 22'h0007da; 
        10'b0011100010: data <= 22'h0007b5; 
        10'b0011100011: data <= 22'h001060; 
        10'b0011100100: data <= 22'h00053c; 
        10'b0011100101: data <= 22'h3fff78; 
        10'b0011100110: data <= 22'h3fe9a2; 
        10'b0011100111: data <= 22'h3fde18; 
        10'b0011101000: data <= 22'h3fb9e9; 
        10'b0011101001: data <= 22'h3fb3e7; 
        10'b0011101010: data <= 22'h3fb78e; 
        10'b0011101011: data <= 22'h3fd904; 
        10'b0011101100: data <= 22'h3fee1b; 
        10'b0011101101: data <= 22'h3fe9fd; 
        10'b0011101110: data <= 22'h3fee08; 
        10'b0011101111: data <= 22'h0007dd; 
        10'b0011110000: data <= 22'h3fe022; 
        10'b0011110001: data <= 22'h3ff532; 
        10'b0011110010: data <= 22'h3ffe33; 
        10'b0011110011: data <= 22'h000421; 
        10'b0011110100: data <= 22'h3fe806; 
        10'b0011110101: data <= 22'h3fe8d2; 
        10'b0011110110: data <= 22'h3fdae4; 
        10'b0011110111: data <= 22'h3fcf4a; 
        10'b0011111000: data <= 22'h3fd941; 
        10'b0011111001: data <= 22'h3ff67d; 
        10'b0011111010: data <= 22'h000e6f; 
        10'b0011111011: data <= 22'h001300; 
        10'b0011111100: data <= 22'h001330; 
        10'b0011111101: data <= 22'h00046e; 
        10'b0011111110: data <= 22'h0007de; 
        10'b0011111111: data <= 22'h0006b8; 
        10'b0100000000: data <= 22'h3ffeca; 
        10'b0100000001: data <= 22'h3ffde1; 
        10'b0100000010: data <= 22'h3fe385; 
        10'b0100000011: data <= 22'h3fe507; 
        10'b0100000100: data <= 22'h3fcfc4; 
        10'b0100000101: data <= 22'h3fb678; 
        10'b0100000110: data <= 22'h3fbca1; 
        10'b0100000111: data <= 22'h3fe561; 
        10'b0100001000: data <= 22'h3fec1d; 
        10'b0100001001: data <= 22'h000f1c; 
        10'b0100001010: data <= 22'h002f94; 
        10'b0100001011: data <= 22'h004426; 
        10'b0100001100: data <= 22'h001940; 
        10'b0100001101: data <= 22'h3ffe3d; 
        10'b0100001110: data <= 22'h3ff49d; 
        10'b0100001111: data <= 22'h3fd1c8; 
        10'b0100010000: data <= 22'h3fc726; 
        10'b0100010001: data <= 22'h3fc7ea; 
        10'b0100010010: data <= 22'h3fb957; 
        10'b0100010011: data <= 22'h3fc2c6; 
        10'b0100010100: data <= 22'h3fdf27; 
        10'b0100010101: data <= 22'h0003d0; 
        10'b0100010110: data <= 22'h000fda; 
        10'b0100010111: data <= 22'h000b7e; 
        10'b0100011000: data <= 22'h00117c; 
        10'b0100011001: data <= 22'h00135e; 
        10'b0100011010: data <= 22'h001008; 
        10'b0100011011: data <= 22'h000219; 
        10'b0100011100: data <= 22'h000d15; 
        10'b0100011101: data <= 22'h3ff0d6; 
        10'b0100011110: data <= 22'h3fe510; 
        10'b0100011111: data <= 22'h3ff383; 
        10'b0100100000: data <= 22'h3fda95; 
        10'b0100100001: data <= 22'h3fda0c; 
        10'b0100100010: data <= 22'h3fe448; 
        10'b0100100011: data <= 22'h3fed79; 
        10'b0100100100: data <= 22'h3ff385; 
        10'b0100100101: data <= 22'h002600; 
        10'b0100100110: data <= 22'h007afc; 
        10'b0100100111: data <= 22'h0081d8; 
        10'b0100101000: data <= 22'h003da8; 
        10'b0100101001: data <= 22'h3ffeaa; 
        10'b0100101010: data <= 22'h3fdb18; 
        10'b0100101011: data <= 22'h3fd382; 
        10'b0100101100: data <= 22'h3fca25; 
        10'b0100101101: data <= 22'h3fcf6c; 
        10'b0100101110: data <= 22'h3fd23d; 
        10'b0100101111: data <= 22'h3fe395; 
        10'b0100110000: data <= 22'h3ff67b; 
        10'b0100110001: data <= 22'h3ffe59; 
        10'b0100110010: data <= 22'h001078; 
        10'b0100110011: data <= 22'h0006c2; 
        10'b0100110100: data <= 22'h00034c; 
        10'b0100110101: data <= 22'h0002f8; 
        10'b0100110110: data <= 22'h000d54; 
        10'b0100110111: data <= 22'h000e31; 
        10'b0100111000: data <= 22'h00000d; 
        10'b0100111001: data <= 22'h3ffbb6; 
        10'b0100111010: data <= 22'h3ffdc4; 
        10'b0100111011: data <= 22'h3fe89b; 
        10'b0100111100: data <= 22'h3ff0e1; 
        10'b0100111101: data <= 22'h3fe8a7; 
        10'b0100111110: data <= 22'h3fdda8; 
        10'b0100111111: data <= 22'h3fcc1f; 
        10'b0101000000: data <= 22'h3ffa0e; 
        10'b0101000001: data <= 22'h0040fe; 
        10'b0101000010: data <= 22'h009446; 
        10'b0101000011: data <= 22'h009d18; 
        10'b0101000100: data <= 22'h003a30; 
        10'b0101000101: data <= 22'h3ff347; 
        10'b0101000110: data <= 22'h3ff44c; 
        10'b0101000111: data <= 22'h3fe10a; 
        10'b0101001000: data <= 22'h3fdf3d; 
        10'b0101001001: data <= 22'h3fe193; 
        10'b0101001010: data <= 22'h3fe3d8; 
        10'b0101001011: data <= 22'h3ff2d2; 
        10'b0101001100: data <= 22'h3ffa6b; 
        10'b0101001101: data <= 22'h000d0b; 
        10'b0101001110: data <= 22'h00124b; 
        10'b0101001111: data <= 22'h000cdc; 
        10'b0101010000: data <= 22'h000206; 
        10'b0101010001: data <= 22'h001182; 
        10'b0101010010: data <= 22'h000864; 
        10'b0101010011: data <= 22'h0005af; 
        10'b0101010100: data <= 22'h0011e6; 
        10'b0101010101: data <= 22'h3ffc92; 
        10'b0101010110: data <= 22'h3ffa88; 
        10'b0101010111: data <= 22'h3ff83e; 
        10'b0101011000: data <= 22'h3fe9b6; 
        10'b0101011001: data <= 22'h3fe2c6; 
        10'b0101011010: data <= 22'h3fc218; 
        10'b0101011011: data <= 22'h3fa92a; 
        10'b0101011100: data <= 22'h3ffd35; 
        10'b0101011101: data <= 22'h0041f9; 
        10'b0101011110: data <= 22'h00ae86; 
        10'b0101011111: data <= 22'h00790d; 
        10'b0101100000: data <= 22'h0017f8; 
        10'b0101100001: data <= 22'h000caf; 
        10'b0101100010: data <= 22'h3ff88b; 
        10'b0101100011: data <= 22'h3fdca2; 
        10'b0101100100: data <= 22'h3fe9ac; 
        10'b0101100101: data <= 22'h3ff529; 
        10'b0101100110: data <= 22'h3ff9e7; 
        10'b0101100111: data <= 22'h3ff87c; 
        10'b0101101000: data <= 22'h000124; 
        10'b0101101001: data <= 22'h0011c7; 
        10'b0101101010: data <= 22'h0002ab; 
        10'b0101101011: data <= 22'h000c80; 
        10'b0101101100: data <= 22'h0001ca; 
        10'b0101101101: data <= 22'h000be1; 
        10'b0101101110: data <= 22'h000b15; 
        10'b0101101111: data <= 22'h000bd5; 
        10'b0101110000: data <= 22'h0013b8; 
        10'b0101110001: data <= 22'h00001e; 
        10'b0101110010: data <= 22'h0001aa; 
        10'b0101110011: data <= 22'h3ff72c; 
        10'b0101110100: data <= 22'h3ff417; 
        10'b0101110101: data <= 22'h3fcf4c; 
        10'b0101110110: data <= 22'h3f98b2; 
        10'b0101110111: data <= 22'h3f9735; 
        10'b0101111000: data <= 22'h000024; 
        10'b0101111001: data <= 22'h003708; 
        10'b0101111010: data <= 22'h008fd3; 
        10'b0101111011: data <= 22'h005146; 
        10'b0101111100: data <= 22'h00157c; 
        10'b0101111101: data <= 22'h000a6f; 
        10'b0101111110: data <= 22'h3fdf2e; 
        10'b0101111111: data <= 22'h3fd04f; 
        10'b0110000000: data <= 22'h3feeaf; 
        10'b0110000001: data <= 22'h3ff9e8; 
        10'b0110000010: data <= 22'h3ff9a6; 
        10'b0110000011: data <= 22'h3ffdb5; 
        10'b0110000100: data <= 22'h00080b; 
        10'b0110000101: data <= 22'h000c05; 
        10'b0110000110: data <= 22'h001157; 
        10'b0110000111: data <= 22'h000b38; 
        10'b0110001000: data <= 22'h0008c1; 
        10'b0110001001: data <= 22'h0012b9; 
        10'b0110001010: data <= 22'h000a89; 
        10'b0110001011: data <= 22'h000efe; 
        10'b0110001100: data <= 22'h000f0e; 
        10'b0110001101: data <= 22'h3ffff0; 
        10'b0110001110: data <= 22'h000294; 
        10'b0110001111: data <= 22'h3ffa3f; 
        10'b0110010000: data <= 22'h3fdfc8; 
        10'b0110010001: data <= 22'h3fc8b0; 
        10'b0110010010: data <= 22'h3f9912; 
        10'b0110010011: data <= 22'h3fb1e2; 
        10'b0110010100: data <= 22'h3ffe42; 
        10'b0110010101: data <= 22'h0037db; 
        10'b0110010110: data <= 22'h007aab; 
        10'b0110010111: data <= 22'h004efe; 
        10'b0110011000: data <= 22'h00179c; 
        10'b0110011001: data <= 22'h3fd42c; 
        10'b0110011010: data <= 22'h3fc4a0; 
        10'b0110011011: data <= 22'h3fd2e8; 
        10'b0110011100: data <= 22'h3fe552; 
        10'b0110011101: data <= 22'h3ff849; 
        10'b0110011110: data <= 22'h3ff79d; 
        10'b0110011111: data <= 22'h3ffa45; 
        10'b0110100000: data <= 22'h000d5e; 
        10'b0110100001: data <= 22'h00020c; 
        10'b0110100010: data <= 22'h0003b3; 
        10'b0110100011: data <= 22'h000aa7; 
        10'b0110100100: data <= 22'h0013da; 
        10'b0110100101: data <= 22'h000342; 
        10'b0110100110: data <= 22'h000cbb; 
        10'b0110100111: data <= 22'h000811; 
        10'b0110101000: data <= 22'h00048e; 
        10'b0110101001: data <= 22'h000b8d; 
        10'b0110101010: data <= 22'h3ff4be; 
        10'b0110101011: data <= 22'h3ff32f; 
        10'b0110101100: data <= 22'h3febb1; 
        10'b0110101101: data <= 22'h3fc380; 
        10'b0110101110: data <= 22'h3fbc2a; 
        10'b0110101111: data <= 22'h3feee9; 
        10'b0110110000: data <= 22'h0018e3; 
        10'b0110110001: data <= 22'h004e87; 
        10'b0110110010: data <= 22'h008345; 
        10'b0110110011: data <= 22'h002e6d; 
        10'b0110110100: data <= 22'h000880; 
        10'b0110110101: data <= 22'h3fad5e; 
        10'b0110110110: data <= 22'h3fb6c9; 
        10'b0110110111: data <= 22'h3fd32f; 
        10'b0110111000: data <= 22'h3fe506; 
        10'b0110111001: data <= 22'h3feca2; 
        10'b0110111010: data <= 22'h3ffb1d; 
        10'b0110111011: data <= 22'h000179; 
        10'b0110111100: data <= 22'h0006fe; 
        10'b0110111101: data <= 22'h0008f6; 
        10'b0110111110: data <= 22'h001279; 
        10'b0110111111: data <= 22'h000315; 
        10'b0111000000: data <= 22'h001337; 
        10'b0111000001: data <= 22'h000965; 
        10'b0111000010: data <= 22'h00118f; 
        10'b0111000011: data <= 22'h000ab4; 
        10'b0111000100: data <= 22'h0005ac; 
        10'b0111000101: data <= 22'h3ff833; 
        10'b0111000110: data <= 22'h3fee2a; 
        10'b0111000111: data <= 22'h3fecd6; 
        10'b0111001000: data <= 22'h3fd123; 
        10'b0111001001: data <= 22'h3fe3f1; 
        10'b0111001010: data <= 22'h3fe9a7; 
        10'b0111001011: data <= 22'h3ff399; 
        10'b0111001100: data <= 22'h3ffcda; 
        10'b0111001101: data <= 22'h006748; 
        10'b0111001110: data <= 22'h007beb; 
        10'b0111001111: data <= 22'h00071a; 
        10'b0111010000: data <= 22'h3fd9a3; 
        10'b0111010001: data <= 22'h3fa69b; 
        10'b0111010010: data <= 22'h3fb60c; 
        10'b0111010011: data <= 22'h3fd063; 
        10'b0111010100: data <= 22'h3fdbd5; 
        10'b0111010101: data <= 22'h3ff093; 
        10'b0111010110: data <= 22'h3ff057; 
        10'b0111010111: data <= 22'h000031; 
        10'b0111011000: data <= 22'h3ff916; 
        10'b0111011001: data <= 22'h000113; 
        10'b0111011010: data <= 22'h0004b5; 
        10'b0111011011: data <= 22'h0009f7; 
        10'b0111011100: data <= 22'h0007f7; 
        10'b0111011101: data <= 22'h0012f9; 
        10'b0111011110: data <= 22'h000437; 
        10'b0111011111: data <= 22'h0012b7; 
        10'b0111100000: data <= 22'h000dd5; 
        10'b0111100001: data <= 22'h3ff520; 
        10'b0111100010: data <= 22'h3fd8c1; 
        10'b0111100011: data <= 22'h3fd57e; 
        10'b0111100100: data <= 22'h3fe193; 
        10'b0111100101: data <= 22'h3fec8a; 
        10'b0111100110: data <= 22'h000df8; 
        10'b0111100111: data <= 22'h000028; 
        10'b0111101000: data <= 22'h0021bf; 
        10'b0111101001: data <= 22'h00764b; 
        10'b0111101010: data <= 22'h006574; 
        10'b0111101011: data <= 22'h3feb66; 
        10'b0111101100: data <= 22'h3fb981; 
        10'b0111101101: data <= 22'h3fa649; 
        10'b0111101110: data <= 22'h3fb681; 
        10'b0111101111: data <= 22'h3fd18b; 
        10'b0111110000: data <= 22'h3fee88; 
        10'b0111110001: data <= 22'h3ff739; 
        10'b0111110010: data <= 22'h3ff9b3; 
        10'b0111110011: data <= 22'h3ff790; 
        10'b0111110100: data <= 22'h3ff187; 
        10'b0111110101: data <= 22'h000427; 
        10'b0111110110: data <= 22'h000b0f; 
        10'b0111110111: data <= 22'h000cef; 
        10'b0111111000: data <= 22'h000bbb; 
        10'b0111111001: data <= 22'h000ad0; 
        10'b0111111010: data <= 22'h0006a5; 
        10'b0111111011: data <= 22'h000fa0; 
        10'b0111111100: data <= 22'h0008ab; 
        10'b0111111101: data <= 22'h3ff080; 
        10'b0111111110: data <= 22'h3fd624; 
        10'b0111111111: data <= 22'h3fd677; 
        10'b1000000000: data <= 22'h3ff06d; 
        10'b1000000001: data <= 22'h000fec; 
        10'b1000000010: data <= 22'h000d24; 
        10'b1000000011: data <= 22'h00150c; 
        10'b1000000100: data <= 22'h0036e4; 
        10'b1000000101: data <= 22'h00585c; 
        10'b1000000110: data <= 22'h003d19; 
        10'b1000000111: data <= 22'h3fd7d5; 
        10'b1000001000: data <= 22'h3fbe01; 
        10'b1000001001: data <= 22'h3fc776; 
        10'b1000001010: data <= 22'h3fcfb8; 
        10'b1000001011: data <= 22'h3fdfa4; 
        10'b1000001100: data <= 22'h3ff019; 
        10'b1000001101: data <= 22'h3fe51b; 
        10'b1000001110: data <= 22'h3ff410; 
        10'b1000001111: data <= 22'h3fedac; 
        10'b1000010000: data <= 22'h3ff4cd; 
        10'b1000010001: data <= 22'h000a23; 
        10'b1000010010: data <= 22'h001197; 
        10'b1000010011: data <= 22'h0011f8; 
        10'b1000010100: data <= 22'h001278; 
        10'b1000010101: data <= 22'h000d03; 
        10'b1000010110: data <= 22'h000d8c; 
        10'b1000010111: data <= 22'h000f01; 
        10'b1000011000: data <= 22'h0001c0; 
        10'b1000011001: data <= 22'h3fe8be; 
        10'b1000011010: data <= 22'h3fcc0f; 
        10'b1000011011: data <= 22'h3fdcf4; 
        10'b1000011100: data <= 22'h3ff1b1; 
        10'b1000011101: data <= 22'h00083f; 
        10'b1000011110: data <= 22'h000423; 
        10'b1000011111: data <= 22'h0002df; 
        10'b1000100000: data <= 22'h000746; 
        10'b1000100001: data <= 22'h0028b1; 
        10'b1000100010: data <= 22'h0008f7; 
        10'b1000100011: data <= 22'h3fdec9; 
        10'b1000100100: data <= 22'h3fe456; 
        10'b1000100101: data <= 22'h3fe7eb; 
        10'b1000100110: data <= 22'h3fe1c1; 
        10'b1000100111: data <= 22'h3fe88b; 
        10'b1000101000: data <= 22'h3fddaa; 
        10'b1000101001: data <= 22'h3fe365; 
        10'b1000101010: data <= 22'h3feebe; 
        10'b1000101011: data <= 22'h3ff0cb; 
        10'b1000101100: data <= 22'h0000d4; 
        10'b1000101101: data <= 22'h0005d4; 
        10'b1000101110: data <= 22'h000666; 
        10'b1000101111: data <= 22'h00028d; 
        10'b1000110000: data <= 22'h0002f1; 
        10'b1000110001: data <= 22'h00136b; 
        10'b1000110010: data <= 22'h000a77; 
        10'b1000110011: data <= 22'h0006b4; 
        10'b1000110100: data <= 22'h3ffacb; 
        10'b1000110101: data <= 22'h3fef72; 
        10'b1000110110: data <= 22'h3ffce4; 
        10'b1000110111: data <= 22'h3ff49d; 
        10'b1000111000: data <= 22'h3fffb8; 
        10'b1000111001: data <= 22'h0004dd; 
        10'b1000111010: data <= 22'h3ff33a; 
        10'b1000111011: data <= 22'h3ffb66; 
        10'b1000111100: data <= 22'h3feb27; 
        10'b1000111101: data <= 22'h3ff8e0; 
        10'b1000111110: data <= 22'h3fface; 
        10'b1000111111: data <= 22'h000154; 
        10'b1001000000: data <= 22'h0013ca; 
        10'b1001000001: data <= 22'h00071d; 
        10'b1001000010: data <= 22'h3ff886; 
        10'b1001000011: data <= 22'h3fe435; 
        10'b1001000100: data <= 22'h3fddda; 
        10'b1001000101: data <= 22'h3fe062; 
        10'b1001000110: data <= 22'h3fe72b; 
        10'b1001000111: data <= 22'h3ffa68; 
        10'b1001001000: data <= 22'h0002a0; 
        10'b1001001001: data <= 22'h000fdb; 
        10'b1001001010: data <= 22'h000655; 
        10'b1001001011: data <= 22'h001385; 
        10'b1001001100: data <= 22'h000ddf; 
        10'b1001001101: data <= 22'h00074e; 
        10'b1001001110: data <= 22'h000b59; 
        10'b1001001111: data <= 22'h000d94; 
        10'b1001010000: data <= 22'h000ac9; 
        10'b1001010001: data <= 22'h001d1d; 
        10'b1001010010: data <= 22'h0017ef; 
        10'b1001010011: data <= 22'h000b42; 
        10'b1001010100: data <= 22'h0001e0; 
        10'b1001010101: data <= 22'h3ff7b7; 
        10'b1001010110: data <= 22'h000059; 
        10'b1001010111: data <= 22'h3fef34; 
        10'b1001011000: data <= 22'h3fd9d9; 
        10'b1001011001: data <= 22'h3fd475; 
        10'b1001011010: data <= 22'h3ffc15; 
        10'b1001011011: data <= 22'h000d16; 
        10'b1001011100: data <= 22'h0014e4; 
        10'b1001011101: data <= 22'h0017cb; 
        10'b1001011110: data <= 22'h001069; 
        10'b1001011111: data <= 22'h3fe45c; 
        10'b1001100000: data <= 22'h3fe4cf; 
        10'b1001100001: data <= 22'h3fe0f8; 
        10'b1001100010: data <= 22'h3feaa6; 
        10'b1001100011: data <= 22'h3ff3ae; 
        10'b1001100100: data <= 22'h0002c3; 
        10'b1001100101: data <= 22'h000870; 
        10'b1001100110: data <= 22'h0001a8; 
        10'b1001100111: data <= 22'h000264; 
        10'b1001101000: data <= 22'h000ac8; 
        10'b1001101001: data <= 22'h000b00; 
        10'b1001101010: data <= 22'h000c66; 
        10'b1001101011: data <= 22'h00028a; 
        10'b1001101100: data <= 22'h001939; 
        10'b1001101101: data <= 22'h00384f; 
        10'b1001101110: data <= 22'h003a52; 
        10'b1001101111: data <= 22'h002332; 
        10'b1001110000: data <= 22'h0004ca; 
        10'b1001110001: data <= 22'h3ffc16; 
        10'b1001110010: data <= 22'h3ff2a2; 
        10'b1001110011: data <= 22'h3fc86b; 
        10'b1001110100: data <= 22'h3fa5c4; 
        10'b1001110101: data <= 22'h3fbb03; 
        10'b1001110110: data <= 22'h000035; 
        10'b1001110111: data <= 22'h000d85; 
        10'b1001111000: data <= 22'h0033b6; 
        10'b1001111001: data <= 22'h0054c9; 
        10'b1001111010: data <= 22'h002518; 
        10'b1001111011: data <= 22'h0007bb; 
        10'b1001111100: data <= 22'h3fece6; 
        10'b1001111101: data <= 22'h3ff120; 
        10'b1001111110: data <= 22'h3ffeac; 
        10'b1001111111: data <= 22'h000282; 
        10'b1010000000: data <= 22'h000131; 
        10'b1010000001: data <= 22'h000839; 
        10'b1010000010: data <= 22'h0012c3; 
        10'b1010000011: data <= 22'h000908; 
        10'b1010000100: data <= 22'h001174; 
        10'b1010000101: data <= 22'h000aea; 
        10'b1010000110: data <= 22'h000df8; 
        10'b1010000111: data <= 22'h0007c5; 
        10'b1010001000: data <= 22'h001686; 
        10'b1010001001: data <= 22'h00306c; 
        10'b1010001010: data <= 22'h003397; 
        10'b1010001011: data <= 22'h0017ad; 
        10'b1010001100: data <= 22'h000685; 
        10'b1010001101: data <= 22'h3ff3fd; 
        10'b1010001110: data <= 22'h3ff7d2; 
        10'b1010001111: data <= 22'h3fe091; 
        10'b1010010000: data <= 22'h3fea10; 
        10'b1010010001: data <= 22'h3fec66; 
        10'b1010010010: data <= 22'h3fe5cd; 
        10'b1010010011: data <= 22'h000a41; 
        10'b1010010100: data <= 22'h003c26; 
        10'b1010010101: data <= 22'h00488c; 
        10'b1010010110: data <= 22'h002098; 
        10'b1010010111: data <= 22'h3ffa34; 
        10'b1010011000: data <= 22'h3ff224; 
        10'b1010011001: data <= 22'h3fea8e; 
        10'b1010011010: data <= 22'h3ff89c; 
        10'b1010011011: data <= 22'h3ff930; 
        10'b1010011100: data <= 22'h000444; 
        10'b1010011101: data <= 22'h000227; 
        10'b1010011110: data <= 22'h000402; 
        10'b1010011111: data <= 22'h0001fb; 
        10'b1010100000: data <= 22'h000440; 
        10'b1010100001: data <= 22'h0002b1; 
        10'b1010100010: data <= 22'h000714; 
        10'b1010100011: data <= 22'h000238; 
        10'b1010100100: data <= 22'h000afe; 
        10'b1010100101: data <= 22'h001569; 
        10'b1010100110: data <= 22'h00161c; 
        10'b1010100111: data <= 22'h3ff8df; 
        10'b1010101000: data <= 22'h3fdfeb; 
        10'b1010101001: data <= 22'h3fdfc3; 
        10'b1010101010: data <= 22'h3fc753; 
        10'b1010101011: data <= 22'h3fc9bc; 
        10'b1010101100: data <= 22'h3fcf51; 
        10'b1010101101: data <= 22'h3fd64c; 
        10'b1010101110: data <= 22'h3fd67b; 
        10'b1010101111: data <= 22'h3fd663; 
        10'b1010110000: data <= 22'h3ff3f6; 
        10'b1010110001: data <= 22'h00050a; 
        10'b1010110010: data <= 22'h00092f; 
        10'b1010110011: data <= 22'h000d4f; 
        10'b1010110100: data <= 22'h000b27; 
        10'b1010110101: data <= 22'h0002b1; 
        10'b1010110110: data <= 22'h0005c9; 
        10'b1010110111: data <= 22'h000f72; 
        10'b1010111000: data <= 22'h0004ae; 
        10'b1010111001: data <= 22'h00079c; 
        10'b1010111010: data <= 22'h000ea7; 
        10'b1010111011: data <= 22'h0004d6; 
        10'b1010111100: data <= 22'h0012f4; 
        10'b1010111101: data <= 22'h000609; 
        10'b1010111110: data <= 22'h00073b; 
        10'b1010111111: data <= 22'h000a3b; 
        10'b1011000000: data <= 22'h000ea2; 
        10'b1011000001: data <= 22'h000d59; 
        10'b1011000010: data <= 22'h000034; 
        10'b1011000011: data <= 22'h3ff7b9; 
        10'b1011000100: data <= 22'h3ffcb9; 
        10'b1011000101: data <= 22'h3ff860; 
        10'b1011000110: data <= 22'h3fe051; 
        10'b1011000111: data <= 22'h3fd96d; 
        10'b1011001000: data <= 22'h3fe37c; 
        10'b1011001001: data <= 22'h3fd802; 
        10'b1011001010: data <= 22'h3fe78e; 
        10'b1011001011: data <= 22'h3fe10d; 
        10'b1011001100: data <= 22'h3fee2e; 
        10'b1011001101: data <= 22'h3ffcca; 
        10'b1011001110: data <= 22'h000629; 
        10'b1011001111: data <= 22'h000cc9; 
        10'b1011010000: data <= 22'h000138; 
        10'b1011010001: data <= 22'h000b9e; 
        10'b1011010010: data <= 22'h0006e7; 
        10'b1011010011: data <= 22'h001094; 
        10'b1011010100: data <= 22'h00042c; 
        10'b1011010101: data <= 22'h0004f1; 
        10'b1011010110: data <= 22'h000716; 
        10'b1011010111: data <= 22'h00061d; 
        10'b1011011000: data <= 22'h0006f9; 
        10'b1011011001: data <= 22'h000d6d; 
        10'b1011011010: data <= 22'h000bf2; 
        10'b1011011011: data <= 22'h0003a6; 
        10'b1011011100: data <= 22'h000ced; 
        10'b1011011101: data <= 22'h001130; 
        10'b1011011110: data <= 22'h000ba7; 
        10'b1011011111: data <= 22'h000abe; 
        10'b1011100000: data <= 22'h000f59; 
        10'b1011100001: data <= 22'h000cff; 
        10'b1011100010: data <= 22'h0001cf; 
        10'b1011100011: data <= 22'h000a92; 
        10'b1011100100: data <= 22'h0009a0; 
        10'b1011100101: data <= 22'h000592; 
        10'b1011100110: data <= 22'h3fffac; 
        10'b1011100111: data <= 22'h000501; 
        10'b1011101000: data <= 22'h000b43; 
        10'b1011101001: data <= 22'h00116f; 
        10'b1011101010: data <= 22'h000cdb; 
        10'b1011101011: data <= 22'h00020d; 
        10'b1011101100: data <= 22'h000bf4; 
        10'b1011101101: data <= 22'h000b39; 
        10'b1011101110: data <= 22'h000ab3; 
        10'b1011101111: data <= 22'h00051a; 
        10'b1011110000: data <= 22'h00047f; 
        10'b1011110001: data <= 22'h000cf7; 
        10'b1011110010: data <= 22'h0011ba; 
        10'b1011110011: data <= 22'h000e64; 
        10'b1011110100: data <= 22'h000e76; 
        10'b1011110101: data <= 22'h00124d; 
        10'b1011110110: data <= 22'h0002e4; 
        10'b1011110111: data <= 22'h000a1f; 
        10'b1011111000: data <= 22'h001334; 
        10'b1011111001: data <= 22'h000f43; 
        10'b1011111010: data <= 22'h00114c; 
        10'b1011111011: data <= 22'h000ff6; 
        10'b1011111100: data <= 22'h00114e; 
        10'b1011111101: data <= 22'h00082d; 
        10'b1011111110: data <= 22'h000f2a; 
        10'b1011111111: data <= 22'h000fc0; 
        10'b1100000000: data <= 22'h000194; 
        10'b1100000001: data <= 22'h00034a; 
        10'b1100000010: data <= 22'h0012d6; 
        10'b1100000011: data <= 22'h000c4a; 
        10'b1100000100: data <= 22'h000b52; 
        10'b1100000101: data <= 22'h0001a4; 
        10'b1100000110: data <= 22'h000836; 
        10'b1100000111: data <= 22'h00039e; 
        10'b1100001000: data <= 22'h00035e; 
        10'b1100001001: data <= 22'h000628; 
        10'b1100001010: data <= 22'h000b1a; 
        10'b1100001011: data <= 22'h000ffd; 
        10'b1100001100: data <= 22'h0011bd; 
        10'b1100001101: data <= 22'h00114f; 
        10'b1100001110: data <= 22'h00110e; 
        10'b1100001111: data <= 22'h0005b1; 
      endcase 
    end 
  end 
endgenerate 
assign dout = data; 
endmodule
