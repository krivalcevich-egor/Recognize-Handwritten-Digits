`timescale 1ns / 1ps 
 
////////////////////////////////////////////////////////////////////////////////// 
// WEIGHT MEMORY (ROM) 
////////////////////////////////////////////////////////////////////////////////// 
module ROM_weights_6 #( 
    parameter int WGHT_INT = 6, // integer part 
    parameter int WGHT_FRC = 16 // fractional part 
)( 
    input logic clk, // clock 
    input logic [9:0] address,
    output [WGHT_INT + WGHT_FRC-1:0] dout 
); 

(* rom_style = "block" *) reg [WGHT_INT + WGHT_FRC-1:0] data;
generate 
  if (WGHT_FRC == 1) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 7'h00; 
        10'b0000000001: data <= 7'h00; 
        10'b0000000010: data <= 7'h00; 
        10'b0000000011: data <= 7'h00; 
        10'b0000000100: data <= 7'h00; 
        10'b0000000101: data <= 7'h00; 
        10'b0000000110: data <= 7'h00; 
        10'b0000000111: data <= 7'h00; 
        10'b0000001000: data <= 7'h00; 
        10'b0000001001: data <= 7'h00; 
        10'b0000001010: data <= 7'h00; 
        10'b0000001011: data <= 7'h00; 
        10'b0000001100: data <= 7'h00; 
        10'b0000001101: data <= 7'h00; 
        10'b0000001110: data <= 7'h00; 
        10'b0000001111: data <= 7'h00; 
        10'b0000010000: data <= 7'h00; 
        10'b0000010001: data <= 7'h00; 
        10'b0000010010: data <= 7'h00; 
        10'b0000010011: data <= 7'h00; 
        10'b0000010100: data <= 7'h00; 
        10'b0000010101: data <= 7'h00; 
        10'b0000010110: data <= 7'h00; 
        10'b0000010111: data <= 7'h00; 
        10'b0000011000: data <= 7'h00; 
        10'b0000011001: data <= 7'h00; 
        10'b0000011010: data <= 7'h00; 
        10'b0000011011: data <= 7'h00; 
        10'b0000011100: data <= 7'h00; 
        10'b0000011101: data <= 7'h00; 
        10'b0000011110: data <= 7'h00; 
        10'b0000011111: data <= 7'h00; 
        10'b0000100000: data <= 7'h00; 
        10'b0000100001: data <= 7'h00; 
        10'b0000100010: data <= 7'h00; 
        10'b0000100011: data <= 7'h00; 
        10'b0000100100: data <= 7'h00; 
        10'b0000100101: data <= 7'h00; 
        10'b0000100110: data <= 7'h00; 
        10'b0000100111: data <= 7'h00; 
        10'b0000101000: data <= 7'h00; 
        10'b0000101001: data <= 7'h00; 
        10'b0000101010: data <= 7'h00; 
        10'b0000101011: data <= 7'h00; 
        10'b0000101100: data <= 7'h00; 
        10'b0000101101: data <= 7'h00; 
        10'b0000101110: data <= 7'h00; 
        10'b0000101111: data <= 7'h00; 
        10'b0000110000: data <= 7'h00; 
        10'b0000110001: data <= 7'h00; 
        10'b0000110010: data <= 7'h00; 
        10'b0000110011: data <= 7'h00; 
        10'b0000110100: data <= 7'h00; 
        10'b0000110101: data <= 7'h00; 
        10'b0000110110: data <= 7'h00; 
        10'b0000110111: data <= 7'h00; 
        10'b0000111000: data <= 7'h00; 
        10'b0000111001: data <= 7'h00; 
        10'b0000111010: data <= 7'h00; 
        10'b0000111011: data <= 7'h00; 
        10'b0000111100: data <= 7'h00; 
        10'b0000111101: data <= 7'h00; 
        10'b0000111110: data <= 7'h00; 
        10'b0000111111: data <= 7'h00; 
        10'b0001000000: data <= 7'h00; 
        10'b0001000001: data <= 7'h00; 
        10'b0001000010: data <= 7'h00; 
        10'b0001000011: data <= 7'h00; 
        10'b0001000100: data <= 7'h00; 
        10'b0001000101: data <= 7'h00; 
        10'b0001000110: data <= 7'h00; 
        10'b0001000111: data <= 7'h00; 
        10'b0001001000: data <= 7'h00; 
        10'b0001001001: data <= 7'h00; 
        10'b0001001010: data <= 7'h00; 
        10'b0001001011: data <= 7'h00; 
        10'b0001001100: data <= 7'h00; 
        10'b0001001101: data <= 7'h00; 
        10'b0001001110: data <= 7'h00; 
        10'b0001001111: data <= 7'h00; 
        10'b0001010000: data <= 7'h00; 
        10'b0001010001: data <= 7'h00; 
        10'b0001010010: data <= 7'h00; 
        10'b0001010011: data <= 7'h00; 
        10'b0001010100: data <= 7'h00; 
        10'b0001010101: data <= 7'h00; 
        10'b0001010110: data <= 7'h00; 
        10'b0001010111: data <= 7'h00; 
        10'b0001011000: data <= 7'h00; 
        10'b0001011001: data <= 7'h00; 
        10'b0001011010: data <= 7'h00; 
        10'b0001011011: data <= 7'h00; 
        10'b0001011100: data <= 7'h00; 
        10'b0001011101: data <= 7'h00; 
        10'b0001011110: data <= 7'h00; 
        10'b0001011111: data <= 7'h00; 
        10'b0001100000: data <= 7'h00; 
        10'b0001100001: data <= 7'h00; 
        10'b0001100010: data <= 7'h00; 
        10'b0001100011: data <= 7'h00; 
        10'b0001100100: data <= 7'h00; 
        10'b0001100101: data <= 7'h00; 
        10'b0001100110: data <= 7'h00; 
        10'b0001100111: data <= 7'h00; 
        10'b0001101000: data <= 7'h00; 
        10'b0001101001: data <= 7'h00; 
        10'b0001101010: data <= 7'h00; 
        10'b0001101011: data <= 7'h00; 
        10'b0001101100: data <= 7'h00; 
        10'b0001101101: data <= 7'h00; 
        10'b0001101110: data <= 7'h00; 
        10'b0001101111: data <= 7'h00; 
        10'b0001110000: data <= 7'h00; 
        10'b0001110001: data <= 7'h00; 
        10'b0001110010: data <= 7'h00; 
        10'b0001110011: data <= 7'h00; 
        10'b0001110100: data <= 7'h00; 
        10'b0001110101: data <= 7'h00; 
        10'b0001110110: data <= 7'h00; 
        10'b0001110111: data <= 7'h00; 
        10'b0001111000: data <= 7'h00; 
        10'b0001111001: data <= 7'h00; 
        10'b0001111010: data <= 7'h00; 
        10'b0001111011: data <= 7'h00; 
        10'b0001111100: data <= 7'h00; 
        10'b0001111101: data <= 7'h00; 
        10'b0001111110: data <= 7'h00; 
        10'b0001111111: data <= 7'h00; 
        10'b0010000000: data <= 7'h00; 
        10'b0010000001: data <= 7'h00; 
        10'b0010000010: data <= 7'h00; 
        10'b0010000011: data <= 7'h00; 
        10'b0010000100: data <= 7'h00; 
        10'b0010000101: data <= 7'h01; 
        10'b0010000110: data <= 7'h00; 
        10'b0010000111: data <= 7'h00; 
        10'b0010001000: data <= 7'h00; 
        10'b0010001001: data <= 7'h00; 
        10'b0010001010: data <= 7'h00; 
        10'b0010001011: data <= 7'h00; 
        10'b0010001100: data <= 7'h00; 
        10'b0010001101: data <= 7'h00; 
        10'b0010001110: data <= 7'h00; 
        10'b0010001111: data <= 7'h00; 
        10'b0010010000: data <= 7'h00; 
        10'b0010010001: data <= 7'h00; 
        10'b0010010010: data <= 7'h00; 
        10'b0010010011: data <= 7'h00; 
        10'b0010010100: data <= 7'h00; 
        10'b0010010101: data <= 7'h00; 
        10'b0010010110: data <= 7'h00; 
        10'b0010010111: data <= 7'h00; 
        10'b0010011000: data <= 7'h00; 
        10'b0010011001: data <= 7'h00; 
        10'b0010011010: data <= 7'h00; 
        10'b0010011011: data <= 7'h00; 
        10'b0010011100: data <= 7'h00; 
        10'b0010011101: data <= 7'h00; 
        10'b0010011110: data <= 7'h00; 
        10'b0010011111: data <= 7'h00; 
        10'b0010100000: data <= 7'h00; 
        10'b0010100001: data <= 7'h00; 
        10'b0010100010: data <= 7'h00; 
        10'b0010100011: data <= 7'h00; 
        10'b0010100100: data <= 7'h00; 
        10'b0010100101: data <= 7'h00; 
        10'b0010100110: data <= 7'h00; 
        10'b0010100111: data <= 7'h00; 
        10'b0010101000: data <= 7'h00; 
        10'b0010101001: data <= 7'h00; 
        10'b0010101010: data <= 7'h00; 
        10'b0010101011: data <= 7'h00; 
        10'b0010101100: data <= 7'h00; 
        10'b0010101101: data <= 7'h00; 
        10'b0010101110: data <= 7'h00; 
        10'b0010101111: data <= 7'h00; 
        10'b0010110000: data <= 7'h00; 
        10'b0010110001: data <= 7'h00; 
        10'b0010110010: data <= 7'h00; 
        10'b0010110011: data <= 7'h00; 
        10'b0010110100: data <= 7'h00; 
        10'b0010110101: data <= 7'h00; 
        10'b0010110110: data <= 7'h00; 
        10'b0010110111: data <= 7'h00; 
        10'b0010111000: data <= 7'h00; 
        10'b0010111001: data <= 7'h00; 
        10'b0010111010: data <= 7'h00; 
        10'b0010111011: data <= 7'h00; 
        10'b0010111100: data <= 7'h00; 
        10'b0010111101: data <= 7'h00; 
        10'b0010111110: data <= 7'h00; 
        10'b0010111111: data <= 7'h00; 
        10'b0011000000: data <= 7'h00; 
        10'b0011000001: data <= 7'h00; 
        10'b0011000010: data <= 7'h00; 
        10'b0011000011: data <= 7'h00; 
        10'b0011000100: data <= 7'h00; 
        10'b0011000101: data <= 7'h00; 
        10'b0011000110: data <= 7'h00; 
        10'b0011000111: data <= 7'h00; 
        10'b0011001000: data <= 7'h00; 
        10'b0011001001: data <= 7'h00; 
        10'b0011001010: data <= 7'h00; 
        10'b0011001011: data <= 7'h00; 
        10'b0011001100: data <= 7'h00; 
        10'b0011001101: data <= 7'h00; 
        10'b0011001110: data <= 7'h00; 
        10'b0011001111: data <= 7'h00; 
        10'b0011010000: data <= 7'h00; 
        10'b0011010001: data <= 7'h7f; 
        10'b0011010010: data <= 7'h00; 
        10'b0011010011: data <= 7'h00; 
        10'b0011010100: data <= 7'h00; 
        10'b0011010101: data <= 7'h00; 
        10'b0011010110: data <= 7'h00; 
        10'b0011010111: data <= 7'h7f; 
        10'b0011011000: data <= 7'h7f; 
        10'b0011011001: data <= 7'h7f; 
        10'b0011011010: data <= 7'h7f; 
        10'b0011011011: data <= 7'h00; 
        10'b0011011100: data <= 7'h00; 
        10'b0011011101: data <= 7'h00; 
        10'b0011011110: data <= 7'h00; 
        10'b0011011111: data <= 7'h00; 
        10'b0011100000: data <= 7'h00; 
        10'b0011100001: data <= 7'h00; 
        10'b0011100010: data <= 7'h00; 
        10'b0011100011: data <= 7'h00; 
        10'b0011100100: data <= 7'h00; 
        10'b0011100101: data <= 7'h00; 
        10'b0011100110: data <= 7'h00; 
        10'b0011100111: data <= 7'h00; 
        10'b0011101000: data <= 7'h00; 
        10'b0011101001: data <= 7'h00; 
        10'b0011101010: data <= 7'h00; 
        10'b0011101011: data <= 7'h00; 
        10'b0011101100: data <= 7'h00; 
        10'b0011101101: data <= 7'h00; 
        10'b0011101110: data <= 7'h00; 
        10'b0011101111: data <= 7'h00; 
        10'b0011110000: data <= 7'h7f; 
        10'b0011110001: data <= 7'h7f; 
        10'b0011110010: data <= 7'h7f; 
        10'b0011110011: data <= 7'h7f; 
        10'b0011110100: data <= 7'h7f; 
        10'b0011110101: data <= 7'h7f; 
        10'b0011110110: data <= 7'h7f; 
        10'b0011110111: data <= 7'h00; 
        10'b0011111000: data <= 7'h00; 
        10'b0011111001: data <= 7'h00; 
        10'b0011111010: data <= 7'h00; 
        10'b0011111011: data <= 7'h00; 
        10'b0011111100: data <= 7'h00; 
        10'b0011111101: data <= 7'h00; 
        10'b0011111110: data <= 7'h00; 
        10'b0011111111: data <= 7'h00; 
        10'b0100000000: data <= 7'h00; 
        10'b0100000001: data <= 7'h00; 
        10'b0100000010: data <= 7'h00; 
        10'b0100000011: data <= 7'h00; 
        10'b0100000100: data <= 7'h00; 
        10'b0100000101: data <= 7'h00; 
        10'b0100000110: data <= 7'h00; 
        10'b0100000111: data <= 7'h00; 
        10'b0100001000: data <= 7'h00; 
        10'b0100001001: data <= 7'h00; 
        10'b0100001010: data <= 7'h00; 
        10'b0100001011: data <= 7'h7f; 
        10'b0100001100: data <= 7'h7f; 
        10'b0100001101: data <= 7'h7f; 
        10'b0100001110: data <= 7'h7f; 
        10'b0100001111: data <= 7'h7f; 
        10'b0100010000: data <= 7'h7f; 
        10'b0100010001: data <= 7'h7f; 
        10'b0100010010: data <= 7'h7f; 
        10'b0100010011: data <= 7'h00; 
        10'b0100010100: data <= 7'h00; 
        10'b0100010101: data <= 7'h00; 
        10'b0100010110: data <= 7'h00; 
        10'b0100010111: data <= 7'h00; 
        10'b0100011000: data <= 7'h00; 
        10'b0100011001: data <= 7'h00; 
        10'b0100011010: data <= 7'h00; 
        10'b0100011011: data <= 7'h00; 
        10'b0100011100: data <= 7'h00; 
        10'b0100011101: data <= 7'h00; 
        10'b0100011110: data <= 7'h00; 
        10'b0100011111: data <= 7'h00; 
        10'b0100100000: data <= 7'h00; 
        10'b0100100001: data <= 7'h00; 
        10'b0100100010: data <= 7'h00; 
        10'b0100100011: data <= 7'h00; 
        10'b0100100100: data <= 7'h00; 
        10'b0100100101: data <= 7'h00; 
        10'b0100100110: data <= 7'h00; 
        10'b0100100111: data <= 7'h7f; 
        10'b0100101000: data <= 7'h7f; 
        10'b0100101001: data <= 7'h7f; 
        10'b0100101010: data <= 7'h7f; 
        10'b0100101011: data <= 7'h7f; 
        10'b0100101100: data <= 7'h00; 
        10'b0100101101: data <= 7'h00; 
        10'b0100101110: data <= 7'h00; 
        10'b0100101111: data <= 7'h00; 
        10'b0100110000: data <= 7'h00; 
        10'b0100110001: data <= 7'h00; 
        10'b0100110010: data <= 7'h00; 
        10'b0100110011: data <= 7'h00; 
        10'b0100110100: data <= 7'h00; 
        10'b0100110101: data <= 7'h00; 
        10'b0100110110: data <= 7'h00; 
        10'b0100110111: data <= 7'h00; 
        10'b0100111000: data <= 7'h00; 
        10'b0100111001: data <= 7'h00; 
        10'b0100111010: data <= 7'h00; 
        10'b0100111011: data <= 7'h00; 
        10'b0100111100: data <= 7'h00; 
        10'b0100111101: data <= 7'h00; 
        10'b0100111110: data <= 7'h00; 
        10'b0100111111: data <= 7'h00; 
        10'b0101000000: data <= 7'h00; 
        10'b0101000001: data <= 7'h00; 
        10'b0101000010: data <= 7'h00; 
        10'b0101000011: data <= 7'h00; 
        10'b0101000100: data <= 7'h00; 
        10'b0101000101: data <= 7'h00; 
        10'b0101000110: data <= 7'h00; 
        10'b0101000111: data <= 7'h00; 
        10'b0101001000: data <= 7'h00; 
        10'b0101001001: data <= 7'h00; 
        10'b0101001010: data <= 7'h00; 
        10'b0101001011: data <= 7'h00; 
        10'b0101001100: data <= 7'h00; 
        10'b0101001101: data <= 7'h00; 
        10'b0101001110: data <= 7'h00; 
        10'b0101001111: data <= 7'h00; 
        10'b0101010000: data <= 7'h00; 
        10'b0101010001: data <= 7'h00; 
        10'b0101010010: data <= 7'h00; 
        10'b0101010011: data <= 7'h00; 
        10'b0101010100: data <= 7'h00; 
        10'b0101010101: data <= 7'h00; 
        10'b0101010110: data <= 7'h00; 
        10'b0101010111: data <= 7'h00; 
        10'b0101011000: data <= 7'h00; 
        10'b0101011001: data <= 7'h00; 
        10'b0101011010: data <= 7'h00; 
        10'b0101011011: data <= 7'h00; 
        10'b0101011100: data <= 7'h00; 
        10'b0101011101: data <= 7'h00; 
        10'b0101011110: data <= 7'h00; 
        10'b0101011111: data <= 7'h00; 
        10'b0101100000: data <= 7'h00; 
        10'b0101100001: data <= 7'h00; 
        10'b0101100010: data <= 7'h00; 
        10'b0101100011: data <= 7'h00; 
        10'b0101100100: data <= 7'h00; 
        10'b0101100101: data <= 7'h00; 
        10'b0101100110: data <= 7'h00; 
        10'b0101100111: data <= 7'h01; 
        10'b0101101000: data <= 7'h00; 
        10'b0101101001: data <= 7'h00; 
        10'b0101101010: data <= 7'h00; 
        10'b0101101011: data <= 7'h00; 
        10'b0101101100: data <= 7'h00; 
        10'b0101101101: data <= 7'h00; 
        10'b0101101110: data <= 7'h00; 
        10'b0101101111: data <= 7'h00; 
        10'b0101110000: data <= 7'h00; 
        10'b0101110001: data <= 7'h00; 
        10'b0101110010: data <= 7'h00; 
        10'b0101110011: data <= 7'h00; 
        10'b0101110100: data <= 7'h00; 
        10'b0101110101: data <= 7'h00; 
        10'b0101110110: data <= 7'h00; 
        10'b0101110111: data <= 7'h00; 
        10'b0101111000: data <= 7'h00; 
        10'b0101111001: data <= 7'h00; 
        10'b0101111010: data <= 7'h00; 
        10'b0101111011: data <= 7'h00; 
        10'b0101111100: data <= 7'h00; 
        10'b0101111101: data <= 7'h00; 
        10'b0101111110: data <= 7'h00; 
        10'b0101111111: data <= 7'h00; 
        10'b0110000000: data <= 7'h00; 
        10'b0110000001: data <= 7'h00; 
        10'b0110000010: data <= 7'h01; 
        10'b0110000011: data <= 7'h01; 
        10'b0110000100: data <= 7'h00; 
        10'b0110000101: data <= 7'h00; 
        10'b0110000110: data <= 7'h00; 
        10'b0110000111: data <= 7'h00; 
        10'b0110001000: data <= 7'h00; 
        10'b0110001001: data <= 7'h00; 
        10'b0110001010: data <= 7'h00; 
        10'b0110001011: data <= 7'h00; 
        10'b0110001100: data <= 7'h00; 
        10'b0110001101: data <= 7'h00; 
        10'b0110001110: data <= 7'h00; 
        10'b0110001111: data <= 7'h00; 
        10'b0110010000: data <= 7'h00; 
        10'b0110010001: data <= 7'h00; 
        10'b0110010010: data <= 7'h00; 
        10'b0110010011: data <= 7'h00; 
        10'b0110010100: data <= 7'h00; 
        10'b0110010101: data <= 7'h00; 
        10'b0110010110: data <= 7'h00; 
        10'b0110010111: data <= 7'h00; 
        10'b0110011000: data <= 7'h00; 
        10'b0110011001: data <= 7'h00; 
        10'b0110011010: data <= 7'h00; 
        10'b0110011011: data <= 7'h00; 
        10'b0110011100: data <= 7'h00; 
        10'b0110011101: data <= 7'h00; 
        10'b0110011110: data <= 7'h01; 
        10'b0110011111: data <= 7'h01; 
        10'b0110100000: data <= 7'h00; 
        10'b0110100001: data <= 7'h00; 
        10'b0110100010: data <= 7'h00; 
        10'b0110100011: data <= 7'h00; 
        10'b0110100100: data <= 7'h00; 
        10'b0110100101: data <= 7'h00; 
        10'b0110100110: data <= 7'h00; 
        10'b0110100111: data <= 7'h00; 
        10'b0110101000: data <= 7'h00; 
        10'b0110101001: data <= 7'h00; 
        10'b0110101010: data <= 7'h00; 
        10'b0110101011: data <= 7'h00; 
        10'b0110101100: data <= 7'h00; 
        10'b0110101101: data <= 7'h00; 
        10'b0110101110: data <= 7'h00; 
        10'b0110101111: data <= 7'h01; 
        10'b0110110000: data <= 7'h00; 
        10'b0110110001: data <= 7'h00; 
        10'b0110110010: data <= 7'h00; 
        10'b0110110011: data <= 7'h00; 
        10'b0110110100: data <= 7'h00; 
        10'b0110110101: data <= 7'h00; 
        10'b0110110110: data <= 7'h00; 
        10'b0110110111: data <= 7'h00; 
        10'b0110111000: data <= 7'h00; 
        10'b0110111001: data <= 7'h00; 
        10'b0110111010: data <= 7'h00; 
        10'b0110111011: data <= 7'h00; 
        10'b0110111100: data <= 7'h00; 
        10'b0110111101: data <= 7'h00; 
        10'b0110111110: data <= 7'h00; 
        10'b0110111111: data <= 7'h00; 
        10'b0111000000: data <= 7'h00; 
        10'b0111000001: data <= 7'h00; 
        10'b0111000010: data <= 7'h00; 
        10'b0111000011: data <= 7'h00; 
        10'b0111000100: data <= 7'h00; 
        10'b0111000101: data <= 7'h00; 
        10'b0111000110: data <= 7'h00; 
        10'b0111000111: data <= 7'h00; 
        10'b0111001000: data <= 7'h00; 
        10'b0111001001: data <= 7'h00; 
        10'b0111001010: data <= 7'h01; 
        10'b0111001011: data <= 7'h01; 
        10'b0111001100: data <= 7'h00; 
        10'b0111001101: data <= 7'h00; 
        10'b0111001110: data <= 7'h00; 
        10'b0111001111: data <= 7'h00; 
        10'b0111010000: data <= 7'h00; 
        10'b0111010001: data <= 7'h00; 
        10'b0111010010: data <= 7'h00; 
        10'b0111010011: data <= 7'h00; 
        10'b0111010100: data <= 7'h00; 
        10'b0111010101: data <= 7'h00; 
        10'b0111010110: data <= 7'h00; 
        10'b0111010111: data <= 7'h00; 
        10'b0111011000: data <= 7'h00; 
        10'b0111011001: data <= 7'h00; 
        10'b0111011010: data <= 7'h00; 
        10'b0111011011: data <= 7'h00; 
        10'b0111011100: data <= 7'h00; 
        10'b0111011101: data <= 7'h00; 
        10'b0111011110: data <= 7'h00; 
        10'b0111011111: data <= 7'h00; 
        10'b0111100000: data <= 7'h00; 
        10'b0111100001: data <= 7'h00; 
        10'b0111100010: data <= 7'h00; 
        10'b0111100011: data <= 7'h00; 
        10'b0111100100: data <= 7'h00; 
        10'b0111100101: data <= 7'h00; 
        10'b0111100110: data <= 7'h01; 
        10'b0111100111: data <= 7'h01; 
        10'b0111101000: data <= 7'h00; 
        10'b0111101001: data <= 7'h00; 
        10'b0111101010: data <= 7'h00; 
        10'b0111101011: data <= 7'h00; 
        10'b0111101100: data <= 7'h00; 
        10'b0111101101: data <= 7'h00; 
        10'b0111101110: data <= 7'h00; 
        10'b0111101111: data <= 7'h00; 
        10'b0111110000: data <= 7'h00; 
        10'b0111110001: data <= 7'h00; 
        10'b0111110010: data <= 7'h00; 
        10'b0111110011: data <= 7'h00; 
        10'b0111110100: data <= 7'h00; 
        10'b0111110101: data <= 7'h00; 
        10'b0111110110: data <= 7'h00; 
        10'b0111110111: data <= 7'h00; 
        10'b0111111000: data <= 7'h00; 
        10'b0111111001: data <= 7'h00; 
        10'b0111111010: data <= 7'h00; 
        10'b0111111011: data <= 7'h00; 
        10'b0111111100: data <= 7'h00; 
        10'b0111111101: data <= 7'h00; 
        10'b0111111110: data <= 7'h00; 
        10'b0111111111: data <= 7'h00; 
        10'b1000000000: data <= 7'h00; 
        10'b1000000001: data <= 7'h00; 
        10'b1000000010: data <= 7'h01; 
        10'b1000000011: data <= 7'h01; 
        10'b1000000100: data <= 7'h01; 
        10'b1000000101: data <= 7'h00; 
        10'b1000000110: data <= 7'h00; 
        10'b1000000111: data <= 7'h00; 
        10'b1000001000: data <= 7'h00; 
        10'b1000001001: data <= 7'h00; 
        10'b1000001010: data <= 7'h00; 
        10'b1000001011: data <= 7'h00; 
        10'b1000001100: data <= 7'h00; 
        10'b1000001101: data <= 7'h00; 
        10'b1000001110: data <= 7'h00; 
        10'b1000001111: data <= 7'h00; 
        10'b1000010000: data <= 7'h00; 
        10'b1000010001: data <= 7'h00; 
        10'b1000010010: data <= 7'h00; 
        10'b1000010011: data <= 7'h00; 
        10'b1000010100: data <= 7'h00; 
        10'b1000010101: data <= 7'h00; 
        10'b1000010110: data <= 7'h00; 
        10'b1000010111: data <= 7'h00; 
        10'b1000011000: data <= 7'h00; 
        10'b1000011001: data <= 7'h00; 
        10'b1000011010: data <= 7'h00; 
        10'b1000011011: data <= 7'h00; 
        10'b1000011100: data <= 7'h00; 
        10'b1000011101: data <= 7'h00; 
        10'b1000011110: data <= 7'h00; 
        10'b1000011111: data <= 7'h01; 
        10'b1000100000: data <= 7'h01; 
        10'b1000100001: data <= 7'h00; 
        10'b1000100010: data <= 7'h00; 
        10'b1000100011: data <= 7'h00; 
        10'b1000100100: data <= 7'h00; 
        10'b1000100101: data <= 7'h00; 
        10'b1000100110: data <= 7'h00; 
        10'b1000100111: data <= 7'h00; 
        10'b1000101000: data <= 7'h00; 
        10'b1000101001: data <= 7'h00; 
        10'b1000101010: data <= 7'h00; 
        10'b1000101011: data <= 7'h00; 
        10'b1000101100: data <= 7'h00; 
        10'b1000101101: data <= 7'h00; 
        10'b1000101110: data <= 7'h00; 
        10'b1000101111: data <= 7'h00; 
        10'b1000110000: data <= 7'h00; 
        10'b1000110001: data <= 7'h00; 
        10'b1000110010: data <= 7'h00; 
        10'b1000110011: data <= 7'h00; 
        10'b1000110100: data <= 7'h00; 
        10'b1000110101: data <= 7'h00; 
        10'b1000110110: data <= 7'h00; 
        10'b1000110111: data <= 7'h00; 
        10'b1000111000: data <= 7'h00; 
        10'b1000111001: data <= 7'h00; 
        10'b1000111010: data <= 7'h00; 
        10'b1000111011: data <= 7'h00; 
        10'b1000111100: data <= 7'h01; 
        10'b1000111101: data <= 7'h01; 
        10'b1000111110: data <= 7'h01; 
        10'b1000111111: data <= 7'h01; 
        10'b1001000000: data <= 7'h00; 
        10'b1001000001: data <= 7'h00; 
        10'b1001000010: data <= 7'h00; 
        10'b1001000011: data <= 7'h00; 
        10'b1001000100: data <= 7'h00; 
        10'b1001000101: data <= 7'h00; 
        10'b1001000110: data <= 7'h00; 
        10'b1001000111: data <= 7'h00; 
        10'b1001001000: data <= 7'h00; 
        10'b1001001001: data <= 7'h00; 
        10'b1001001010: data <= 7'h00; 
        10'b1001001011: data <= 7'h00; 
        10'b1001001100: data <= 7'h00; 
        10'b1001001101: data <= 7'h00; 
        10'b1001001110: data <= 7'h00; 
        10'b1001001111: data <= 7'h00; 
        10'b1001010000: data <= 7'h00; 
        10'b1001010001: data <= 7'h00; 
        10'b1001010010: data <= 7'h00; 
        10'b1001010011: data <= 7'h00; 
        10'b1001010100: data <= 7'h00; 
        10'b1001010101: data <= 7'h00; 
        10'b1001010110: data <= 7'h00; 
        10'b1001010111: data <= 7'h00; 
        10'b1001011000: data <= 7'h01; 
        10'b1001011001: data <= 7'h01; 
        10'b1001011010: data <= 7'h01; 
        10'b1001011011: data <= 7'h00; 
        10'b1001011100: data <= 7'h00; 
        10'b1001011101: data <= 7'h00; 
        10'b1001011110: data <= 7'h00; 
        10'b1001011111: data <= 7'h00; 
        10'b1001100000: data <= 7'h00; 
        10'b1001100001: data <= 7'h00; 
        10'b1001100010: data <= 7'h00; 
        10'b1001100011: data <= 7'h00; 
        10'b1001100100: data <= 7'h00; 
        10'b1001100101: data <= 7'h00; 
        10'b1001100110: data <= 7'h00; 
        10'b1001100111: data <= 7'h00; 
        10'b1001101000: data <= 7'h00; 
        10'b1001101001: data <= 7'h00; 
        10'b1001101010: data <= 7'h00; 
        10'b1001101011: data <= 7'h00; 
        10'b1001101100: data <= 7'h00; 
        10'b1001101101: data <= 7'h00; 
        10'b1001101110: data <= 7'h00; 
        10'b1001101111: data <= 7'h00; 
        10'b1001110000: data <= 7'h00; 
        10'b1001110001: data <= 7'h00; 
        10'b1001110010: data <= 7'h00; 
        10'b1001110011: data <= 7'h00; 
        10'b1001110100: data <= 7'h00; 
        10'b1001110101: data <= 7'h00; 
        10'b1001110110: data <= 7'h00; 
        10'b1001110111: data <= 7'h00; 
        10'b1001111000: data <= 7'h00; 
        10'b1001111001: data <= 7'h00; 
        10'b1001111010: data <= 7'h00; 
        10'b1001111011: data <= 7'h00; 
        10'b1001111100: data <= 7'h00; 
        10'b1001111101: data <= 7'h00; 
        10'b1001111110: data <= 7'h00; 
        10'b1001111111: data <= 7'h00; 
        10'b1010000000: data <= 7'h00; 
        10'b1010000001: data <= 7'h00; 
        10'b1010000010: data <= 7'h00; 
        10'b1010000011: data <= 7'h00; 
        10'b1010000100: data <= 7'h00; 
        10'b1010000101: data <= 7'h00; 
        10'b1010000110: data <= 7'h00; 
        10'b1010000111: data <= 7'h00; 
        10'b1010001000: data <= 7'h00; 
        10'b1010001001: data <= 7'h00; 
        10'b1010001010: data <= 7'h00; 
        10'b1010001011: data <= 7'h00; 
        10'b1010001100: data <= 7'h00; 
        10'b1010001101: data <= 7'h7f; 
        10'b1010001110: data <= 7'h7f; 
        10'b1010001111: data <= 7'h7f; 
        10'b1010010000: data <= 7'h00; 
        10'b1010010001: data <= 7'h00; 
        10'b1010010010: data <= 7'h00; 
        10'b1010010011: data <= 7'h00; 
        10'b1010010100: data <= 7'h00; 
        10'b1010010101: data <= 7'h7f; 
        10'b1010010110: data <= 7'h00; 
        10'b1010010111: data <= 7'h00; 
        10'b1010011000: data <= 7'h00; 
        10'b1010011001: data <= 7'h00; 
        10'b1010011010: data <= 7'h00; 
        10'b1010011011: data <= 7'h00; 
        10'b1010011100: data <= 7'h00; 
        10'b1010011101: data <= 7'h00; 
        10'b1010011110: data <= 7'h00; 
        10'b1010011111: data <= 7'h00; 
        10'b1010100000: data <= 7'h00; 
        10'b1010100001: data <= 7'h00; 
        10'b1010100010: data <= 7'h00; 
        10'b1010100011: data <= 7'h00; 
        10'b1010100100: data <= 7'h00; 
        10'b1010100101: data <= 7'h00; 
        10'b1010100110: data <= 7'h00; 
        10'b1010100111: data <= 7'h00; 
        10'b1010101000: data <= 7'h00; 
        10'b1010101001: data <= 7'h00; 
        10'b1010101010: data <= 7'h00; 
        10'b1010101011: data <= 7'h00; 
        10'b1010101100: data <= 7'h00; 
        10'b1010101101: data <= 7'h00; 
        10'b1010101110: data <= 7'h00; 
        10'b1010101111: data <= 7'h00; 
        10'b1010110000: data <= 7'h00; 
        10'b1010110001: data <= 7'h00; 
        10'b1010110010: data <= 7'h00; 
        10'b1010110011: data <= 7'h00; 
        10'b1010110100: data <= 7'h00; 
        10'b1010110101: data <= 7'h00; 
        10'b1010110110: data <= 7'h00; 
        10'b1010110111: data <= 7'h00; 
        10'b1010111000: data <= 7'h00; 
        10'b1010111001: data <= 7'h00; 
        10'b1010111010: data <= 7'h00; 
        10'b1010111011: data <= 7'h00; 
        10'b1010111100: data <= 7'h00; 
        10'b1010111101: data <= 7'h00; 
        10'b1010111110: data <= 7'h00; 
        10'b1010111111: data <= 7'h00; 
        10'b1011000000: data <= 7'h00; 
        10'b1011000001: data <= 7'h00; 
        10'b1011000010: data <= 7'h00; 
        10'b1011000011: data <= 7'h00; 
        10'b1011000100: data <= 7'h00; 
        10'b1011000101: data <= 7'h00; 
        10'b1011000110: data <= 7'h00; 
        10'b1011000111: data <= 7'h00; 
        10'b1011001000: data <= 7'h00; 
        10'b1011001001: data <= 7'h00; 
        10'b1011001010: data <= 7'h00; 
        10'b1011001011: data <= 7'h00; 
        10'b1011001100: data <= 7'h00; 
        10'b1011001101: data <= 7'h00; 
        10'b1011001110: data <= 7'h00; 
        10'b1011001111: data <= 7'h00; 
        10'b1011010000: data <= 7'h00; 
        10'b1011010001: data <= 7'h00; 
        10'b1011010010: data <= 7'h00; 
        10'b1011010011: data <= 7'h00; 
        10'b1011010100: data <= 7'h00; 
        10'b1011010101: data <= 7'h00; 
        10'b1011010110: data <= 7'h00; 
        10'b1011010111: data <= 7'h00; 
        10'b1011011000: data <= 7'h00; 
        10'b1011011001: data <= 7'h00; 
        10'b1011011010: data <= 7'h00; 
        10'b1011011011: data <= 7'h00; 
        10'b1011011100: data <= 7'h00; 
        10'b1011011101: data <= 7'h00; 
        10'b1011011110: data <= 7'h00; 
        10'b1011011111: data <= 7'h00; 
        10'b1011100000: data <= 7'h00; 
        10'b1011100001: data <= 7'h00; 
        10'b1011100010: data <= 7'h00; 
        10'b1011100011: data <= 7'h00; 
        10'b1011100100: data <= 7'h00; 
        10'b1011100101: data <= 7'h00; 
        10'b1011100110: data <= 7'h00; 
        10'b1011100111: data <= 7'h00; 
        10'b1011101000: data <= 7'h00; 
        10'b1011101001: data <= 7'h00; 
        10'b1011101010: data <= 7'h00; 
        10'b1011101011: data <= 7'h00; 
        10'b1011101100: data <= 7'h00; 
        10'b1011101101: data <= 7'h00; 
        10'b1011101110: data <= 7'h00; 
        10'b1011101111: data <= 7'h00; 
        10'b1011110000: data <= 7'h00; 
        10'b1011110001: data <= 7'h00; 
        10'b1011110010: data <= 7'h00; 
        10'b1011110011: data <= 7'h00; 
        10'b1011110100: data <= 7'h00; 
        10'b1011110101: data <= 7'h00; 
        10'b1011110110: data <= 7'h00; 
        10'b1011110111: data <= 7'h00; 
        10'b1011111000: data <= 7'h00; 
        10'b1011111001: data <= 7'h00; 
        10'b1011111010: data <= 7'h00; 
        10'b1011111011: data <= 7'h00; 
        10'b1011111100: data <= 7'h00; 
        10'b1011111101: data <= 7'h00; 
        10'b1011111110: data <= 7'h00; 
        10'b1011111111: data <= 7'h00; 
        10'b1100000000: data <= 7'h00; 
        10'b1100000001: data <= 7'h00; 
        10'b1100000010: data <= 7'h00; 
        10'b1100000011: data <= 7'h00; 
        10'b1100000100: data <= 7'h00; 
        10'b1100000101: data <= 7'h00; 
        10'b1100000110: data <= 7'h00; 
        10'b1100000111: data <= 7'h00; 
        10'b1100001000: data <= 7'h00; 
        10'b1100001001: data <= 7'h00; 
        10'b1100001010: data <= 7'h00; 
        10'b1100001011: data <= 7'h00; 
        10'b1100001100: data <= 7'h00; 
        10'b1100001101: data <= 7'h00; 
        10'b1100001110: data <= 7'h00; 
        10'b1100001111: data <= 7'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 2) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 8'h00; 
        10'b0000000001: data <= 8'h00; 
        10'b0000000010: data <= 8'h00; 
        10'b0000000011: data <= 8'h00; 
        10'b0000000100: data <= 8'h00; 
        10'b0000000101: data <= 8'h00; 
        10'b0000000110: data <= 8'h00; 
        10'b0000000111: data <= 8'h00; 
        10'b0000001000: data <= 8'h00; 
        10'b0000001001: data <= 8'h00; 
        10'b0000001010: data <= 8'h00; 
        10'b0000001011: data <= 8'h00; 
        10'b0000001100: data <= 8'h00; 
        10'b0000001101: data <= 8'h00; 
        10'b0000001110: data <= 8'h00; 
        10'b0000001111: data <= 8'h00; 
        10'b0000010000: data <= 8'h00; 
        10'b0000010001: data <= 8'h00; 
        10'b0000010010: data <= 8'h00; 
        10'b0000010011: data <= 8'h00; 
        10'b0000010100: data <= 8'h00; 
        10'b0000010101: data <= 8'h00; 
        10'b0000010110: data <= 8'h00; 
        10'b0000010111: data <= 8'h00; 
        10'b0000011000: data <= 8'h00; 
        10'b0000011001: data <= 8'h00; 
        10'b0000011010: data <= 8'h00; 
        10'b0000011011: data <= 8'h00; 
        10'b0000011100: data <= 8'h00; 
        10'b0000011101: data <= 8'h00; 
        10'b0000011110: data <= 8'h00; 
        10'b0000011111: data <= 8'h00; 
        10'b0000100000: data <= 8'h00; 
        10'b0000100001: data <= 8'h00; 
        10'b0000100010: data <= 8'h00; 
        10'b0000100011: data <= 8'h00; 
        10'b0000100100: data <= 8'h00; 
        10'b0000100101: data <= 8'h00; 
        10'b0000100110: data <= 8'h00; 
        10'b0000100111: data <= 8'h00; 
        10'b0000101000: data <= 8'h00; 
        10'b0000101001: data <= 8'h00; 
        10'b0000101010: data <= 8'h00; 
        10'b0000101011: data <= 8'h00; 
        10'b0000101100: data <= 8'h00; 
        10'b0000101101: data <= 8'h00; 
        10'b0000101110: data <= 8'h00; 
        10'b0000101111: data <= 8'h00; 
        10'b0000110000: data <= 8'h00; 
        10'b0000110001: data <= 8'h00; 
        10'b0000110010: data <= 8'h00; 
        10'b0000110011: data <= 8'h00; 
        10'b0000110100: data <= 8'h00; 
        10'b0000110101: data <= 8'h00; 
        10'b0000110110: data <= 8'h00; 
        10'b0000110111: data <= 8'h00; 
        10'b0000111000: data <= 8'h00; 
        10'b0000111001: data <= 8'h00; 
        10'b0000111010: data <= 8'h00; 
        10'b0000111011: data <= 8'h00; 
        10'b0000111100: data <= 8'h00; 
        10'b0000111101: data <= 8'h00; 
        10'b0000111110: data <= 8'h00; 
        10'b0000111111: data <= 8'h00; 
        10'b0001000000: data <= 8'h00; 
        10'b0001000001: data <= 8'h00; 
        10'b0001000010: data <= 8'h00; 
        10'b0001000011: data <= 8'h00; 
        10'b0001000100: data <= 8'h00; 
        10'b0001000101: data <= 8'h00; 
        10'b0001000110: data <= 8'h00; 
        10'b0001000111: data <= 8'h00; 
        10'b0001001000: data <= 8'h00; 
        10'b0001001001: data <= 8'h00; 
        10'b0001001010: data <= 8'h00; 
        10'b0001001011: data <= 8'h00; 
        10'b0001001100: data <= 8'h00; 
        10'b0001001101: data <= 8'h00; 
        10'b0001001110: data <= 8'h00; 
        10'b0001001111: data <= 8'h00; 
        10'b0001010000: data <= 8'h00; 
        10'b0001010001: data <= 8'h00; 
        10'b0001010010: data <= 8'h00; 
        10'b0001010011: data <= 8'h00; 
        10'b0001010100: data <= 8'h00; 
        10'b0001010101: data <= 8'h00; 
        10'b0001010110: data <= 8'h00; 
        10'b0001010111: data <= 8'h00; 
        10'b0001011000: data <= 8'h00; 
        10'b0001011001: data <= 8'h00; 
        10'b0001011010: data <= 8'h00; 
        10'b0001011011: data <= 8'h00; 
        10'b0001011100: data <= 8'h00; 
        10'b0001011101: data <= 8'h00; 
        10'b0001011110: data <= 8'h00; 
        10'b0001011111: data <= 8'h00; 
        10'b0001100000: data <= 8'h00; 
        10'b0001100001: data <= 8'h00; 
        10'b0001100010: data <= 8'h01; 
        10'b0001100011: data <= 8'h01; 
        10'b0001100100: data <= 8'h00; 
        10'b0001100101: data <= 8'h00; 
        10'b0001100110: data <= 8'h01; 
        10'b0001100111: data <= 8'h01; 
        10'b0001101000: data <= 8'h01; 
        10'b0001101001: data <= 8'h01; 
        10'b0001101010: data <= 8'h01; 
        10'b0001101011: data <= 8'h00; 
        10'b0001101100: data <= 8'h00; 
        10'b0001101101: data <= 8'h00; 
        10'b0001101110: data <= 8'h00; 
        10'b0001101111: data <= 8'h00; 
        10'b0001110000: data <= 8'h00; 
        10'b0001110001: data <= 8'h00; 
        10'b0001110010: data <= 8'h00; 
        10'b0001110011: data <= 8'h00; 
        10'b0001110100: data <= 8'h00; 
        10'b0001110101: data <= 8'h00; 
        10'b0001110110: data <= 8'h00; 
        10'b0001110111: data <= 8'h00; 
        10'b0001111000: data <= 8'h00; 
        10'b0001111001: data <= 8'h00; 
        10'b0001111010: data <= 8'h00; 
        10'b0001111011: data <= 8'h00; 
        10'b0001111100: data <= 8'h00; 
        10'b0001111101: data <= 8'h00; 
        10'b0001111110: data <= 8'h00; 
        10'b0001111111: data <= 8'h00; 
        10'b0010000000: data <= 8'h00; 
        10'b0010000001: data <= 8'h00; 
        10'b0010000010: data <= 8'h01; 
        10'b0010000011: data <= 8'h01; 
        10'b0010000100: data <= 8'h01; 
        10'b0010000101: data <= 8'h01; 
        10'b0010000110: data <= 8'h01; 
        10'b0010000111: data <= 8'h01; 
        10'b0010001000: data <= 8'h00; 
        10'b0010001001: data <= 8'h00; 
        10'b0010001010: data <= 8'h00; 
        10'b0010001011: data <= 8'h00; 
        10'b0010001100: data <= 8'h00; 
        10'b0010001101: data <= 8'h00; 
        10'b0010001110: data <= 8'h00; 
        10'b0010001111: data <= 8'h00; 
        10'b0010010000: data <= 8'h00; 
        10'b0010010001: data <= 8'h00; 
        10'b0010010010: data <= 8'h00; 
        10'b0010010011: data <= 8'h00; 
        10'b0010010100: data <= 8'h00; 
        10'b0010010101: data <= 8'h00; 
        10'b0010010110: data <= 8'h00; 
        10'b0010010111: data <= 8'hff; 
        10'b0010011000: data <= 8'h00; 
        10'b0010011001: data <= 8'h00; 
        10'b0010011010: data <= 8'h00; 
        10'b0010011011: data <= 8'h00; 
        10'b0010011100: data <= 8'h00; 
        10'b0010011101: data <= 8'h00; 
        10'b0010011110: data <= 8'h00; 
        10'b0010011111: data <= 8'h01; 
        10'b0010100000: data <= 8'h01; 
        10'b0010100001: data <= 8'h01; 
        10'b0010100010: data <= 8'h00; 
        10'b0010100011: data <= 8'h00; 
        10'b0010100100: data <= 8'h00; 
        10'b0010100101: data <= 8'h00; 
        10'b0010100110: data <= 8'h00; 
        10'b0010100111: data <= 8'h00; 
        10'b0010101000: data <= 8'h00; 
        10'b0010101001: data <= 8'h00; 
        10'b0010101010: data <= 8'h00; 
        10'b0010101011: data <= 8'h00; 
        10'b0010101100: data <= 8'h00; 
        10'b0010101101: data <= 8'h00; 
        10'b0010101110: data <= 8'h00; 
        10'b0010101111: data <= 8'h00; 
        10'b0010110000: data <= 8'h00; 
        10'b0010110001: data <= 8'h00; 
        10'b0010110010: data <= 8'hff; 
        10'b0010110011: data <= 8'hff; 
        10'b0010110100: data <= 8'h00; 
        10'b0010110101: data <= 8'hff; 
        10'b0010110110: data <= 8'h00; 
        10'b0010110111: data <= 8'h00; 
        10'b0010111000: data <= 8'h00; 
        10'b0010111001: data <= 8'h00; 
        10'b0010111010: data <= 8'h00; 
        10'b0010111011: data <= 8'h00; 
        10'b0010111100: data <= 8'h00; 
        10'b0010111101: data <= 8'h00; 
        10'b0010111110: data <= 8'hff; 
        10'b0010111111: data <= 8'h00; 
        10'b0011000000: data <= 8'h00; 
        10'b0011000001: data <= 8'h00; 
        10'b0011000010: data <= 8'h00; 
        10'b0011000011: data <= 8'h00; 
        10'b0011000100: data <= 8'h00; 
        10'b0011000101: data <= 8'h00; 
        10'b0011000110: data <= 8'h00; 
        10'b0011000111: data <= 8'h00; 
        10'b0011001000: data <= 8'h00; 
        10'b0011001001: data <= 8'h00; 
        10'b0011001010: data <= 8'h00; 
        10'b0011001011: data <= 8'h00; 
        10'b0011001100: data <= 8'h00; 
        10'b0011001101: data <= 8'h00; 
        10'b0011001110: data <= 8'hff; 
        10'b0011001111: data <= 8'hff; 
        10'b0011010000: data <= 8'hff; 
        10'b0011010001: data <= 8'hff; 
        10'b0011010010: data <= 8'hff; 
        10'b0011010011: data <= 8'hff; 
        10'b0011010100: data <= 8'hff; 
        10'b0011010101: data <= 8'hff; 
        10'b0011010110: data <= 8'hff; 
        10'b0011010111: data <= 8'hff; 
        10'b0011011000: data <= 8'hff; 
        10'b0011011001: data <= 8'hff; 
        10'b0011011010: data <= 8'hff; 
        10'b0011011011: data <= 8'hff; 
        10'b0011011100: data <= 8'h00; 
        10'b0011011101: data <= 8'h00; 
        10'b0011011110: data <= 8'h00; 
        10'b0011011111: data <= 8'h00; 
        10'b0011100000: data <= 8'h00; 
        10'b0011100001: data <= 8'h00; 
        10'b0011100010: data <= 8'h00; 
        10'b0011100011: data <= 8'h00; 
        10'b0011100100: data <= 8'h00; 
        10'b0011100101: data <= 8'h00; 
        10'b0011100110: data <= 8'h00; 
        10'b0011100111: data <= 8'h00; 
        10'b0011101000: data <= 8'h00; 
        10'b0011101001: data <= 8'hff; 
        10'b0011101010: data <= 8'hff; 
        10'b0011101011: data <= 8'hff; 
        10'b0011101100: data <= 8'hff; 
        10'b0011101101: data <= 8'hff; 
        10'b0011101110: data <= 8'hff; 
        10'b0011101111: data <= 8'hff; 
        10'b0011110000: data <= 8'hff; 
        10'b0011110001: data <= 8'hff; 
        10'b0011110010: data <= 8'hfe; 
        10'b0011110011: data <= 8'hfe; 
        10'b0011110100: data <= 8'hfe; 
        10'b0011110101: data <= 8'hfe; 
        10'b0011110110: data <= 8'hff; 
        10'b0011110111: data <= 8'hff; 
        10'b0011111000: data <= 8'hff; 
        10'b0011111001: data <= 8'h00; 
        10'b0011111010: data <= 8'h00; 
        10'b0011111011: data <= 8'h00; 
        10'b0011111100: data <= 8'h00; 
        10'b0011111101: data <= 8'h00; 
        10'b0011111110: data <= 8'h00; 
        10'b0011111111: data <= 8'h00; 
        10'b0100000000: data <= 8'h00; 
        10'b0100000001: data <= 8'h00; 
        10'b0100000010: data <= 8'h00; 
        10'b0100000011: data <= 8'h00; 
        10'b0100000100: data <= 8'h00; 
        10'b0100000101: data <= 8'h00; 
        10'b0100000110: data <= 8'hff; 
        10'b0100000111: data <= 8'h00; 
        10'b0100001000: data <= 8'h00; 
        10'b0100001001: data <= 8'hff; 
        10'b0100001010: data <= 8'h00; 
        10'b0100001011: data <= 8'hff; 
        10'b0100001100: data <= 8'hff; 
        10'b0100001101: data <= 8'hfe; 
        10'b0100001110: data <= 8'hfe; 
        10'b0100001111: data <= 8'hfe; 
        10'b0100010000: data <= 8'hff; 
        10'b0100010001: data <= 8'hff; 
        10'b0100010010: data <= 8'hff; 
        10'b0100010011: data <= 8'hff; 
        10'b0100010100: data <= 8'hff; 
        10'b0100010101: data <= 8'h00; 
        10'b0100010110: data <= 8'h00; 
        10'b0100010111: data <= 8'h00; 
        10'b0100011000: data <= 8'h00; 
        10'b0100011001: data <= 8'h00; 
        10'b0100011010: data <= 8'h00; 
        10'b0100011011: data <= 8'h00; 
        10'b0100011100: data <= 8'h00; 
        10'b0100011101: data <= 8'h00; 
        10'b0100011110: data <= 8'h00; 
        10'b0100011111: data <= 8'h00; 
        10'b0100100000: data <= 8'h01; 
        10'b0100100001: data <= 8'h00; 
        10'b0100100010: data <= 8'h00; 
        10'b0100100011: data <= 8'h00; 
        10'b0100100100: data <= 8'h00; 
        10'b0100100101: data <= 8'h00; 
        10'b0100100110: data <= 8'hff; 
        10'b0100100111: data <= 8'hff; 
        10'b0100101000: data <= 8'hff; 
        10'b0100101001: data <= 8'hff; 
        10'b0100101010: data <= 8'hff; 
        10'b0100101011: data <= 8'hff; 
        10'b0100101100: data <= 8'hff; 
        10'b0100101101: data <= 8'hff; 
        10'b0100101110: data <= 8'hff; 
        10'b0100101111: data <= 8'h00; 
        10'b0100110000: data <= 8'h00; 
        10'b0100110001: data <= 8'h00; 
        10'b0100110010: data <= 8'h00; 
        10'b0100110011: data <= 8'h00; 
        10'b0100110100: data <= 8'h00; 
        10'b0100110101: data <= 8'h00; 
        10'b0100110110: data <= 8'h00; 
        10'b0100110111: data <= 8'h00; 
        10'b0100111000: data <= 8'h00; 
        10'b0100111001: data <= 8'h00; 
        10'b0100111010: data <= 8'h00; 
        10'b0100111011: data <= 8'h00; 
        10'b0100111100: data <= 8'h00; 
        10'b0100111101: data <= 8'h00; 
        10'b0100111110: data <= 8'h00; 
        10'b0100111111: data <= 8'h00; 
        10'b0101000000: data <= 8'h00; 
        10'b0101000001: data <= 8'h00; 
        10'b0101000010: data <= 8'h00; 
        10'b0101000011: data <= 8'hff; 
        10'b0101000100: data <= 8'hff; 
        10'b0101000101: data <= 8'hff; 
        10'b0101000110: data <= 8'hff; 
        10'b0101000111: data <= 8'hff; 
        10'b0101001000: data <= 8'h00; 
        10'b0101001001: data <= 8'h00; 
        10'b0101001010: data <= 8'h00; 
        10'b0101001011: data <= 8'h01; 
        10'b0101001100: data <= 8'h00; 
        10'b0101001101: data <= 8'h00; 
        10'b0101001110: data <= 8'h00; 
        10'b0101001111: data <= 8'h00; 
        10'b0101010000: data <= 8'h00; 
        10'b0101010001: data <= 8'h00; 
        10'b0101010010: data <= 8'h00; 
        10'b0101010011: data <= 8'h00; 
        10'b0101010100: data <= 8'h00; 
        10'b0101010101: data <= 8'h00; 
        10'b0101010110: data <= 8'h00; 
        10'b0101010111: data <= 8'h00; 
        10'b0101011000: data <= 8'h00; 
        10'b0101011001: data <= 8'h00; 
        10'b0101011010: data <= 8'h00; 
        10'b0101011011: data <= 8'h01; 
        10'b0101011100: data <= 8'h01; 
        10'b0101011101: data <= 8'h00; 
        10'b0101011110: data <= 8'h00; 
        10'b0101011111: data <= 8'hff; 
        10'b0101100000: data <= 8'h00; 
        10'b0101100001: data <= 8'h00; 
        10'b0101100010: data <= 8'hff; 
        10'b0101100011: data <= 8'hff; 
        10'b0101100100: data <= 8'h00; 
        10'b0101100101: data <= 8'h00; 
        10'b0101100110: data <= 8'h01; 
        10'b0101100111: data <= 8'h01; 
        10'b0101101000: data <= 8'h01; 
        10'b0101101001: data <= 8'h00; 
        10'b0101101010: data <= 8'h00; 
        10'b0101101011: data <= 8'h00; 
        10'b0101101100: data <= 8'h00; 
        10'b0101101101: data <= 8'h00; 
        10'b0101101110: data <= 8'h00; 
        10'b0101101111: data <= 8'h00; 
        10'b0101110000: data <= 8'h00; 
        10'b0101110001: data <= 8'h00; 
        10'b0101110010: data <= 8'h01; 
        10'b0101110011: data <= 8'h00; 
        10'b0101110100: data <= 8'h00; 
        10'b0101110101: data <= 8'h00; 
        10'b0101110110: data <= 8'h01; 
        10'b0101110111: data <= 8'h00; 
        10'b0101111000: data <= 8'h00; 
        10'b0101111001: data <= 8'h00; 
        10'b0101111010: data <= 8'h00; 
        10'b0101111011: data <= 8'h00; 
        10'b0101111100: data <= 8'h00; 
        10'b0101111101: data <= 8'h00; 
        10'b0101111110: data <= 8'hff; 
        10'b0101111111: data <= 8'h00; 
        10'b0110000000: data <= 8'h00; 
        10'b0110000001: data <= 8'h00; 
        10'b0110000010: data <= 8'h01; 
        10'b0110000011: data <= 8'h02; 
        10'b0110000100: data <= 8'h01; 
        10'b0110000101: data <= 8'h00; 
        10'b0110000110: data <= 8'h00; 
        10'b0110000111: data <= 8'h00; 
        10'b0110001000: data <= 8'h00; 
        10'b0110001001: data <= 8'h00; 
        10'b0110001010: data <= 8'h00; 
        10'b0110001011: data <= 8'h00; 
        10'b0110001100: data <= 8'h00; 
        10'b0110001101: data <= 8'h00; 
        10'b0110001110: data <= 8'h01; 
        10'b0110001111: data <= 8'h00; 
        10'b0110010000: data <= 8'h01; 
        10'b0110010001: data <= 8'h01; 
        10'b0110010010: data <= 8'h01; 
        10'b0110010011: data <= 8'h01; 
        10'b0110010100: data <= 8'h00; 
        10'b0110010101: data <= 8'h00; 
        10'b0110010110: data <= 8'h00; 
        10'b0110010111: data <= 8'h00; 
        10'b0110011000: data <= 8'h00; 
        10'b0110011001: data <= 8'h00; 
        10'b0110011010: data <= 8'h00; 
        10'b0110011011: data <= 8'h00; 
        10'b0110011100: data <= 8'h00; 
        10'b0110011101: data <= 8'h00; 
        10'b0110011110: data <= 8'h01; 
        10'b0110011111: data <= 8'h01; 
        10'b0110100000: data <= 8'h01; 
        10'b0110100001: data <= 8'h00; 
        10'b0110100010: data <= 8'h00; 
        10'b0110100011: data <= 8'h00; 
        10'b0110100100: data <= 8'h00; 
        10'b0110100101: data <= 8'h00; 
        10'b0110100110: data <= 8'h00; 
        10'b0110100111: data <= 8'h00; 
        10'b0110101000: data <= 8'h00; 
        10'b0110101001: data <= 8'h00; 
        10'b0110101010: data <= 8'h01; 
        10'b0110101011: data <= 8'h01; 
        10'b0110101100: data <= 8'h00; 
        10'b0110101101: data <= 8'h01; 
        10'b0110101110: data <= 8'h01; 
        10'b0110101111: data <= 8'h01; 
        10'b0110110000: data <= 8'h00; 
        10'b0110110001: data <= 8'h00; 
        10'b0110110010: data <= 8'h00; 
        10'b0110110011: data <= 8'h00; 
        10'b0110110100: data <= 8'h00; 
        10'b0110110101: data <= 8'h00; 
        10'b0110110110: data <= 8'h00; 
        10'b0110110111: data <= 8'h00; 
        10'b0110111000: data <= 8'h01; 
        10'b0110111001: data <= 8'h01; 
        10'b0110111010: data <= 8'h01; 
        10'b0110111011: data <= 8'h01; 
        10'b0110111100: data <= 8'h00; 
        10'b0110111101: data <= 8'h00; 
        10'b0110111110: data <= 8'h00; 
        10'b0110111111: data <= 8'h00; 
        10'b0111000000: data <= 8'h00; 
        10'b0111000001: data <= 8'h00; 
        10'b0111000010: data <= 8'h00; 
        10'b0111000011: data <= 8'h00; 
        10'b0111000100: data <= 8'hff; 
        10'b0111000101: data <= 8'h00; 
        10'b0111000110: data <= 8'h01; 
        10'b0111000111: data <= 8'h01; 
        10'b0111001000: data <= 8'h01; 
        10'b0111001001: data <= 8'h01; 
        10'b0111001010: data <= 8'h01; 
        10'b0111001011: data <= 8'h01; 
        10'b0111001100: data <= 8'h00; 
        10'b0111001101: data <= 8'h00; 
        10'b0111001110: data <= 8'h01; 
        10'b0111001111: data <= 8'h00; 
        10'b0111010000: data <= 8'h00; 
        10'b0111010001: data <= 8'h00; 
        10'b0111010010: data <= 8'h00; 
        10'b0111010011: data <= 8'h00; 
        10'b0111010100: data <= 8'h00; 
        10'b0111010101: data <= 8'h00; 
        10'b0111010110: data <= 8'h00; 
        10'b0111010111: data <= 8'h00; 
        10'b0111011000: data <= 8'h00; 
        10'b0111011001: data <= 8'h00; 
        10'b0111011010: data <= 8'h00; 
        10'b0111011011: data <= 8'h00; 
        10'b0111011100: data <= 8'h00; 
        10'b0111011101: data <= 8'h00; 
        10'b0111011110: data <= 8'h00; 
        10'b0111011111: data <= 8'h00; 
        10'b0111100000: data <= 8'hff; 
        10'b0111100001: data <= 8'h00; 
        10'b0111100010: data <= 8'h00; 
        10'b0111100011: data <= 8'h01; 
        10'b0111100100: data <= 8'h01; 
        10'b0111100101: data <= 8'h01; 
        10'b0111100110: data <= 8'h02; 
        10'b0111100111: data <= 8'h02; 
        10'b0111101000: data <= 8'h01; 
        10'b0111101001: data <= 8'h00; 
        10'b0111101010: data <= 8'h00; 
        10'b0111101011: data <= 8'h00; 
        10'b0111101100: data <= 8'h00; 
        10'b0111101101: data <= 8'h00; 
        10'b0111101110: data <= 8'h01; 
        10'b0111101111: data <= 8'h00; 
        10'b0111110000: data <= 8'h00; 
        10'b0111110001: data <= 8'h00; 
        10'b0111110010: data <= 8'h00; 
        10'b0111110011: data <= 8'h00; 
        10'b0111110100: data <= 8'h00; 
        10'b0111110101: data <= 8'h00; 
        10'b0111110110: data <= 8'h00; 
        10'b0111110111: data <= 8'h00; 
        10'b0111111000: data <= 8'h00; 
        10'b0111111001: data <= 8'h00; 
        10'b0111111010: data <= 8'h00; 
        10'b0111111011: data <= 8'h00; 
        10'b0111111100: data <= 8'hff; 
        10'b0111111101: data <= 8'hff; 
        10'b0111111110: data <= 8'h00; 
        10'b0111111111: data <= 8'h00; 
        10'b1000000000: data <= 8'h01; 
        10'b1000000001: data <= 8'h01; 
        10'b1000000010: data <= 8'h01; 
        10'b1000000011: data <= 8'h01; 
        10'b1000000100: data <= 8'h02; 
        10'b1000000101: data <= 8'h01; 
        10'b1000000110: data <= 8'h00; 
        10'b1000000111: data <= 8'h00; 
        10'b1000001000: data <= 8'h01; 
        10'b1000001001: data <= 8'h00; 
        10'b1000001010: data <= 8'h01; 
        10'b1000001011: data <= 8'h00; 
        10'b1000001100: data <= 8'h00; 
        10'b1000001101: data <= 8'h00; 
        10'b1000001110: data <= 8'h00; 
        10'b1000001111: data <= 8'h00; 
        10'b1000010000: data <= 8'h00; 
        10'b1000010001: data <= 8'h00; 
        10'b1000010010: data <= 8'h00; 
        10'b1000010011: data <= 8'h00; 
        10'b1000010100: data <= 8'h00; 
        10'b1000010101: data <= 8'h00; 
        10'b1000010110: data <= 8'h00; 
        10'b1000010111: data <= 8'h00; 
        10'b1000011000: data <= 8'h00; 
        10'b1000011001: data <= 8'hff; 
        10'b1000011010: data <= 8'hff; 
        10'b1000011011: data <= 8'h00; 
        10'b1000011100: data <= 8'h00; 
        10'b1000011101: data <= 8'h01; 
        10'b1000011110: data <= 8'h01; 
        10'b1000011111: data <= 8'h02; 
        10'b1000100000: data <= 8'h02; 
        10'b1000100001: data <= 8'h01; 
        10'b1000100010: data <= 8'h01; 
        10'b1000100011: data <= 8'h01; 
        10'b1000100100: data <= 8'h01; 
        10'b1000100101: data <= 8'h01; 
        10'b1000100110: data <= 8'h01; 
        10'b1000100111: data <= 8'h01; 
        10'b1000101000: data <= 8'h00; 
        10'b1000101001: data <= 8'h00; 
        10'b1000101010: data <= 8'h00; 
        10'b1000101011: data <= 8'h00; 
        10'b1000101100: data <= 8'h00; 
        10'b1000101101: data <= 8'h00; 
        10'b1000101110: data <= 8'h00; 
        10'b1000101111: data <= 8'h00; 
        10'b1000110000: data <= 8'h00; 
        10'b1000110001: data <= 8'h00; 
        10'b1000110010: data <= 8'h00; 
        10'b1000110011: data <= 8'h00; 
        10'b1000110100: data <= 8'hff; 
        10'b1000110101: data <= 8'hff; 
        10'b1000110110: data <= 8'hff; 
        10'b1000110111: data <= 8'h00; 
        10'b1000111000: data <= 8'h00; 
        10'b1000111001: data <= 8'h00; 
        10'b1000111010: data <= 8'h01; 
        10'b1000111011: data <= 8'h01; 
        10'b1000111100: data <= 8'h01; 
        10'b1000111101: data <= 8'h01; 
        10'b1000111110: data <= 8'h02; 
        10'b1000111111: data <= 8'h01; 
        10'b1001000000: data <= 8'h01; 
        10'b1001000001: data <= 8'h00; 
        10'b1001000010: data <= 8'h01; 
        10'b1001000011: data <= 8'h01; 
        10'b1001000100: data <= 8'h00; 
        10'b1001000101: data <= 8'h00; 
        10'b1001000110: data <= 8'h00; 
        10'b1001000111: data <= 8'h00; 
        10'b1001001000: data <= 8'h00; 
        10'b1001001001: data <= 8'h00; 
        10'b1001001010: data <= 8'h00; 
        10'b1001001011: data <= 8'h00; 
        10'b1001001100: data <= 8'h00; 
        10'b1001001101: data <= 8'h00; 
        10'b1001001110: data <= 8'h00; 
        10'b1001001111: data <= 8'h00; 
        10'b1001010000: data <= 8'h00; 
        10'b1001010001: data <= 8'h00; 
        10'b1001010010: data <= 8'hff; 
        10'b1001010011: data <= 8'h00; 
        10'b1001010100: data <= 8'h00; 
        10'b1001010101: data <= 8'h00; 
        10'b1001010110: data <= 8'h01; 
        10'b1001010111: data <= 8'h01; 
        10'b1001011000: data <= 8'h01; 
        10'b1001011001: data <= 8'h01; 
        10'b1001011010: data <= 8'h01; 
        10'b1001011011: data <= 8'h01; 
        10'b1001011100: data <= 8'h01; 
        10'b1001011101: data <= 8'h01; 
        10'b1001011110: data <= 8'h01; 
        10'b1001011111: data <= 8'h00; 
        10'b1001100000: data <= 8'h00; 
        10'b1001100001: data <= 8'h00; 
        10'b1001100010: data <= 8'h00; 
        10'b1001100011: data <= 8'h00; 
        10'b1001100100: data <= 8'h00; 
        10'b1001100101: data <= 8'h00; 
        10'b1001100110: data <= 8'h00; 
        10'b1001100111: data <= 8'h00; 
        10'b1001101000: data <= 8'h00; 
        10'b1001101001: data <= 8'h00; 
        10'b1001101010: data <= 8'h00; 
        10'b1001101011: data <= 8'h00; 
        10'b1001101100: data <= 8'h00; 
        10'b1001101101: data <= 8'h00; 
        10'b1001101110: data <= 8'h00; 
        10'b1001101111: data <= 8'hff; 
        10'b1001110000: data <= 8'h00; 
        10'b1001110001: data <= 8'h00; 
        10'b1001110010: data <= 8'h00; 
        10'b1001110011: data <= 8'h00; 
        10'b1001110100: data <= 8'h00; 
        10'b1001110101: data <= 8'h00; 
        10'b1001110110: data <= 8'h00; 
        10'b1001110111: data <= 8'h00; 
        10'b1001111000: data <= 8'h00; 
        10'b1001111001: data <= 8'h00; 
        10'b1001111010: data <= 8'h00; 
        10'b1001111011: data <= 8'h00; 
        10'b1001111100: data <= 8'h00; 
        10'b1001111101: data <= 8'h00; 
        10'b1001111110: data <= 8'h00; 
        10'b1001111111: data <= 8'h00; 
        10'b1010000000: data <= 8'h00; 
        10'b1010000001: data <= 8'h00; 
        10'b1010000010: data <= 8'h00; 
        10'b1010000011: data <= 8'h00; 
        10'b1010000100: data <= 8'h00; 
        10'b1010000101: data <= 8'h00; 
        10'b1010000110: data <= 8'h00; 
        10'b1010000111: data <= 8'h00; 
        10'b1010001000: data <= 8'h00; 
        10'b1010001001: data <= 8'h00; 
        10'b1010001010: data <= 8'h00; 
        10'b1010001011: data <= 8'hff; 
        10'b1010001100: data <= 8'hff; 
        10'b1010001101: data <= 8'hff; 
        10'b1010001110: data <= 8'hff; 
        10'b1010001111: data <= 8'hff; 
        10'b1010010000: data <= 8'hff; 
        10'b1010010001: data <= 8'hff; 
        10'b1010010010: data <= 8'h00; 
        10'b1010010011: data <= 8'hff; 
        10'b1010010100: data <= 8'hff; 
        10'b1010010101: data <= 8'hff; 
        10'b1010010110: data <= 8'hff; 
        10'b1010010111: data <= 8'h00; 
        10'b1010011000: data <= 8'h00; 
        10'b1010011001: data <= 8'h00; 
        10'b1010011010: data <= 8'h00; 
        10'b1010011011: data <= 8'h00; 
        10'b1010011100: data <= 8'h00; 
        10'b1010011101: data <= 8'h00; 
        10'b1010011110: data <= 8'h00; 
        10'b1010011111: data <= 8'h00; 
        10'b1010100000: data <= 8'h00; 
        10'b1010100001: data <= 8'h00; 
        10'b1010100010: data <= 8'h00; 
        10'b1010100011: data <= 8'h00; 
        10'b1010100100: data <= 8'h00; 
        10'b1010100101: data <= 8'h00; 
        10'b1010100110: data <= 8'h00; 
        10'b1010100111: data <= 8'h00; 
        10'b1010101000: data <= 8'h00; 
        10'b1010101001: data <= 8'h00; 
        10'b1010101010: data <= 8'h00; 
        10'b1010101011: data <= 8'h00; 
        10'b1010101100: data <= 8'hff; 
        10'b1010101101: data <= 8'hff; 
        10'b1010101110: data <= 8'hff; 
        10'b1010101111: data <= 8'hff; 
        10'b1010110000: data <= 8'hff; 
        10'b1010110001: data <= 8'hff; 
        10'b1010110010: data <= 8'h00; 
        10'b1010110011: data <= 8'h00; 
        10'b1010110100: data <= 8'h00; 
        10'b1010110101: data <= 8'h00; 
        10'b1010110110: data <= 8'h00; 
        10'b1010110111: data <= 8'h00; 
        10'b1010111000: data <= 8'h00; 
        10'b1010111001: data <= 8'h00; 
        10'b1010111010: data <= 8'h00; 
        10'b1010111011: data <= 8'h00; 
        10'b1010111100: data <= 8'h00; 
        10'b1010111101: data <= 8'h00; 
        10'b1010111110: data <= 8'h00; 
        10'b1010111111: data <= 8'h00; 
        10'b1011000000: data <= 8'h00; 
        10'b1011000001: data <= 8'h00; 
        10'b1011000010: data <= 8'h00; 
        10'b1011000011: data <= 8'h00; 
        10'b1011000100: data <= 8'h00; 
        10'b1011000101: data <= 8'h00; 
        10'b1011000110: data <= 8'h00; 
        10'b1011000111: data <= 8'h00; 
        10'b1011001000: data <= 8'h00; 
        10'b1011001001: data <= 8'h00; 
        10'b1011001010: data <= 8'h00; 
        10'b1011001011: data <= 8'h00; 
        10'b1011001100: data <= 8'h00; 
        10'b1011001101: data <= 8'h00; 
        10'b1011001110: data <= 8'h00; 
        10'b1011001111: data <= 8'h00; 
        10'b1011010000: data <= 8'h00; 
        10'b1011010001: data <= 8'h00; 
        10'b1011010010: data <= 8'h00; 
        10'b1011010011: data <= 8'h00; 
        10'b1011010100: data <= 8'h00; 
        10'b1011010101: data <= 8'h00; 
        10'b1011010110: data <= 8'h00; 
        10'b1011010111: data <= 8'h00; 
        10'b1011011000: data <= 8'h00; 
        10'b1011011001: data <= 8'h00; 
        10'b1011011010: data <= 8'h00; 
        10'b1011011011: data <= 8'h00; 
        10'b1011011100: data <= 8'h00; 
        10'b1011011101: data <= 8'h00; 
        10'b1011011110: data <= 8'h00; 
        10'b1011011111: data <= 8'h00; 
        10'b1011100000: data <= 8'h00; 
        10'b1011100001: data <= 8'h00; 
        10'b1011100010: data <= 8'h00; 
        10'b1011100011: data <= 8'h00; 
        10'b1011100100: data <= 8'h00; 
        10'b1011100101: data <= 8'h00; 
        10'b1011100110: data <= 8'h00; 
        10'b1011100111: data <= 8'h00; 
        10'b1011101000: data <= 8'h00; 
        10'b1011101001: data <= 8'h00; 
        10'b1011101010: data <= 8'h00; 
        10'b1011101011: data <= 8'h00; 
        10'b1011101100: data <= 8'h00; 
        10'b1011101101: data <= 8'h00; 
        10'b1011101110: data <= 8'h00; 
        10'b1011101111: data <= 8'h00; 
        10'b1011110000: data <= 8'h00; 
        10'b1011110001: data <= 8'h00; 
        10'b1011110010: data <= 8'h00; 
        10'b1011110011: data <= 8'h00; 
        10'b1011110100: data <= 8'h00; 
        10'b1011110101: data <= 8'h00; 
        10'b1011110110: data <= 8'h00; 
        10'b1011110111: data <= 8'h00; 
        10'b1011111000: data <= 8'h00; 
        10'b1011111001: data <= 8'h00; 
        10'b1011111010: data <= 8'h00; 
        10'b1011111011: data <= 8'h00; 
        10'b1011111100: data <= 8'h00; 
        10'b1011111101: data <= 8'h00; 
        10'b1011111110: data <= 8'h00; 
        10'b1011111111: data <= 8'h00; 
        10'b1100000000: data <= 8'h00; 
        10'b1100000001: data <= 8'h00; 
        10'b1100000010: data <= 8'h00; 
        10'b1100000011: data <= 8'h00; 
        10'b1100000100: data <= 8'h00; 
        10'b1100000101: data <= 8'h00; 
        10'b1100000110: data <= 8'h00; 
        10'b1100000111: data <= 8'h00; 
        10'b1100001000: data <= 8'h00; 
        10'b1100001001: data <= 8'h00; 
        10'b1100001010: data <= 8'h00; 
        10'b1100001011: data <= 8'h00; 
        10'b1100001100: data <= 8'h00; 
        10'b1100001101: data <= 8'h00; 
        10'b1100001110: data <= 8'h00; 
        10'b1100001111: data <= 8'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 3) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 9'h000; 
        10'b0000000001: data <= 9'h000; 
        10'b0000000010: data <= 9'h000; 
        10'b0000000011: data <= 9'h000; 
        10'b0000000100: data <= 9'h000; 
        10'b0000000101: data <= 9'h000; 
        10'b0000000110: data <= 9'h000; 
        10'b0000000111: data <= 9'h000; 
        10'b0000001000: data <= 9'h000; 
        10'b0000001001: data <= 9'h000; 
        10'b0000001010: data <= 9'h000; 
        10'b0000001011: data <= 9'h000; 
        10'b0000001100: data <= 9'h000; 
        10'b0000001101: data <= 9'h000; 
        10'b0000001110: data <= 9'h000; 
        10'b0000001111: data <= 9'h000; 
        10'b0000010000: data <= 9'h000; 
        10'b0000010001: data <= 9'h000; 
        10'b0000010010: data <= 9'h000; 
        10'b0000010011: data <= 9'h000; 
        10'b0000010100: data <= 9'h000; 
        10'b0000010101: data <= 9'h000; 
        10'b0000010110: data <= 9'h000; 
        10'b0000010111: data <= 9'h000; 
        10'b0000011000: data <= 9'h000; 
        10'b0000011001: data <= 9'h000; 
        10'b0000011010: data <= 9'h000; 
        10'b0000011011: data <= 9'h000; 
        10'b0000011100: data <= 9'h000; 
        10'b0000011101: data <= 9'h000; 
        10'b0000011110: data <= 9'h000; 
        10'b0000011111: data <= 9'h000; 
        10'b0000100000: data <= 9'h000; 
        10'b0000100001: data <= 9'h000; 
        10'b0000100010: data <= 9'h000; 
        10'b0000100011: data <= 9'h000; 
        10'b0000100100: data <= 9'h000; 
        10'b0000100101: data <= 9'h000; 
        10'b0000100110: data <= 9'h000; 
        10'b0000100111: data <= 9'h000; 
        10'b0000101000: data <= 9'h000; 
        10'b0000101001: data <= 9'h000; 
        10'b0000101010: data <= 9'h000; 
        10'b0000101011: data <= 9'h000; 
        10'b0000101100: data <= 9'h000; 
        10'b0000101101: data <= 9'h000; 
        10'b0000101110: data <= 9'h000; 
        10'b0000101111: data <= 9'h000; 
        10'b0000110000: data <= 9'h000; 
        10'b0000110001: data <= 9'h000; 
        10'b0000110010: data <= 9'h000; 
        10'b0000110011: data <= 9'h000; 
        10'b0000110100: data <= 9'h000; 
        10'b0000110101: data <= 9'h000; 
        10'b0000110110: data <= 9'h000; 
        10'b0000110111: data <= 9'h000; 
        10'b0000111000: data <= 9'h000; 
        10'b0000111001: data <= 9'h000; 
        10'b0000111010: data <= 9'h000; 
        10'b0000111011: data <= 9'h000; 
        10'b0000111100: data <= 9'h000; 
        10'b0000111101: data <= 9'h000; 
        10'b0000111110: data <= 9'h000; 
        10'b0000111111: data <= 9'h000; 
        10'b0001000000: data <= 9'h000; 
        10'b0001000001: data <= 9'h001; 
        10'b0001000010: data <= 9'h001; 
        10'b0001000011: data <= 9'h001; 
        10'b0001000100: data <= 9'h001; 
        10'b0001000101: data <= 9'h001; 
        10'b0001000110: data <= 9'h000; 
        10'b0001000111: data <= 9'h000; 
        10'b0001001000: data <= 9'h001; 
        10'b0001001001: data <= 9'h000; 
        10'b0001001010: data <= 9'h000; 
        10'b0001001011: data <= 9'h000; 
        10'b0001001100: data <= 9'h000; 
        10'b0001001101: data <= 9'h000; 
        10'b0001001110: data <= 9'h000; 
        10'b0001001111: data <= 9'h000; 
        10'b0001010000: data <= 9'h000; 
        10'b0001010001: data <= 9'h000; 
        10'b0001010010: data <= 9'h000; 
        10'b0001010011: data <= 9'h000; 
        10'b0001010100: data <= 9'h000; 
        10'b0001010101: data <= 9'h000; 
        10'b0001010110: data <= 9'h000; 
        10'b0001010111: data <= 9'h000; 
        10'b0001011000: data <= 9'h000; 
        10'b0001011001: data <= 9'h000; 
        10'b0001011010: data <= 9'h000; 
        10'b0001011011: data <= 9'h000; 
        10'b0001011100: data <= 9'h000; 
        10'b0001011101: data <= 9'h001; 
        10'b0001011110: data <= 9'h001; 
        10'b0001011111: data <= 9'h001; 
        10'b0001100000: data <= 9'h001; 
        10'b0001100001: data <= 9'h001; 
        10'b0001100010: data <= 9'h001; 
        10'b0001100011: data <= 9'h001; 
        10'b0001100100: data <= 9'h001; 
        10'b0001100101: data <= 9'h001; 
        10'b0001100110: data <= 9'h001; 
        10'b0001100111: data <= 9'h001; 
        10'b0001101000: data <= 9'h002; 
        10'b0001101001: data <= 9'h001; 
        10'b0001101010: data <= 9'h001; 
        10'b0001101011: data <= 9'h001; 
        10'b0001101100: data <= 9'h001; 
        10'b0001101101: data <= 9'h000; 
        10'b0001101110: data <= 9'h000; 
        10'b0001101111: data <= 9'h000; 
        10'b0001110000: data <= 9'h000; 
        10'b0001110001: data <= 9'h000; 
        10'b0001110010: data <= 9'h000; 
        10'b0001110011: data <= 9'h000; 
        10'b0001110100: data <= 9'h000; 
        10'b0001110101: data <= 9'h000; 
        10'b0001110110: data <= 9'h000; 
        10'b0001110111: data <= 9'h000; 
        10'b0001111000: data <= 9'h000; 
        10'b0001111001: data <= 9'h000; 
        10'b0001111010: data <= 9'h000; 
        10'b0001111011: data <= 9'h000; 
        10'b0001111100: data <= 9'h000; 
        10'b0001111101: data <= 9'h000; 
        10'b0001111110: data <= 9'h000; 
        10'b0001111111: data <= 9'h000; 
        10'b0010000000: data <= 9'h001; 
        10'b0010000001: data <= 9'h001; 
        10'b0010000010: data <= 9'h001; 
        10'b0010000011: data <= 9'h002; 
        10'b0010000100: data <= 9'h002; 
        10'b0010000101: data <= 9'h002; 
        10'b0010000110: data <= 9'h002; 
        10'b0010000111: data <= 9'h001; 
        10'b0010001000: data <= 9'h000; 
        10'b0010001001: data <= 9'h000; 
        10'b0010001010: data <= 9'h000; 
        10'b0010001011: data <= 9'h000; 
        10'b0010001100: data <= 9'h000; 
        10'b0010001101: data <= 9'h000; 
        10'b0010001110: data <= 9'h000; 
        10'b0010001111: data <= 9'h000; 
        10'b0010010000: data <= 9'h000; 
        10'b0010010001: data <= 9'h000; 
        10'b0010010010: data <= 9'h000; 
        10'b0010010011: data <= 9'h000; 
        10'b0010010100: data <= 9'h000; 
        10'b0010010101: data <= 9'h000; 
        10'b0010010110: data <= 9'h000; 
        10'b0010010111: data <= 9'h1ff; 
        10'b0010011000: data <= 9'h1ff; 
        10'b0010011001: data <= 9'h000; 
        10'b0010011010: data <= 9'h000; 
        10'b0010011011: data <= 9'h1ff; 
        10'b0010011100: data <= 9'h1ff; 
        10'b0010011101: data <= 9'h000; 
        10'b0010011110: data <= 9'h001; 
        10'b0010011111: data <= 9'h001; 
        10'b0010100000: data <= 9'h001; 
        10'b0010100001: data <= 9'h001; 
        10'b0010100010: data <= 9'h001; 
        10'b0010100011: data <= 9'h001; 
        10'b0010100100: data <= 9'h000; 
        10'b0010100101: data <= 9'h000; 
        10'b0010100110: data <= 9'h000; 
        10'b0010100111: data <= 9'h000; 
        10'b0010101000: data <= 9'h000; 
        10'b0010101001: data <= 9'h000; 
        10'b0010101010: data <= 9'h000; 
        10'b0010101011: data <= 9'h000; 
        10'b0010101100: data <= 9'h000; 
        10'b0010101101: data <= 9'h000; 
        10'b0010101110: data <= 9'h000; 
        10'b0010101111: data <= 9'h000; 
        10'b0010110000: data <= 9'h000; 
        10'b0010110001: data <= 9'h1ff; 
        10'b0010110010: data <= 9'h1ff; 
        10'b0010110011: data <= 9'h1fe; 
        10'b0010110100: data <= 9'h1ff; 
        10'b0010110101: data <= 9'h1fe; 
        10'b0010110110: data <= 9'h1ff; 
        10'b0010110111: data <= 9'h1ff; 
        10'b0010111000: data <= 9'h1ff; 
        10'b0010111001: data <= 9'h1ff; 
        10'b0010111010: data <= 9'h000; 
        10'b0010111011: data <= 9'h1ff; 
        10'b0010111100: data <= 9'h1ff; 
        10'b0010111101: data <= 9'h1ff; 
        10'b0010111110: data <= 9'h1ff; 
        10'b0010111111: data <= 9'h1ff; 
        10'b0011000000: data <= 9'h1ff; 
        10'b0011000001: data <= 9'h1ff; 
        10'b0011000010: data <= 9'h000; 
        10'b0011000011: data <= 9'h000; 
        10'b0011000100: data <= 9'h000; 
        10'b0011000101: data <= 9'h000; 
        10'b0011000110: data <= 9'h000; 
        10'b0011000111: data <= 9'h000; 
        10'b0011001000: data <= 9'h000; 
        10'b0011001001: data <= 9'h000; 
        10'b0011001010: data <= 9'h1ff; 
        10'b0011001011: data <= 9'h000; 
        10'b0011001100: data <= 9'h1ff; 
        10'b0011001101: data <= 9'h1ff; 
        10'b0011001110: data <= 9'h1ff; 
        10'b0011001111: data <= 9'h1ff; 
        10'b0011010000: data <= 9'h1fe; 
        10'b0011010001: data <= 9'h1fe; 
        10'b0011010010: data <= 9'h1ff; 
        10'b0011010011: data <= 9'h1ff; 
        10'b0011010100: data <= 9'h1fe; 
        10'b0011010101: data <= 9'h1fe; 
        10'b0011010110: data <= 9'h1fe; 
        10'b0011010111: data <= 9'h1fd; 
        10'b0011011000: data <= 9'h1fd; 
        10'b0011011001: data <= 9'h1fe; 
        10'b0011011010: data <= 9'h1fe; 
        10'b0011011011: data <= 9'h1fe; 
        10'b0011011100: data <= 9'h1ff; 
        10'b0011011101: data <= 9'h1ff; 
        10'b0011011110: data <= 9'h000; 
        10'b0011011111: data <= 9'h000; 
        10'b0011100000: data <= 9'h000; 
        10'b0011100001: data <= 9'h000; 
        10'b0011100010: data <= 9'h000; 
        10'b0011100011: data <= 9'h000; 
        10'b0011100100: data <= 9'h000; 
        10'b0011100101: data <= 9'h000; 
        10'b0011100110: data <= 9'h1ff; 
        10'b0011100111: data <= 9'h000; 
        10'b0011101000: data <= 9'h000; 
        10'b0011101001: data <= 9'h1ff; 
        10'b0011101010: data <= 9'h1ff; 
        10'b0011101011: data <= 9'h1ff; 
        10'b0011101100: data <= 9'h1fe; 
        10'b0011101101: data <= 9'h1fe; 
        10'b0011101110: data <= 9'h1fe; 
        10'b0011101111: data <= 9'h1fe; 
        10'b0011110000: data <= 9'h1fe; 
        10'b0011110001: data <= 9'h1fd; 
        10'b0011110010: data <= 9'h1fc; 
        10'b0011110011: data <= 9'h1fc; 
        10'b0011110100: data <= 9'h1fd; 
        10'b0011110101: data <= 9'h1fd; 
        10'b0011110110: data <= 9'h1fe; 
        10'b0011110111: data <= 9'h1fe; 
        10'b0011111000: data <= 9'h1ff; 
        10'b0011111001: data <= 9'h1ff; 
        10'b0011111010: data <= 9'h1ff; 
        10'b0011111011: data <= 9'h000; 
        10'b0011111100: data <= 9'h000; 
        10'b0011111101: data <= 9'h000; 
        10'b0011111110: data <= 9'h000; 
        10'b0011111111: data <= 9'h000; 
        10'b0100000000: data <= 9'h000; 
        10'b0100000001: data <= 9'h000; 
        10'b0100000010: data <= 9'h000; 
        10'b0100000011: data <= 9'h000; 
        10'b0100000100: data <= 9'h000; 
        10'b0100000101: data <= 9'h1ff; 
        10'b0100000110: data <= 9'h1ff; 
        10'b0100000111: data <= 9'h1ff; 
        10'b0100001000: data <= 9'h1ff; 
        10'b0100001001: data <= 9'h1ff; 
        10'b0100001010: data <= 9'h1ff; 
        10'b0100001011: data <= 9'h1fe; 
        10'b0100001100: data <= 9'h1fd; 
        10'b0100001101: data <= 9'h1fc; 
        10'b0100001110: data <= 9'h1fc; 
        10'b0100001111: data <= 9'h1fd; 
        10'b0100010000: data <= 9'h1fd; 
        10'b0100010001: data <= 9'h1fe; 
        10'b0100010010: data <= 9'h1fe; 
        10'b0100010011: data <= 9'h1fe; 
        10'b0100010100: data <= 9'h1ff; 
        10'b0100010101: data <= 9'h1ff; 
        10'b0100010110: data <= 9'h000; 
        10'b0100010111: data <= 9'h000; 
        10'b0100011000: data <= 9'h000; 
        10'b0100011001: data <= 9'h000; 
        10'b0100011010: data <= 9'h000; 
        10'b0100011011: data <= 9'h000; 
        10'b0100011100: data <= 9'h000; 
        10'b0100011101: data <= 9'h000; 
        10'b0100011110: data <= 9'h000; 
        10'b0100011111: data <= 9'h000; 
        10'b0100100000: data <= 9'h001; 
        10'b0100100001: data <= 9'h000; 
        10'b0100100010: data <= 9'h000; 
        10'b0100100011: data <= 9'h000; 
        10'b0100100100: data <= 9'h1ff; 
        10'b0100100101: data <= 9'h000; 
        10'b0100100110: data <= 9'h1ff; 
        10'b0100100111: data <= 9'h1fe; 
        10'b0100101000: data <= 9'h1fe; 
        10'b0100101001: data <= 9'h1fd; 
        10'b0100101010: data <= 9'h1fd; 
        10'b0100101011: data <= 9'h1fe; 
        10'b0100101100: data <= 9'h1fe; 
        10'b0100101101: data <= 9'h1ff; 
        10'b0100101110: data <= 9'h1ff; 
        10'b0100101111: data <= 9'h000; 
        10'b0100110000: data <= 9'h1ff; 
        10'b0100110001: data <= 9'h1ff; 
        10'b0100110010: data <= 9'h000; 
        10'b0100110011: data <= 9'h000; 
        10'b0100110100: data <= 9'h000; 
        10'b0100110101: data <= 9'h000; 
        10'b0100110110: data <= 9'h000; 
        10'b0100110111: data <= 9'h000; 
        10'b0100111000: data <= 9'h000; 
        10'b0100111001: data <= 9'h000; 
        10'b0100111010: data <= 9'h000; 
        10'b0100111011: data <= 9'h001; 
        10'b0100111100: data <= 9'h001; 
        10'b0100111101: data <= 9'h000; 
        10'b0100111110: data <= 9'h000; 
        10'b0100111111: data <= 9'h000; 
        10'b0101000000: data <= 9'h000; 
        10'b0101000001: data <= 9'h000; 
        10'b0101000010: data <= 9'h1ff; 
        10'b0101000011: data <= 9'h1fe; 
        10'b0101000100: data <= 9'h1fe; 
        10'b0101000101: data <= 9'h1ff; 
        10'b0101000110: data <= 9'h1ff; 
        10'b0101000111: data <= 9'h1ff; 
        10'b0101001000: data <= 9'h1ff; 
        10'b0101001001: data <= 9'h000; 
        10'b0101001010: data <= 9'h001; 
        10'b0101001011: data <= 9'h001; 
        10'b0101001100: data <= 9'h000; 
        10'b0101001101: data <= 9'h1ff; 
        10'b0101001110: data <= 9'h000; 
        10'b0101001111: data <= 9'h000; 
        10'b0101010000: data <= 9'h000; 
        10'b0101010001: data <= 9'h000; 
        10'b0101010010: data <= 9'h000; 
        10'b0101010011: data <= 9'h000; 
        10'b0101010100: data <= 9'h000; 
        10'b0101010101: data <= 9'h000; 
        10'b0101010110: data <= 9'h001; 
        10'b0101010111: data <= 9'h001; 
        10'b0101011000: data <= 9'h000; 
        10'b0101011001: data <= 9'h001; 
        10'b0101011010: data <= 9'h000; 
        10'b0101011011: data <= 9'h001; 
        10'b0101011100: data <= 9'h001; 
        10'b0101011101: data <= 9'h001; 
        10'b0101011110: data <= 9'h1ff; 
        10'b0101011111: data <= 9'h1ff; 
        10'b0101100000: data <= 9'h000; 
        10'b0101100001: data <= 9'h000; 
        10'b0101100010: data <= 9'h1ff; 
        10'b0101100011: data <= 9'h1ff; 
        10'b0101100100: data <= 9'h000; 
        10'b0101100101: data <= 9'h001; 
        10'b0101100110: data <= 9'h002; 
        10'b0101100111: data <= 9'h003; 
        10'b0101101000: data <= 9'h001; 
        10'b0101101001: data <= 9'h000; 
        10'b0101101010: data <= 9'h000; 
        10'b0101101011: data <= 9'h000; 
        10'b0101101100: data <= 9'h000; 
        10'b0101101101: data <= 9'h000; 
        10'b0101101110: data <= 9'h000; 
        10'b0101101111: data <= 9'h000; 
        10'b0101110000: data <= 9'h000; 
        10'b0101110001: data <= 9'h000; 
        10'b0101110010: data <= 9'h001; 
        10'b0101110011: data <= 9'h001; 
        10'b0101110100: data <= 9'h001; 
        10'b0101110101: data <= 9'h000; 
        10'b0101110110: data <= 9'h001; 
        10'b0101110111: data <= 9'h001; 
        10'b0101111000: data <= 9'h001; 
        10'b0101111001: data <= 9'h000; 
        10'b0101111010: data <= 9'h000; 
        10'b0101111011: data <= 9'h000; 
        10'b0101111100: data <= 9'h000; 
        10'b0101111101: data <= 9'h000; 
        10'b0101111110: data <= 9'h1ff; 
        10'b0101111111: data <= 9'h000; 
        10'b0110000000: data <= 9'h000; 
        10'b0110000001: data <= 9'h001; 
        10'b0110000010: data <= 9'h002; 
        10'b0110000011: data <= 9'h003; 
        10'b0110000100: data <= 9'h002; 
        10'b0110000101: data <= 9'h000; 
        10'b0110000110: data <= 9'h000; 
        10'b0110000111: data <= 9'h000; 
        10'b0110001000: data <= 9'h000; 
        10'b0110001001: data <= 9'h000; 
        10'b0110001010: data <= 9'h000; 
        10'b0110001011: data <= 9'h000; 
        10'b0110001100: data <= 9'h000; 
        10'b0110001101: data <= 9'h000; 
        10'b0110001110: data <= 9'h001; 
        10'b0110001111: data <= 9'h001; 
        10'b0110010000: data <= 9'h001; 
        10'b0110010001: data <= 9'h001; 
        10'b0110010010: data <= 9'h001; 
        10'b0110010011: data <= 9'h001; 
        10'b0110010100: data <= 9'h000; 
        10'b0110010101: data <= 9'h1ff; 
        10'b0110010110: data <= 9'h000; 
        10'b0110010111: data <= 9'h001; 
        10'b0110011000: data <= 9'h000; 
        10'b0110011001: data <= 9'h000; 
        10'b0110011010: data <= 9'h000; 
        10'b0110011011: data <= 9'h000; 
        10'b0110011100: data <= 9'h001; 
        10'b0110011101: data <= 9'h001; 
        10'b0110011110: data <= 9'h002; 
        10'b0110011111: data <= 9'h003; 
        10'b0110100000: data <= 9'h002; 
        10'b0110100001: data <= 9'h000; 
        10'b0110100010: data <= 9'h1ff; 
        10'b0110100011: data <= 9'h000; 
        10'b0110100100: data <= 9'h000; 
        10'b0110100101: data <= 9'h000; 
        10'b0110100110: data <= 9'h000; 
        10'b0110100111: data <= 9'h000; 
        10'b0110101000: data <= 9'h1ff; 
        10'b0110101001: data <= 9'h000; 
        10'b0110101010: data <= 9'h001; 
        10'b0110101011: data <= 9'h001; 
        10'b0110101100: data <= 9'h001; 
        10'b0110101101: data <= 9'h002; 
        10'b0110101110: data <= 9'h002; 
        10'b0110101111: data <= 9'h002; 
        10'b0110110000: data <= 9'h001; 
        10'b0110110001: data <= 9'h000; 
        10'b0110110010: data <= 9'h001; 
        10'b0110110011: data <= 9'h001; 
        10'b0110110100: data <= 9'h000; 
        10'b0110110101: data <= 9'h000; 
        10'b0110110110: data <= 9'h000; 
        10'b0110110111: data <= 9'h000; 
        10'b0110111000: data <= 9'h001; 
        10'b0110111001: data <= 9'h001; 
        10'b0110111010: data <= 9'h001; 
        10'b0110111011: data <= 9'h002; 
        10'b0110111100: data <= 9'h001; 
        10'b0110111101: data <= 9'h000; 
        10'b0110111110: data <= 9'h000; 
        10'b0110111111: data <= 9'h000; 
        10'b0111000000: data <= 9'h000; 
        10'b0111000001: data <= 9'h000; 
        10'b0111000010: data <= 9'h000; 
        10'b0111000011: data <= 9'h000; 
        10'b0111000100: data <= 9'h1ff; 
        10'b0111000101: data <= 9'h1ff; 
        10'b0111000110: data <= 9'h002; 
        10'b0111000111: data <= 9'h002; 
        10'b0111001000: data <= 9'h001; 
        10'b0111001001: data <= 9'h002; 
        10'b0111001010: data <= 9'h003; 
        10'b0111001011: data <= 9'h003; 
        10'b0111001100: data <= 9'h001; 
        10'b0111001101: data <= 9'h001; 
        10'b0111001110: data <= 9'h001; 
        10'b0111001111: data <= 9'h001; 
        10'b0111010000: data <= 9'h000; 
        10'b0111010001: data <= 9'h1ff; 
        10'b0111010010: data <= 9'h000; 
        10'b0111010011: data <= 9'h001; 
        10'b0111010100: data <= 9'h000; 
        10'b0111010101: data <= 9'h000; 
        10'b0111010110: data <= 9'h001; 
        10'b0111010111: data <= 9'h000; 
        10'b0111011000: data <= 9'h000; 
        10'b0111011001: data <= 9'h1ff; 
        10'b0111011010: data <= 9'h000; 
        10'b0111011011: data <= 9'h000; 
        10'b0111011100: data <= 9'h000; 
        10'b0111011101: data <= 9'h000; 
        10'b0111011110: data <= 9'h000; 
        10'b0111011111: data <= 9'h000; 
        10'b0111100000: data <= 9'h1ff; 
        10'b0111100001: data <= 9'h1ff; 
        10'b0111100010: data <= 9'h001; 
        10'b0111100011: data <= 9'h001; 
        10'b0111100100: data <= 9'h002; 
        10'b0111100101: data <= 9'h002; 
        10'b0111100110: data <= 9'h003; 
        10'b0111100111: data <= 9'h003; 
        10'b0111101000: data <= 9'h002; 
        10'b0111101001: data <= 9'h001; 
        10'b0111101010: data <= 9'h001; 
        10'b0111101011: data <= 9'h001; 
        10'b0111101100: data <= 9'h000; 
        10'b0111101101: data <= 9'h000; 
        10'b0111101110: data <= 9'h001; 
        10'b0111101111: data <= 9'h000; 
        10'b0111110000: data <= 9'h000; 
        10'b0111110001: data <= 9'h000; 
        10'b0111110010: data <= 9'h000; 
        10'b0111110011: data <= 9'h000; 
        10'b0111110100: data <= 9'h000; 
        10'b0111110101: data <= 9'h1ff; 
        10'b0111110110: data <= 9'h000; 
        10'b0111110111: data <= 9'h000; 
        10'b0111111000: data <= 9'h000; 
        10'b0111111001: data <= 9'h000; 
        10'b0111111010: data <= 9'h000; 
        10'b0111111011: data <= 9'h000; 
        10'b0111111100: data <= 9'h1ff; 
        10'b0111111101: data <= 9'h1ff; 
        10'b0111111110: data <= 9'h1ff; 
        10'b0111111111: data <= 9'h001; 
        10'b1000000000: data <= 9'h001; 
        10'b1000000001: data <= 9'h001; 
        10'b1000000010: data <= 9'h002; 
        10'b1000000011: data <= 9'h003; 
        10'b1000000100: data <= 9'h003; 
        10'b1000000101: data <= 9'h002; 
        10'b1000000110: data <= 9'h000; 
        10'b1000000111: data <= 9'h001; 
        10'b1000001000: data <= 9'h001; 
        10'b1000001001: data <= 9'h001; 
        10'b1000001010: data <= 9'h001; 
        10'b1000001011: data <= 9'h001; 
        10'b1000001100: data <= 9'h000; 
        10'b1000001101: data <= 9'h000; 
        10'b1000001110: data <= 9'h000; 
        10'b1000001111: data <= 9'h000; 
        10'b1000010000: data <= 9'h000; 
        10'b1000010001: data <= 9'h000; 
        10'b1000010010: data <= 9'h000; 
        10'b1000010011: data <= 9'h000; 
        10'b1000010100: data <= 9'h000; 
        10'b1000010101: data <= 9'h000; 
        10'b1000010110: data <= 9'h000; 
        10'b1000010111: data <= 9'h1ff; 
        10'b1000011000: data <= 9'h1ff; 
        10'b1000011001: data <= 9'h1ff; 
        10'b1000011010: data <= 9'h1ff; 
        10'b1000011011: data <= 9'h000; 
        10'b1000011100: data <= 9'h001; 
        10'b1000011101: data <= 9'h001; 
        10'b1000011110: data <= 9'h002; 
        10'b1000011111: data <= 9'h003; 
        10'b1000100000: data <= 9'h004; 
        10'b1000100001: data <= 9'h002; 
        10'b1000100010: data <= 9'h002; 
        10'b1000100011: data <= 9'h002; 
        10'b1000100100: data <= 9'h001; 
        10'b1000100101: data <= 9'h001; 
        10'b1000100110: data <= 9'h002; 
        10'b1000100111: data <= 9'h001; 
        10'b1000101000: data <= 9'h001; 
        10'b1000101001: data <= 9'h000; 
        10'b1000101010: data <= 9'h000; 
        10'b1000101011: data <= 9'h000; 
        10'b1000101100: data <= 9'h000; 
        10'b1000101101: data <= 9'h000; 
        10'b1000101110: data <= 9'h000; 
        10'b1000101111: data <= 9'h000; 
        10'b1000110000: data <= 9'h000; 
        10'b1000110001: data <= 9'h000; 
        10'b1000110010: data <= 9'h000; 
        10'b1000110011: data <= 9'h000; 
        10'b1000110100: data <= 9'h1ff; 
        10'b1000110101: data <= 9'h1ff; 
        10'b1000110110: data <= 9'h1ff; 
        10'b1000110111: data <= 9'h000; 
        10'b1000111000: data <= 9'h000; 
        10'b1000111001: data <= 9'h001; 
        10'b1000111010: data <= 9'h002; 
        10'b1000111011: data <= 9'h001; 
        10'b1000111100: data <= 9'h002; 
        10'b1000111101: data <= 9'h003; 
        10'b1000111110: data <= 9'h003; 
        10'b1000111111: data <= 9'h003; 
        10'b1001000000: data <= 9'h001; 
        10'b1001000001: data <= 9'h001; 
        10'b1001000010: data <= 9'h002; 
        10'b1001000011: data <= 9'h001; 
        10'b1001000100: data <= 9'h001; 
        10'b1001000101: data <= 9'h000; 
        10'b1001000110: data <= 9'h1ff; 
        10'b1001000111: data <= 9'h000; 
        10'b1001001000: data <= 9'h000; 
        10'b1001001001: data <= 9'h000; 
        10'b1001001010: data <= 9'h000; 
        10'b1001001011: data <= 9'h000; 
        10'b1001001100: data <= 9'h000; 
        10'b1001001101: data <= 9'h000; 
        10'b1001001110: data <= 9'h000; 
        10'b1001001111: data <= 9'h000; 
        10'b1001010000: data <= 9'h000; 
        10'b1001010001: data <= 9'h1ff; 
        10'b1001010010: data <= 9'h1fe; 
        10'b1001010011: data <= 9'h1ff; 
        10'b1001010100: data <= 9'h000; 
        10'b1001010101: data <= 9'h001; 
        10'b1001010110: data <= 9'h001; 
        10'b1001010111: data <= 9'h002; 
        10'b1001011000: data <= 9'h002; 
        10'b1001011001: data <= 9'h003; 
        10'b1001011010: data <= 9'h002; 
        10'b1001011011: data <= 9'h002; 
        10'b1001011100: data <= 9'h001; 
        10'b1001011101: data <= 9'h002; 
        10'b1001011110: data <= 9'h001; 
        10'b1001011111: data <= 9'h001; 
        10'b1001100000: data <= 9'h000; 
        10'b1001100001: data <= 9'h000; 
        10'b1001100010: data <= 9'h1ff; 
        10'b1001100011: data <= 9'h000; 
        10'b1001100100: data <= 9'h000; 
        10'b1001100101: data <= 9'h000; 
        10'b1001100110: data <= 9'h000; 
        10'b1001100111: data <= 9'h000; 
        10'b1001101000: data <= 9'h000; 
        10'b1001101001: data <= 9'h000; 
        10'b1001101010: data <= 9'h000; 
        10'b1001101011: data <= 9'h000; 
        10'b1001101100: data <= 9'h000; 
        10'b1001101101: data <= 9'h1ff; 
        10'b1001101110: data <= 9'h1ff; 
        10'b1001101111: data <= 9'h1ff; 
        10'b1001110000: data <= 9'h1ff; 
        10'b1001110001: data <= 9'h000; 
        10'b1001110010: data <= 9'h000; 
        10'b1001110011: data <= 9'h000; 
        10'b1001110100: data <= 9'h001; 
        10'b1001110101: data <= 9'h000; 
        10'b1001110110: data <= 9'h000; 
        10'b1001110111: data <= 9'h001; 
        10'b1001111000: data <= 9'h001; 
        10'b1001111001: data <= 9'h000; 
        10'b1001111010: data <= 9'h000; 
        10'b1001111011: data <= 9'h1ff; 
        10'b1001111100: data <= 9'h1ff; 
        10'b1001111101: data <= 9'h1ff; 
        10'b1001111110: data <= 9'h1ff; 
        10'b1001111111: data <= 9'h000; 
        10'b1010000000: data <= 9'h000; 
        10'b1010000001: data <= 9'h000; 
        10'b1010000010: data <= 9'h000; 
        10'b1010000011: data <= 9'h000; 
        10'b1010000100: data <= 9'h000; 
        10'b1010000101: data <= 9'h000; 
        10'b1010000110: data <= 9'h000; 
        10'b1010000111: data <= 9'h000; 
        10'b1010001000: data <= 9'h000; 
        10'b1010001001: data <= 9'h000; 
        10'b1010001010: data <= 9'h1ff; 
        10'b1010001011: data <= 9'h1ff; 
        10'b1010001100: data <= 9'h1ff; 
        10'b1010001101: data <= 9'h1fe; 
        10'b1010001110: data <= 9'h1fe; 
        10'b1010001111: data <= 9'h1fe; 
        10'b1010010000: data <= 9'h1ff; 
        10'b1010010001: data <= 9'h1ff; 
        10'b1010010010: data <= 9'h1ff; 
        10'b1010010011: data <= 9'h1ff; 
        10'b1010010100: data <= 9'h1fe; 
        10'b1010010101: data <= 9'h1fe; 
        10'b1010010110: data <= 9'h1fe; 
        10'b1010010111: data <= 9'h1ff; 
        10'b1010011000: data <= 9'h1ff; 
        10'b1010011001: data <= 9'h1ff; 
        10'b1010011010: data <= 9'h000; 
        10'b1010011011: data <= 9'h000; 
        10'b1010011100: data <= 9'h000; 
        10'b1010011101: data <= 9'h000; 
        10'b1010011110: data <= 9'h000; 
        10'b1010011111: data <= 9'h000; 
        10'b1010100000: data <= 9'h000; 
        10'b1010100001: data <= 9'h000; 
        10'b1010100010: data <= 9'h000; 
        10'b1010100011: data <= 9'h000; 
        10'b1010100100: data <= 9'h000; 
        10'b1010100101: data <= 9'h000; 
        10'b1010100110: data <= 9'h000; 
        10'b1010100111: data <= 9'h000; 
        10'b1010101000: data <= 9'h000; 
        10'b1010101001: data <= 9'h000; 
        10'b1010101010: data <= 9'h1ff; 
        10'b1010101011: data <= 9'h1ff; 
        10'b1010101100: data <= 9'h1ff; 
        10'b1010101101: data <= 9'h1ff; 
        10'b1010101110: data <= 9'h1ff; 
        10'b1010101111: data <= 9'h1ff; 
        10'b1010110000: data <= 9'h1ff; 
        10'b1010110001: data <= 9'h1ff; 
        10'b1010110010: data <= 9'h000; 
        10'b1010110011: data <= 9'h000; 
        10'b1010110100: data <= 9'h000; 
        10'b1010110101: data <= 9'h000; 
        10'b1010110110: data <= 9'h000; 
        10'b1010110111: data <= 9'h000; 
        10'b1010111000: data <= 9'h000; 
        10'b1010111001: data <= 9'h000; 
        10'b1010111010: data <= 9'h000; 
        10'b1010111011: data <= 9'h000; 
        10'b1010111100: data <= 9'h000; 
        10'b1010111101: data <= 9'h000; 
        10'b1010111110: data <= 9'h000; 
        10'b1010111111: data <= 9'h000; 
        10'b1011000000: data <= 9'h000; 
        10'b1011000001: data <= 9'h000; 
        10'b1011000010: data <= 9'h000; 
        10'b1011000011: data <= 9'h000; 
        10'b1011000100: data <= 9'h000; 
        10'b1011000101: data <= 9'h000; 
        10'b1011000110: data <= 9'h000; 
        10'b1011000111: data <= 9'h000; 
        10'b1011001000: data <= 9'h000; 
        10'b1011001001: data <= 9'h000; 
        10'b1011001010: data <= 9'h000; 
        10'b1011001011: data <= 9'h000; 
        10'b1011001100: data <= 9'h000; 
        10'b1011001101: data <= 9'h000; 
        10'b1011001110: data <= 9'h000; 
        10'b1011001111: data <= 9'h000; 
        10'b1011010000: data <= 9'h000; 
        10'b1011010001: data <= 9'h000; 
        10'b1011010010: data <= 9'h000; 
        10'b1011010011: data <= 9'h000; 
        10'b1011010100: data <= 9'h000; 
        10'b1011010101: data <= 9'h000; 
        10'b1011010110: data <= 9'h000; 
        10'b1011010111: data <= 9'h000; 
        10'b1011011000: data <= 9'h000; 
        10'b1011011001: data <= 9'h000; 
        10'b1011011010: data <= 9'h000; 
        10'b1011011011: data <= 9'h000; 
        10'b1011011100: data <= 9'h000; 
        10'b1011011101: data <= 9'h000; 
        10'b1011011110: data <= 9'h000; 
        10'b1011011111: data <= 9'h000; 
        10'b1011100000: data <= 9'h000; 
        10'b1011100001: data <= 9'h000; 
        10'b1011100010: data <= 9'h000; 
        10'b1011100011: data <= 9'h000; 
        10'b1011100100: data <= 9'h000; 
        10'b1011100101: data <= 9'h000; 
        10'b1011100110: data <= 9'h000; 
        10'b1011100111: data <= 9'h000; 
        10'b1011101000: data <= 9'h000; 
        10'b1011101001: data <= 9'h000; 
        10'b1011101010: data <= 9'h000; 
        10'b1011101011: data <= 9'h000; 
        10'b1011101100: data <= 9'h000; 
        10'b1011101101: data <= 9'h000; 
        10'b1011101110: data <= 9'h000; 
        10'b1011101111: data <= 9'h000; 
        10'b1011110000: data <= 9'h000; 
        10'b1011110001: data <= 9'h000; 
        10'b1011110010: data <= 9'h000; 
        10'b1011110011: data <= 9'h000; 
        10'b1011110100: data <= 9'h000; 
        10'b1011110101: data <= 9'h000; 
        10'b1011110110: data <= 9'h000; 
        10'b1011110111: data <= 9'h000; 
        10'b1011111000: data <= 9'h000; 
        10'b1011111001: data <= 9'h000; 
        10'b1011111010: data <= 9'h000; 
        10'b1011111011: data <= 9'h000; 
        10'b1011111100: data <= 9'h000; 
        10'b1011111101: data <= 9'h000; 
        10'b1011111110: data <= 9'h000; 
        10'b1011111111: data <= 9'h000; 
        10'b1100000000: data <= 9'h000; 
        10'b1100000001: data <= 9'h000; 
        10'b1100000010: data <= 9'h000; 
        10'b1100000011: data <= 9'h000; 
        10'b1100000100: data <= 9'h000; 
        10'b1100000101: data <= 9'h000; 
        10'b1100000110: data <= 9'h000; 
        10'b1100000111: data <= 9'h000; 
        10'b1100001000: data <= 9'h000; 
        10'b1100001001: data <= 9'h000; 
        10'b1100001010: data <= 9'h000; 
        10'b1100001011: data <= 9'h000; 
        10'b1100001100: data <= 9'h000; 
        10'b1100001101: data <= 9'h000; 
        10'b1100001110: data <= 9'h000; 
        10'b1100001111: data <= 9'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 4) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 10'h000; 
        10'b0000000001: data <= 10'h000; 
        10'b0000000010: data <= 10'h000; 
        10'b0000000011: data <= 10'h000; 
        10'b0000000100: data <= 10'h000; 
        10'b0000000101: data <= 10'h000; 
        10'b0000000110: data <= 10'h000; 
        10'b0000000111: data <= 10'h001; 
        10'b0000001000: data <= 10'h000; 
        10'b0000001001: data <= 10'h000; 
        10'b0000001010: data <= 10'h000; 
        10'b0000001011: data <= 10'h000; 
        10'b0000001100: data <= 10'h000; 
        10'b0000001101: data <= 10'h001; 
        10'b0000001110: data <= 10'h000; 
        10'b0000001111: data <= 10'h000; 
        10'b0000010000: data <= 10'h000; 
        10'b0000010001: data <= 10'h001; 
        10'b0000010010: data <= 10'h000; 
        10'b0000010011: data <= 10'h000; 
        10'b0000010100: data <= 10'h000; 
        10'b0000010101: data <= 10'h000; 
        10'b0000010110: data <= 10'h000; 
        10'b0000010111: data <= 10'h001; 
        10'b0000011000: data <= 10'h000; 
        10'b0000011001: data <= 10'h000; 
        10'b0000011010: data <= 10'h000; 
        10'b0000011011: data <= 10'h000; 
        10'b0000011100: data <= 10'h000; 
        10'b0000011101: data <= 10'h000; 
        10'b0000011110: data <= 10'h000; 
        10'b0000011111: data <= 10'h000; 
        10'b0000100000: data <= 10'h3ff; 
        10'b0000100001: data <= 10'h000; 
        10'b0000100010: data <= 10'h000; 
        10'b0000100011: data <= 10'h001; 
        10'b0000100100: data <= 10'h001; 
        10'b0000100101: data <= 10'h000; 
        10'b0000100110: data <= 10'h001; 
        10'b0000100111: data <= 10'h001; 
        10'b0000101000: data <= 10'h001; 
        10'b0000101001: data <= 10'h001; 
        10'b0000101010: data <= 10'h000; 
        10'b0000101011: data <= 10'h000; 
        10'b0000101100: data <= 10'h3ff; 
        10'b0000101101: data <= 10'h000; 
        10'b0000101110: data <= 10'h001; 
        10'b0000101111: data <= 10'h000; 
        10'b0000110000: data <= 10'h000; 
        10'b0000110001: data <= 10'h000; 
        10'b0000110010: data <= 10'h001; 
        10'b0000110011: data <= 10'h001; 
        10'b0000110100: data <= 10'h000; 
        10'b0000110101: data <= 10'h001; 
        10'b0000110110: data <= 10'h000; 
        10'b0000110111: data <= 10'h000; 
        10'b0000111000: data <= 10'h000; 
        10'b0000111001: data <= 10'h000; 
        10'b0000111010: data <= 10'h3ff; 
        10'b0000111011: data <= 10'h000; 
        10'b0000111100: data <= 10'h000; 
        10'b0000111101: data <= 10'h000; 
        10'b0000111110: data <= 10'h000; 
        10'b0000111111: data <= 10'h001; 
        10'b0001000000: data <= 10'h001; 
        10'b0001000001: data <= 10'h001; 
        10'b0001000010: data <= 10'h002; 
        10'b0001000011: data <= 10'h002; 
        10'b0001000100: data <= 10'h002; 
        10'b0001000101: data <= 10'h002; 
        10'b0001000110: data <= 10'h001; 
        10'b0001000111: data <= 10'h001; 
        10'b0001001000: data <= 10'h002; 
        10'b0001001001: data <= 10'h001; 
        10'b0001001010: data <= 10'h001; 
        10'b0001001011: data <= 10'h001; 
        10'b0001001100: data <= 10'h001; 
        10'b0001001101: data <= 10'h000; 
        10'b0001001110: data <= 10'h000; 
        10'b0001001111: data <= 10'h000; 
        10'b0001010000: data <= 10'h000; 
        10'b0001010001: data <= 10'h000; 
        10'b0001010010: data <= 10'h3ff; 
        10'b0001010011: data <= 10'h000; 
        10'b0001010100: data <= 10'h000; 
        10'b0001010101: data <= 10'h000; 
        10'b0001010110: data <= 10'h000; 
        10'b0001010111: data <= 10'h000; 
        10'b0001011000: data <= 10'h001; 
        10'b0001011001: data <= 10'h000; 
        10'b0001011010: data <= 10'h001; 
        10'b0001011011: data <= 10'h001; 
        10'b0001011100: data <= 10'h001; 
        10'b0001011101: data <= 10'h002; 
        10'b0001011110: data <= 10'h001; 
        10'b0001011111: data <= 10'h002; 
        10'b0001100000: data <= 10'h002; 
        10'b0001100001: data <= 10'h002; 
        10'b0001100010: data <= 10'h002; 
        10'b0001100011: data <= 10'h002; 
        10'b0001100100: data <= 10'h001; 
        10'b0001100101: data <= 10'h002; 
        10'b0001100110: data <= 10'h003; 
        10'b0001100111: data <= 10'h003; 
        10'b0001101000: data <= 10'h003; 
        10'b0001101001: data <= 10'h003; 
        10'b0001101010: data <= 10'h003; 
        10'b0001101011: data <= 10'h002; 
        10'b0001101100: data <= 10'h001; 
        10'b0001101101: data <= 10'h000; 
        10'b0001101110: data <= 10'h000; 
        10'b0001101111: data <= 10'h000; 
        10'b0001110000: data <= 10'h000; 
        10'b0001110001: data <= 10'h000; 
        10'b0001110010: data <= 10'h000; 
        10'b0001110011: data <= 10'h000; 
        10'b0001110100: data <= 10'h000; 
        10'b0001110101: data <= 10'h000; 
        10'b0001110110: data <= 10'h000; 
        10'b0001110111: data <= 10'h001; 
        10'b0001111000: data <= 10'h000; 
        10'b0001111001: data <= 10'h000; 
        10'b0001111010: data <= 10'h001; 
        10'b0001111011: data <= 10'h000; 
        10'b0001111100: data <= 10'h000; 
        10'b0001111101: data <= 10'h000; 
        10'b0001111110: data <= 10'h000; 
        10'b0001111111: data <= 10'h001; 
        10'b0010000000: data <= 10'h002; 
        10'b0010000001: data <= 10'h002; 
        10'b0010000010: data <= 10'h003; 
        10'b0010000011: data <= 10'h003; 
        10'b0010000100: data <= 10'h004; 
        10'b0010000101: data <= 10'h004; 
        10'b0010000110: data <= 10'h004; 
        10'b0010000111: data <= 10'h002; 
        10'b0010001000: data <= 10'h000; 
        10'b0010001001: data <= 10'h001; 
        10'b0010001010: data <= 10'h000; 
        10'b0010001011: data <= 10'h000; 
        10'b0010001100: data <= 10'h000; 
        10'b0010001101: data <= 10'h000; 
        10'b0010001110: data <= 10'h000; 
        10'b0010001111: data <= 10'h000; 
        10'b0010010000: data <= 10'h000; 
        10'b0010010001: data <= 10'h000; 
        10'b0010010010: data <= 10'h000; 
        10'b0010010011: data <= 10'h3ff; 
        10'b0010010100: data <= 10'h001; 
        10'b0010010101: data <= 10'h3ff; 
        10'b0010010110: data <= 10'h000; 
        10'b0010010111: data <= 10'h3fe; 
        10'b0010011000: data <= 10'h3ff; 
        10'b0010011001: data <= 10'h3ff; 
        10'b0010011010: data <= 10'h000; 
        10'b0010011011: data <= 10'h3ff; 
        10'b0010011100: data <= 10'h3ff; 
        10'b0010011101: data <= 10'h000; 
        10'b0010011110: data <= 10'h001; 
        10'b0010011111: data <= 10'h003; 
        10'b0010100000: data <= 10'h002; 
        10'b0010100001: data <= 10'h002; 
        10'b0010100010: data <= 10'h002; 
        10'b0010100011: data <= 10'h001; 
        10'b0010100100: data <= 10'h000; 
        10'b0010100101: data <= 10'h000; 
        10'b0010100110: data <= 10'h3ff; 
        10'b0010100111: data <= 10'h001; 
        10'b0010101000: data <= 10'h000; 
        10'b0010101001: data <= 10'h000; 
        10'b0010101010: data <= 10'h000; 
        10'b0010101011: data <= 10'h3ff; 
        10'b0010101100: data <= 10'h000; 
        10'b0010101101: data <= 10'h000; 
        10'b0010101110: data <= 10'h000; 
        10'b0010101111: data <= 10'h000; 
        10'b0010110000: data <= 10'h3ff; 
        10'b0010110001: data <= 10'h3ff; 
        10'b0010110010: data <= 10'h3fd; 
        10'b0010110011: data <= 10'h3fd; 
        10'b0010110100: data <= 10'h3fe; 
        10'b0010110101: data <= 10'h3fc; 
        10'b0010110110: data <= 10'h3fe; 
        10'b0010110111: data <= 10'h3ff; 
        10'b0010111000: data <= 10'h3fe; 
        10'b0010111001: data <= 10'h3fe; 
        10'b0010111010: data <= 10'h000; 
        10'b0010111011: data <= 10'h3ff; 
        10'b0010111100: data <= 10'h3fe; 
        10'b0010111101: data <= 10'h3fe; 
        10'b0010111110: data <= 10'h3fd; 
        10'b0010111111: data <= 10'h3fe; 
        10'b0011000000: data <= 10'h3ff; 
        10'b0011000001: data <= 10'h3ff; 
        10'b0011000010: data <= 10'h000; 
        10'b0011000011: data <= 10'h000; 
        10'b0011000100: data <= 10'h000; 
        10'b0011000101: data <= 10'h000; 
        10'b0011000110: data <= 10'h000; 
        10'b0011000111: data <= 10'h000; 
        10'b0011001000: data <= 10'h000; 
        10'b0011001001: data <= 10'h000; 
        10'b0011001010: data <= 10'h3ff; 
        10'b0011001011: data <= 10'h000; 
        10'b0011001100: data <= 10'h3ff; 
        10'b0011001101: data <= 10'h3fe; 
        10'b0011001110: data <= 10'h3fd; 
        10'b0011001111: data <= 10'h3fe; 
        10'b0011010000: data <= 10'h3fc; 
        10'b0011010001: data <= 10'h3fc; 
        10'b0011010010: data <= 10'h3fe; 
        10'b0011010011: data <= 10'h3fe; 
        10'b0011010100: data <= 10'h3fd; 
        10'b0011010101: data <= 10'h3fd; 
        10'b0011010110: data <= 10'h3fc; 
        10'b0011010111: data <= 10'h3fb; 
        10'b0011011000: data <= 10'h3fb; 
        10'b0011011001: data <= 10'h3fc; 
        10'b0011011010: data <= 10'h3fb; 
        10'b0011011011: data <= 10'h3fc; 
        10'b0011011100: data <= 10'h3ff; 
        10'b0011011101: data <= 10'h3ff; 
        10'b0011011110: data <= 10'h000; 
        10'b0011011111: data <= 10'h000; 
        10'b0011100000: data <= 10'h000; 
        10'b0011100001: data <= 10'h000; 
        10'b0011100010: data <= 10'h001; 
        10'b0011100011: data <= 10'h3ff; 
        10'b0011100100: data <= 10'h3ff; 
        10'b0011100101: data <= 10'h3ff; 
        10'b0011100110: data <= 10'h3fe; 
        10'b0011100111: data <= 10'h000; 
        10'b0011101000: data <= 10'h3ff; 
        10'b0011101001: data <= 10'h3fe; 
        10'b0011101010: data <= 10'h3fe; 
        10'b0011101011: data <= 10'h3fd; 
        10'b0011101100: data <= 10'h3fd; 
        10'b0011101101: data <= 10'h3fc; 
        10'b0011101110: data <= 10'h3fc; 
        10'b0011101111: data <= 10'h3fc; 
        10'b0011110000: data <= 10'h3fb; 
        10'b0011110001: data <= 10'h3fb; 
        10'b0011110010: data <= 10'h3f8; 
        10'b0011110011: data <= 10'h3f9; 
        10'b0011110100: data <= 10'h3fa; 
        10'b0011110101: data <= 10'h3fa; 
        10'b0011110110: data <= 10'h3fc; 
        10'b0011110111: data <= 10'h3fc; 
        10'b0011111000: data <= 10'h3fe; 
        10'b0011111001: data <= 10'h3fe; 
        10'b0011111010: data <= 10'h3ff; 
        10'b0011111011: data <= 10'h000; 
        10'b0011111100: data <= 10'h000; 
        10'b0011111101: data <= 10'h000; 
        10'b0011111110: data <= 10'h000; 
        10'b0011111111: data <= 10'h000; 
        10'b0100000000: data <= 10'h000; 
        10'b0100000001: data <= 10'h000; 
        10'b0100000010: data <= 10'h3ff; 
        10'b0100000011: data <= 10'h000; 
        10'b0100000100: data <= 10'h000; 
        10'b0100000101: data <= 10'h3ff; 
        10'b0100000110: data <= 10'h3fe; 
        10'b0100000111: data <= 10'h3fe; 
        10'b0100001000: data <= 10'h3ff; 
        10'b0100001001: data <= 10'h3fe; 
        10'b0100001010: data <= 10'h3fe; 
        10'b0100001011: data <= 10'h3fc; 
        10'b0100001100: data <= 10'h3fb; 
        10'b0100001101: data <= 10'h3f9; 
        10'b0100001110: data <= 10'h3f8; 
        10'b0100001111: data <= 10'h3fa; 
        10'b0100010000: data <= 10'h3fb; 
        10'b0100010001: data <= 10'h3fc; 
        10'b0100010010: data <= 10'h3fb; 
        10'b0100010011: data <= 10'h3fd; 
        10'b0100010100: data <= 10'h3fe; 
        10'b0100010101: data <= 10'h3fe; 
        10'b0100010110: data <= 10'h3ff; 
        10'b0100010111: data <= 10'h000; 
        10'b0100011000: data <= 10'h000; 
        10'b0100011001: data <= 10'h000; 
        10'b0100011010: data <= 10'h000; 
        10'b0100011011: data <= 10'h3ff; 
        10'b0100011100: data <= 10'h3ff; 
        10'b0100011101: data <= 10'h000; 
        10'b0100011110: data <= 10'h001; 
        10'b0100011111: data <= 10'h001; 
        10'b0100100000: data <= 10'h002; 
        10'b0100100001: data <= 10'h000; 
        10'b0100100010: data <= 10'h000; 
        10'b0100100011: data <= 10'h000; 
        10'b0100100100: data <= 10'h3ff; 
        10'b0100100101: data <= 10'h3ff; 
        10'b0100100110: data <= 10'h3fe; 
        10'b0100100111: data <= 10'h3fc; 
        10'b0100101000: data <= 10'h3fb; 
        10'b0100101001: data <= 10'h3fb; 
        10'b0100101010: data <= 10'h3fa; 
        10'b0100101011: data <= 10'h3fc; 
        10'b0100101100: data <= 10'h3fd; 
        10'b0100101101: data <= 10'h3fe; 
        10'b0100101110: data <= 10'h3fd; 
        10'b0100101111: data <= 10'h000; 
        10'b0100110000: data <= 10'h3fe; 
        10'b0100110001: data <= 10'h3ff; 
        10'b0100110010: data <= 10'h000; 
        10'b0100110011: data <= 10'h000; 
        10'b0100110100: data <= 10'h000; 
        10'b0100110101: data <= 10'h000; 
        10'b0100110110: data <= 10'h000; 
        10'b0100110111: data <= 10'h000; 
        10'b0100111000: data <= 10'h000; 
        10'b0100111001: data <= 10'h000; 
        10'b0100111010: data <= 10'h000; 
        10'b0100111011: data <= 10'h002; 
        10'b0100111100: data <= 10'h001; 
        10'b0100111101: data <= 10'h001; 
        10'b0100111110: data <= 10'h001; 
        10'b0100111111: data <= 10'h001; 
        10'b0101000000: data <= 10'h001; 
        10'b0101000001: data <= 10'h000; 
        10'b0101000010: data <= 10'h3ff; 
        10'b0101000011: data <= 10'h3fc; 
        10'b0101000100: data <= 10'h3fd; 
        10'b0101000101: data <= 10'h3fd; 
        10'b0101000110: data <= 10'h3fd; 
        10'b0101000111: data <= 10'h3fe; 
        10'b0101001000: data <= 10'h3ff; 
        10'b0101001001: data <= 10'h000; 
        10'b0101001010: data <= 10'h001; 
        10'b0101001011: data <= 10'h002; 
        10'b0101001100: data <= 10'h000; 
        10'b0101001101: data <= 10'h3ff; 
        10'b0101001110: data <= 10'h000; 
        10'b0101001111: data <= 10'h000; 
        10'b0101010000: data <= 10'h000; 
        10'b0101010001: data <= 10'h000; 
        10'b0101010010: data <= 10'h000; 
        10'b0101010011: data <= 10'h000; 
        10'b0101010100: data <= 10'h000; 
        10'b0101010101: data <= 10'h001; 
        10'b0101010110: data <= 10'h001; 
        10'b0101010111: data <= 10'h002; 
        10'b0101011000: data <= 10'h001; 
        10'b0101011001: data <= 10'h001; 
        10'b0101011010: data <= 10'h001; 
        10'b0101011011: data <= 10'h002; 
        10'b0101011100: data <= 10'h002; 
        10'b0101011101: data <= 10'h002; 
        10'b0101011110: data <= 10'h3ff; 
        10'b0101011111: data <= 10'h3fe; 
        10'b0101100000: data <= 10'h000; 
        10'b0101100001: data <= 10'h000; 
        10'b0101100010: data <= 10'h3fe; 
        10'b0101100011: data <= 10'h3fe; 
        10'b0101100100: data <= 10'h000; 
        10'b0101100101: data <= 10'h001; 
        10'b0101100110: data <= 10'h003; 
        10'b0101100111: data <= 10'h005; 
        10'b0101101000: data <= 10'h003; 
        10'b0101101001: data <= 10'h3ff; 
        10'b0101101010: data <= 10'h3ff; 
        10'b0101101011: data <= 10'h000; 
        10'b0101101100: data <= 10'h000; 
        10'b0101101101: data <= 10'h001; 
        10'b0101101110: data <= 10'h000; 
        10'b0101101111: data <= 10'h3ff; 
        10'b0101110000: data <= 10'h3ff; 
        10'b0101110001: data <= 10'h000; 
        10'b0101110010: data <= 10'h002; 
        10'b0101110011: data <= 10'h001; 
        10'b0101110100: data <= 10'h001; 
        10'b0101110101: data <= 10'h001; 
        10'b0101110110: data <= 10'h002; 
        10'b0101110111: data <= 10'h002; 
        10'b0101111000: data <= 10'h002; 
        10'b0101111001: data <= 10'h000; 
        10'b0101111010: data <= 10'h000; 
        10'b0101111011: data <= 10'h000; 
        10'b0101111100: data <= 10'h000; 
        10'b0101111101: data <= 10'h3ff; 
        10'b0101111110: data <= 10'h3fe; 
        10'b0101111111: data <= 10'h000; 
        10'b0110000000: data <= 10'h3ff; 
        10'b0110000001: data <= 10'h002; 
        10'b0110000010: data <= 10'h004; 
        10'b0110000011: data <= 10'h007; 
        10'b0110000100: data <= 10'h004; 
        10'b0110000101: data <= 10'h000; 
        10'b0110000110: data <= 10'h000; 
        10'b0110000111: data <= 10'h000; 
        10'b0110001000: data <= 10'h000; 
        10'b0110001001: data <= 10'h000; 
        10'b0110001010: data <= 10'h000; 
        10'b0110001011: data <= 10'h000; 
        10'b0110001100: data <= 10'h3ff; 
        10'b0110001101: data <= 10'h001; 
        10'b0110001110: data <= 10'h002; 
        10'b0110001111: data <= 10'h002; 
        10'b0110010000: data <= 10'h003; 
        10'b0110010001: data <= 10'h002; 
        10'b0110010010: data <= 10'h003; 
        10'b0110010011: data <= 10'h003; 
        10'b0110010100: data <= 10'h001; 
        10'b0110010101: data <= 10'h3ff; 
        10'b0110010110: data <= 10'h000; 
        10'b0110010111: data <= 10'h001; 
        10'b0110011000: data <= 10'h001; 
        10'b0110011001: data <= 10'h3ff; 
        10'b0110011010: data <= 10'h3ff; 
        10'b0110011011: data <= 10'h000; 
        10'b0110011100: data <= 10'h002; 
        10'b0110011101: data <= 10'h002; 
        10'b0110011110: data <= 10'h005; 
        10'b0110011111: data <= 10'h006; 
        10'b0110100000: data <= 10'h004; 
        10'b0110100001: data <= 10'h000; 
        10'b0110100010: data <= 10'h3ff; 
        10'b0110100011: data <= 10'h3ff; 
        10'b0110100100: data <= 10'h000; 
        10'b0110100101: data <= 10'h000; 
        10'b0110100110: data <= 10'h000; 
        10'b0110100111: data <= 10'h000; 
        10'b0110101000: data <= 10'h3fe; 
        10'b0110101001: data <= 10'h000; 
        10'b0110101010: data <= 10'h002; 
        10'b0110101011: data <= 10'h003; 
        10'b0110101100: data <= 10'h002; 
        10'b0110101101: data <= 10'h003; 
        10'b0110101110: data <= 10'h004; 
        10'b0110101111: data <= 10'h005; 
        10'b0110110000: data <= 10'h001; 
        10'b0110110001: data <= 10'h000; 
        10'b0110110010: data <= 10'h002; 
        10'b0110110011: data <= 10'h002; 
        10'b0110110100: data <= 10'h000; 
        10'b0110110101: data <= 10'h3ff; 
        10'b0110110110: data <= 10'h000; 
        10'b0110110111: data <= 10'h001; 
        10'b0110111000: data <= 10'h002; 
        10'b0110111001: data <= 10'h003; 
        10'b0110111010: data <= 10'h003; 
        10'b0110111011: data <= 10'h003; 
        10'b0110111100: data <= 10'h002; 
        10'b0110111101: data <= 10'h3ff; 
        10'b0110111110: data <= 10'h3ff; 
        10'b0110111111: data <= 10'h3ff; 
        10'b0111000000: data <= 10'h000; 
        10'b0111000001: data <= 10'h000; 
        10'b0111000010: data <= 10'h000; 
        10'b0111000011: data <= 10'h000; 
        10'b0111000100: data <= 10'h3fe; 
        10'b0111000101: data <= 10'h3ff; 
        10'b0111000110: data <= 10'h003; 
        10'b0111000111: data <= 10'h003; 
        10'b0111001000: data <= 10'h002; 
        10'b0111001001: data <= 10'h003; 
        10'b0111001010: data <= 10'h006; 
        10'b0111001011: data <= 10'h006; 
        10'b0111001100: data <= 10'h002; 
        10'b0111001101: data <= 10'h001; 
        10'b0111001110: data <= 10'h003; 
        10'b0111001111: data <= 10'h001; 
        10'b0111010000: data <= 10'h3ff; 
        10'b0111010001: data <= 10'h3ff; 
        10'b0111010010: data <= 10'h000; 
        10'b0111010011: data <= 10'h001; 
        10'b0111010100: data <= 10'h001; 
        10'b0111010101: data <= 10'h000; 
        10'b0111010110: data <= 10'h001; 
        10'b0111010111: data <= 10'h001; 
        10'b0111011000: data <= 10'h000; 
        10'b0111011001: data <= 10'h3ff; 
        10'b0111011010: data <= 10'h3ff; 
        10'b0111011011: data <= 10'h000; 
        10'b0111011100: data <= 10'h000; 
        10'b0111011101: data <= 10'h000; 
        10'b0111011110: data <= 10'h000; 
        10'b0111011111: data <= 10'h000; 
        10'b0111100000: data <= 10'h3fd; 
        10'b0111100001: data <= 10'h3ff; 
        10'b0111100010: data <= 10'h001; 
        10'b0111100011: data <= 10'h003; 
        10'b0111100100: data <= 10'h003; 
        10'b0111100101: data <= 10'h004; 
        10'b0111100110: data <= 10'h007; 
        10'b0111100111: data <= 10'h007; 
        10'b0111101000: data <= 10'h003; 
        10'b0111101001: data <= 10'h002; 
        10'b0111101010: data <= 10'h002; 
        10'b0111101011: data <= 10'h001; 
        10'b0111101100: data <= 10'h000; 
        10'b0111101101: data <= 10'h000; 
        10'b0111101110: data <= 10'h003; 
        10'b0111101111: data <= 10'h001; 
        10'b0111110000: data <= 10'h000; 
        10'b0111110001: data <= 10'h3ff; 
        10'b0111110010: data <= 10'h001; 
        10'b0111110011: data <= 10'h000; 
        10'b0111110100: data <= 10'h3ff; 
        10'b0111110101: data <= 10'h3fe; 
        10'b0111110110: data <= 10'h000; 
        10'b0111110111: data <= 10'h000; 
        10'b0111111000: data <= 10'h000; 
        10'b0111111001: data <= 10'h000; 
        10'b0111111010: data <= 10'h000; 
        10'b0111111011: data <= 10'h3ff; 
        10'b0111111100: data <= 10'h3fd; 
        10'b0111111101: data <= 10'h3fd; 
        10'b0111111110: data <= 10'h3ff; 
        10'b0111111111: data <= 10'h002; 
        10'b1000000000: data <= 10'h003; 
        10'b1000000001: data <= 10'h003; 
        10'b1000000010: data <= 10'h005; 
        10'b1000000011: data <= 10'h006; 
        10'b1000000100: data <= 10'h007; 
        10'b1000000101: data <= 10'h003; 
        10'b1000000110: data <= 10'h001; 
        10'b1000000111: data <= 10'h002; 
        10'b1000001000: data <= 10'h003; 
        10'b1000001001: data <= 10'h002; 
        10'b1000001010: data <= 10'h002; 
        10'b1000001011: data <= 10'h001; 
        10'b1000001100: data <= 10'h000; 
        10'b1000001101: data <= 10'h000; 
        10'b1000001110: data <= 10'h000; 
        10'b1000001111: data <= 10'h000; 
        10'b1000010000: data <= 10'h3ff; 
        10'b1000010001: data <= 10'h3ff; 
        10'b1000010010: data <= 10'h3ff; 
        10'b1000010011: data <= 10'h3ff; 
        10'b1000010100: data <= 10'h000; 
        10'b1000010101: data <= 10'h000; 
        10'b1000010110: data <= 10'h000; 
        10'b1000010111: data <= 10'h3ff; 
        10'b1000011000: data <= 10'h3fe; 
        10'b1000011001: data <= 10'h3fd; 
        10'b1000011010: data <= 10'h3fe; 
        10'b1000011011: data <= 10'h000; 
        10'b1000011100: data <= 10'h002; 
        10'b1000011101: data <= 10'h003; 
        10'b1000011110: data <= 10'h004; 
        10'b1000011111: data <= 10'h006; 
        10'b1000100000: data <= 10'h007; 
        10'b1000100001: data <= 10'h004; 
        10'b1000100010: data <= 10'h003; 
        10'b1000100011: data <= 10'h003; 
        10'b1000100100: data <= 10'h002; 
        10'b1000100101: data <= 10'h002; 
        10'b1000100110: data <= 10'h003; 
        10'b1000100111: data <= 10'h002; 
        10'b1000101000: data <= 10'h001; 
        10'b1000101001: data <= 10'h000; 
        10'b1000101010: data <= 10'h000; 
        10'b1000101011: data <= 10'h3ff; 
        10'b1000101100: data <= 10'h3ff; 
        10'b1000101101: data <= 10'h000; 
        10'b1000101110: data <= 10'h000; 
        10'b1000101111: data <= 10'h000; 
        10'b1000110000: data <= 10'h000; 
        10'b1000110001: data <= 10'h000; 
        10'b1000110010: data <= 10'h000; 
        10'b1000110011: data <= 10'h000; 
        10'b1000110100: data <= 10'h3fe; 
        10'b1000110101: data <= 10'h3fd; 
        10'b1000110110: data <= 10'h3fe; 
        10'b1000110111: data <= 10'h3ff; 
        10'b1000111000: data <= 10'h001; 
        10'b1000111001: data <= 10'h002; 
        10'b1000111010: data <= 10'h003; 
        10'b1000111011: data <= 10'h002; 
        10'b1000111100: data <= 10'h004; 
        10'b1000111101: data <= 10'h005; 
        10'b1000111110: data <= 10'h006; 
        10'b1000111111: data <= 10'h005; 
        10'b1001000000: data <= 10'h003; 
        10'b1001000001: data <= 10'h002; 
        10'b1001000010: data <= 10'h004; 
        10'b1001000011: data <= 10'h002; 
        10'b1001000100: data <= 10'h002; 
        10'b1001000101: data <= 10'h000; 
        10'b1001000110: data <= 10'h3ff; 
        10'b1001000111: data <= 10'h000; 
        10'b1001001000: data <= 10'h000; 
        10'b1001001001: data <= 10'h000; 
        10'b1001001010: data <= 10'h000; 
        10'b1001001011: data <= 10'h000; 
        10'b1001001100: data <= 10'h000; 
        10'b1001001101: data <= 10'h000; 
        10'b1001001110: data <= 10'h000; 
        10'b1001001111: data <= 10'h000; 
        10'b1001010000: data <= 10'h3ff; 
        10'b1001010001: data <= 10'h3fe; 
        10'b1001010010: data <= 10'h3fd; 
        10'b1001010011: data <= 10'h3ff; 
        10'b1001010100: data <= 10'h3ff; 
        10'b1001010101: data <= 10'h002; 
        10'b1001010110: data <= 10'h003; 
        10'b1001010111: data <= 10'h004; 
        10'b1001011000: data <= 10'h005; 
        10'b1001011001: data <= 10'h005; 
        10'b1001011010: data <= 10'h004; 
        10'b1001011011: data <= 10'h004; 
        10'b1001011100: data <= 10'h002; 
        10'b1001011101: data <= 10'h003; 
        10'b1001011110: data <= 10'h003; 
        10'b1001011111: data <= 10'h002; 
        10'b1001100000: data <= 10'h000; 
        10'b1001100001: data <= 10'h3ff; 
        10'b1001100010: data <= 10'h3ff; 
        10'b1001100011: data <= 10'h3ff; 
        10'b1001100100: data <= 10'h000; 
        10'b1001100101: data <= 10'h3ff; 
        10'b1001100110: data <= 10'h000; 
        10'b1001100111: data <= 10'h000; 
        10'b1001101000: data <= 10'h000; 
        10'b1001101001: data <= 10'h000; 
        10'b1001101010: data <= 10'h000; 
        10'b1001101011: data <= 10'h000; 
        10'b1001101100: data <= 10'h000; 
        10'b1001101101: data <= 10'h3fe; 
        10'b1001101110: data <= 10'h3fe; 
        10'b1001101111: data <= 10'h3fd; 
        10'b1001110000: data <= 10'h3fe; 
        10'b1001110001: data <= 10'h3ff; 
        10'b1001110010: data <= 10'h3ff; 
        10'b1001110011: data <= 10'h000; 
        10'b1001110100: data <= 10'h001; 
        10'b1001110101: data <= 10'h001; 
        10'b1001110110: data <= 10'h001; 
        10'b1001110111: data <= 10'h002; 
        10'b1001111000: data <= 10'h001; 
        10'b1001111001: data <= 10'h000; 
        10'b1001111010: data <= 10'h000; 
        10'b1001111011: data <= 10'h3fe; 
        10'b1001111100: data <= 10'h3fe; 
        10'b1001111101: data <= 10'h3ff; 
        10'b1001111110: data <= 10'h3ff; 
        10'b1001111111: data <= 10'h000; 
        10'b1010000000: data <= 10'h000; 
        10'b1010000001: data <= 10'h000; 
        10'b1010000010: data <= 10'h001; 
        10'b1010000011: data <= 10'h000; 
        10'b1010000100: data <= 10'h000; 
        10'b1010000101: data <= 10'h000; 
        10'b1010000110: data <= 10'h000; 
        10'b1010000111: data <= 10'h000; 
        10'b1010001000: data <= 10'h000; 
        10'b1010001001: data <= 10'h3ff; 
        10'b1010001010: data <= 10'h3ff; 
        10'b1010001011: data <= 10'h3fe; 
        10'b1010001100: data <= 10'h3fd; 
        10'b1010001101: data <= 10'h3fc; 
        10'b1010001110: data <= 10'h3fc; 
        10'b1010001111: data <= 10'h3fb; 
        10'b1010010000: data <= 10'h3fd; 
        10'b1010010001: data <= 10'h3fe; 
        10'b1010010010: data <= 10'h3fe; 
        10'b1010010011: data <= 10'h3fd; 
        10'b1010010100: data <= 10'h3fc; 
        10'b1010010101: data <= 10'h3fc; 
        10'b1010010110: data <= 10'h3fd; 
        10'b1010010111: data <= 10'h3ff; 
        10'b1010011000: data <= 10'h3ff; 
        10'b1010011001: data <= 10'h3ff; 
        10'b1010011010: data <= 10'h000; 
        10'b1010011011: data <= 10'h000; 
        10'b1010011100: data <= 10'h3ff; 
        10'b1010011101: data <= 10'h000; 
        10'b1010011110: data <= 10'h000; 
        10'b1010011111: data <= 10'h000; 
        10'b1010100000: data <= 10'h000; 
        10'b1010100001: data <= 10'h000; 
        10'b1010100010: data <= 10'h000; 
        10'b1010100011: data <= 10'h3ff; 
        10'b1010100100: data <= 10'h000; 
        10'b1010100101: data <= 10'h000; 
        10'b1010100110: data <= 10'h000; 
        10'b1010100111: data <= 10'h3ff; 
        10'b1010101000: data <= 10'h3ff; 
        10'b1010101001: data <= 10'h3ff; 
        10'b1010101010: data <= 10'h3ff; 
        10'b1010101011: data <= 10'h3fe; 
        10'b1010101100: data <= 10'h3fe; 
        10'b1010101101: data <= 10'h3fe; 
        10'b1010101110: data <= 10'h3fd; 
        10'b1010101111: data <= 10'h3fd; 
        10'b1010110000: data <= 10'h3fd; 
        10'b1010110001: data <= 10'h3fe; 
        10'b1010110010: data <= 10'h3ff; 
        10'b1010110011: data <= 10'h3ff; 
        10'b1010110100: data <= 10'h000; 
        10'b1010110101: data <= 10'h000; 
        10'b1010110110: data <= 10'h000; 
        10'b1010110111: data <= 10'h000; 
        10'b1010111000: data <= 10'h3ff; 
        10'b1010111001: data <= 10'h000; 
        10'b1010111010: data <= 10'h000; 
        10'b1010111011: data <= 10'h000; 
        10'b1010111100: data <= 10'h000; 
        10'b1010111101: data <= 10'h000; 
        10'b1010111110: data <= 10'h000; 
        10'b1010111111: data <= 10'h000; 
        10'b1011000000: data <= 10'h000; 
        10'b1011000001: data <= 10'h000; 
        10'b1011000010: data <= 10'h000; 
        10'b1011000011: data <= 10'h000; 
        10'b1011000100: data <= 10'h3ff; 
        10'b1011000101: data <= 10'h000; 
        10'b1011000110: data <= 10'h3ff; 
        10'b1011000111: data <= 10'h000; 
        10'b1011001000: data <= 10'h000; 
        10'b1011001001: data <= 10'h3ff; 
        10'b1011001010: data <= 10'h000; 
        10'b1011001011: data <= 10'h000; 
        10'b1011001100: data <= 10'h000; 
        10'b1011001101: data <= 10'h000; 
        10'b1011001110: data <= 10'h000; 
        10'b1011001111: data <= 10'h3ff; 
        10'b1011010000: data <= 10'h000; 
        10'b1011010001: data <= 10'h000; 
        10'b1011010010: data <= 10'h000; 
        10'b1011010011: data <= 10'h000; 
        10'b1011010100: data <= 10'h001; 
        10'b1011010101: data <= 10'h000; 
        10'b1011010110: data <= 10'h000; 
        10'b1011010111: data <= 10'h000; 
        10'b1011011000: data <= 10'h001; 
        10'b1011011001: data <= 10'h000; 
        10'b1011011010: data <= 10'h000; 
        10'b1011011011: data <= 10'h000; 
        10'b1011011100: data <= 10'h000; 
        10'b1011011101: data <= 10'h000; 
        10'b1011011110: data <= 10'h000; 
        10'b1011011111: data <= 10'h000; 
        10'b1011100000: data <= 10'h000; 
        10'b1011100001: data <= 10'h000; 
        10'b1011100010: data <= 10'h000; 
        10'b1011100011: data <= 10'h000; 
        10'b1011100100: data <= 10'h000; 
        10'b1011100101: data <= 10'h000; 
        10'b1011100110: data <= 10'h000; 
        10'b1011100111: data <= 10'h000; 
        10'b1011101000: data <= 10'h000; 
        10'b1011101001: data <= 10'h000; 
        10'b1011101010: data <= 10'h000; 
        10'b1011101011: data <= 10'h000; 
        10'b1011101100: data <= 10'h000; 
        10'b1011101101: data <= 10'h000; 
        10'b1011101110: data <= 10'h000; 
        10'b1011101111: data <= 10'h000; 
        10'b1011110000: data <= 10'h000; 
        10'b1011110001: data <= 10'h000; 
        10'b1011110010: data <= 10'h000; 
        10'b1011110011: data <= 10'h000; 
        10'b1011110100: data <= 10'h001; 
        10'b1011110101: data <= 10'h000; 
        10'b1011110110: data <= 10'h000; 
        10'b1011110111: data <= 10'h000; 
        10'b1011111000: data <= 10'h000; 
        10'b1011111001: data <= 10'h000; 
        10'b1011111010: data <= 10'h000; 
        10'b1011111011: data <= 10'h000; 
        10'b1011111100: data <= 10'h000; 
        10'b1011111101: data <= 10'h3ff; 
        10'b1011111110: data <= 10'h000; 
        10'b1011111111: data <= 10'h000; 
        10'b1100000000: data <= 10'h3ff; 
        10'b1100000001: data <= 10'h000; 
        10'b1100000010: data <= 10'h000; 
        10'b1100000011: data <= 10'h3ff; 
        10'b1100000100: data <= 10'h000; 
        10'b1100000101: data <= 10'h000; 
        10'b1100000110: data <= 10'h000; 
        10'b1100000111: data <= 10'h000; 
        10'b1100001000: data <= 10'h000; 
        10'b1100001001: data <= 10'h000; 
        10'b1100001010: data <= 10'h000; 
        10'b1100001011: data <= 10'h000; 
        10'b1100001100: data <= 10'h000; 
        10'b1100001101: data <= 10'h000; 
        10'b1100001110: data <= 10'h000; 
        10'b1100001111: data <= 10'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 5) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 11'h000; 
        10'b0000000001: data <= 11'h001; 
        10'b0000000010: data <= 11'h7ff; 
        10'b0000000011: data <= 11'h000; 
        10'b0000000100: data <= 11'h000; 
        10'b0000000101: data <= 11'h000; 
        10'b0000000110: data <= 11'h000; 
        10'b0000000111: data <= 11'h001; 
        10'b0000001000: data <= 11'h7ff; 
        10'b0000001001: data <= 11'h7ff; 
        10'b0000001010: data <= 11'h000; 
        10'b0000001011: data <= 11'h7ff; 
        10'b0000001100: data <= 11'h000; 
        10'b0000001101: data <= 11'h001; 
        10'b0000001110: data <= 11'h001; 
        10'b0000001111: data <= 11'h7ff; 
        10'b0000010000: data <= 11'h000; 
        10'b0000010001: data <= 11'h001; 
        10'b0000010010: data <= 11'h000; 
        10'b0000010011: data <= 11'h000; 
        10'b0000010100: data <= 11'h7ff; 
        10'b0000010101: data <= 11'h7ff; 
        10'b0000010110: data <= 11'h000; 
        10'b0000010111: data <= 11'h001; 
        10'b0000011000: data <= 11'h001; 
        10'b0000011001: data <= 11'h001; 
        10'b0000011010: data <= 11'h7ff; 
        10'b0000011011: data <= 11'h7ff; 
        10'b0000011100: data <= 11'h001; 
        10'b0000011101: data <= 11'h001; 
        10'b0000011110: data <= 11'h001; 
        10'b0000011111: data <= 11'h000; 
        10'b0000100000: data <= 11'h7ff; 
        10'b0000100001: data <= 11'h7ff; 
        10'b0000100010: data <= 11'h001; 
        10'b0000100011: data <= 11'h002; 
        10'b0000100100: data <= 11'h001; 
        10'b0000100101: data <= 11'h000; 
        10'b0000100110: data <= 11'h001; 
        10'b0000100111: data <= 11'h001; 
        10'b0000101000: data <= 11'h002; 
        10'b0000101001: data <= 11'h001; 
        10'b0000101010: data <= 11'h001; 
        10'b0000101011: data <= 11'h001; 
        10'b0000101100: data <= 11'h7ff; 
        10'b0000101101: data <= 11'h001; 
        10'b0000101110: data <= 11'h001; 
        10'b0000101111: data <= 11'h001; 
        10'b0000110000: data <= 11'h000; 
        10'b0000110001: data <= 11'h7ff; 
        10'b0000110010: data <= 11'h001; 
        10'b0000110011: data <= 11'h001; 
        10'b0000110100: data <= 11'h000; 
        10'b0000110101: data <= 11'h001; 
        10'b0000110110: data <= 11'h000; 
        10'b0000110111: data <= 11'h001; 
        10'b0000111000: data <= 11'h7ff; 
        10'b0000111001: data <= 11'h7ff; 
        10'b0000111010: data <= 11'h7ff; 
        10'b0000111011: data <= 11'h000; 
        10'b0000111100: data <= 11'h001; 
        10'b0000111101: data <= 11'h000; 
        10'b0000111110: data <= 11'h001; 
        10'b0000111111: data <= 11'h002; 
        10'b0001000000: data <= 11'h001; 
        10'b0001000001: data <= 11'h002; 
        10'b0001000010: data <= 11'h003; 
        10'b0001000011: data <= 11'h004; 
        10'b0001000100: data <= 11'h004; 
        10'b0001000101: data <= 11'h004; 
        10'b0001000110: data <= 11'h002; 
        10'b0001000111: data <= 11'h001; 
        10'b0001001000: data <= 11'h003; 
        10'b0001001001: data <= 11'h001; 
        10'b0001001010: data <= 11'h001; 
        10'b0001001011: data <= 11'h001; 
        10'b0001001100: data <= 11'h001; 
        10'b0001001101: data <= 11'h001; 
        10'b0001001110: data <= 11'h001; 
        10'b0001001111: data <= 11'h000; 
        10'b0001010000: data <= 11'h001; 
        10'b0001010001: data <= 11'h000; 
        10'b0001010010: data <= 11'h7ff; 
        10'b0001010011: data <= 11'h000; 
        10'b0001010100: data <= 11'h7ff; 
        10'b0001010101: data <= 11'h000; 
        10'b0001010110: data <= 11'h001; 
        10'b0001010111: data <= 11'h000; 
        10'b0001011000: data <= 11'h001; 
        10'b0001011001: data <= 11'h7ff; 
        10'b0001011010: data <= 11'h001; 
        10'b0001011011: data <= 11'h001; 
        10'b0001011100: data <= 11'h002; 
        10'b0001011101: data <= 11'h003; 
        10'b0001011110: data <= 11'h003; 
        10'b0001011111: data <= 11'h004; 
        10'b0001100000: data <= 11'h003; 
        10'b0001100001: data <= 11'h003; 
        10'b0001100010: data <= 11'h005; 
        10'b0001100011: data <= 11'h005; 
        10'b0001100100: data <= 11'h003; 
        10'b0001100101: data <= 11'h004; 
        10'b0001100110: data <= 11'h006; 
        10'b0001100111: data <= 11'h006; 
        10'b0001101000: data <= 11'h006; 
        10'b0001101001: data <= 11'h005; 
        10'b0001101010: data <= 11'h006; 
        10'b0001101011: data <= 11'h003; 
        10'b0001101100: data <= 11'h003; 
        10'b0001101101: data <= 11'h001; 
        10'b0001101110: data <= 11'h000; 
        10'b0001101111: data <= 11'h001; 
        10'b0001110000: data <= 11'h000; 
        10'b0001110001: data <= 11'h000; 
        10'b0001110010: data <= 11'h000; 
        10'b0001110011: data <= 11'h001; 
        10'b0001110100: data <= 11'h001; 
        10'b0001110101: data <= 11'h000; 
        10'b0001110110: data <= 11'h000; 
        10'b0001110111: data <= 11'h002; 
        10'b0001111000: data <= 11'h000; 
        10'b0001111001: data <= 11'h000; 
        10'b0001111010: data <= 11'h002; 
        10'b0001111011: data <= 11'h001; 
        10'b0001111100: data <= 11'h001; 
        10'b0001111101: data <= 11'h000; 
        10'b0001111110: data <= 11'h001; 
        10'b0001111111: data <= 11'h001; 
        10'b0010000000: data <= 11'h004; 
        10'b0010000001: data <= 11'h004; 
        10'b0010000010: data <= 11'h006; 
        10'b0010000011: data <= 11'h006; 
        10'b0010000100: data <= 11'h008; 
        10'b0010000101: data <= 11'h008; 
        10'b0010000110: data <= 11'h007; 
        10'b0010000111: data <= 11'h005; 
        10'b0010001000: data <= 11'h001; 
        10'b0010001001: data <= 11'h001; 
        10'b0010001010: data <= 11'h000; 
        10'b0010001011: data <= 11'h000; 
        10'b0010001100: data <= 11'h000; 
        10'b0010001101: data <= 11'h001; 
        10'b0010001110: data <= 11'h000; 
        10'b0010001111: data <= 11'h000; 
        10'b0010010000: data <= 11'h7ff; 
        10'b0010010001: data <= 11'h000; 
        10'b0010010010: data <= 11'h7ff; 
        10'b0010010011: data <= 11'h7ff; 
        10'b0010010100: data <= 11'h001; 
        10'b0010010101: data <= 11'h7ff; 
        10'b0010010110: data <= 11'h000; 
        10'b0010010111: data <= 11'h7fc; 
        10'b0010011000: data <= 11'h7fe; 
        10'b0010011001: data <= 11'h7fe; 
        10'b0010011010: data <= 11'h7ff; 
        10'b0010011011: data <= 11'h7fe; 
        10'b0010011100: data <= 11'h7fe; 
        10'b0010011101: data <= 11'h000; 
        10'b0010011110: data <= 11'h003; 
        10'b0010011111: data <= 11'h005; 
        10'b0010100000: data <= 11'h005; 
        10'b0010100001: data <= 11'h004; 
        10'b0010100010: data <= 11'h003; 
        10'b0010100011: data <= 11'h002; 
        10'b0010100100: data <= 11'h000; 
        10'b0010100101: data <= 11'h000; 
        10'b0010100110: data <= 11'h7ff; 
        10'b0010100111: data <= 11'h001; 
        10'b0010101000: data <= 11'h000; 
        10'b0010101001: data <= 11'h001; 
        10'b0010101010: data <= 11'h001; 
        10'b0010101011: data <= 11'h7ff; 
        10'b0010101100: data <= 11'h000; 
        10'b0010101101: data <= 11'h000; 
        10'b0010101110: data <= 11'h000; 
        10'b0010101111: data <= 11'h000; 
        10'b0010110000: data <= 11'h7fe; 
        10'b0010110001: data <= 11'h7fe; 
        10'b0010110010: data <= 11'h7fb; 
        10'b0010110011: data <= 11'h7f9; 
        10'b0010110100: data <= 11'h7fc; 
        10'b0010110101: data <= 11'h7f8; 
        10'b0010110110: data <= 11'h7fd; 
        10'b0010110111: data <= 11'h7fe; 
        10'b0010111000: data <= 11'h7fc; 
        10'b0010111001: data <= 11'h7fd; 
        10'b0010111010: data <= 11'h7ff; 
        10'b0010111011: data <= 11'h7fe; 
        10'b0010111100: data <= 11'h7fd; 
        10'b0010111101: data <= 11'h7fd; 
        10'b0010111110: data <= 11'h7fb; 
        10'b0010111111: data <= 11'h7fd; 
        10'b0011000000: data <= 11'h7fd; 
        10'b0011000001: data <= 11'h7fd; 
        10'b0011000010: data <= 11'h000; 
        10'b0011000011: data <= 11'h001; 
        10'b0011000100: data <= 11'h000; 
        10'b0011000101: data <= 11'h001; 
        10'b0011000110: data <= 11'h000; 
        10'b0011000111: data <= 11'h000; 
        10'b0011001000: data <= 11'h000; 
        10'b0011001001: data <= 11'h7ff; 
        10'b0011001010: data <= 11'h7fe; 
        10'b0011001011: data <= 11'h000; 
        10'b0011001100: data <= 11'h7fd; 
        10'b0011001101: data <= 11'h7fc; 
        10'b0011001110: data <= 11'h7fb; 
        10'b0011001111: data <= 11'h7fc; 
        10'b0011010000: data <= 11'h7f9; 
        10'b0011010001: data <= 11'h7f8; 
        10'b0011010010: data <= 11'h7fc; 
        10'b0011010011: data <= 11'h7fc; 
        10'b0011010100: data <= 11'h7fa; 
        10'b0011010101: data <= 11'h7fa; 
        10'b0011010110: data <= 11'h7f9; 
        10'b0011010111: data <= 11'h7f6; 
        10'b0011011000: data <= 11'h7f6; 
        10'b0011011001: data <= 11'h7f7; 
        10'b0011011010: data <= 11'h7f7; 
        10'b0011011011: data <= 11'h7f9; 
        10'b0011011100: data <= 11'h7fd; 
        10'b0011011101: data <= 11'h7fe; 
        10'b0011011110: data <= 11'h7ff; 
        10'b0011011111: data <= 11'h7ff; 
        10'b0011100000: data <= 11'h000; 
        10'b0011100001: data <= 11'h000; 
        10'b0011100010: data <= 11'h001; 
        10'b0011100011: data <= 11'h7ff; 
        10'b0011100100: data <= 11'h7ff; 
        10'b0011100101: data <= 11'h7fe; 
        10'b0011100110: data <= 11'h7fc; 
        10'b0011100111: data <= 11'h7ff; 
        10'b0011101000: data <= 11'h7ff; 
        10'b0011101001: data <= 11'h7fc; 
        10'b0011101010: data <= 11'h7fb; 
        10'b0011101011: data <= 11'h7fb; 
        10'b0011101100: data <= 11'h7f9; 
        10'b0011101101: data <= 11'h7f8; 
        10'b0011101110: data <= 11'h7f9; 
        10'b0011101111: data <= 11'h7f8; 
        10'b0011110000: data <= 11'h7f7; 
        10'b0011110001: data <= 11'h7f5; 
        10'b0011110010: data <= 11'h7f1; 
        10'b0011110011: data <= 11'h7f2; 
        10'b0011110100: data <= 11'h7f3; 
        10'b0011110101: data <= 11'h7f3; 
        10'b0011110110: data <= 11'h7f7; 
        10'b0011110111: data <= 11'h7f8; 
        10'b0011111000: data <= 11'h7fb; 
        10'b0011111001: data <= 11'h7fd; 
        10'b0011111010: data <= 11'h7fe; 
        10'b0011111011: data <= 11'h000; 
        10'b0011111100: data <= 11'h000; 
        10'b0011111101: data <= 11'h7ff; 
        10'b0011111110: data <= 11'h000; 
        10'b0011111111: data <= 11'h7ff; 
        10'b0100000000: data <= 11'h000; 
        10'b0100000001: data <= 11'h7ff; 
        10'b0100000010: data <= 11'h7ff; 
        10'b0100000011: data <= 11'h7ff; 
        10'b0100000100: data <= 11'h001; 
        10'b0100000101: data <= 11'h7fe; 
        10'b0100000110: data <= 11'h7fb; 
        10'b0100000111: data <= 11'h7fc; 
        10'b0100001000: data <= 11'h7fe; 
        10'b0100001001: data <= 11'h7fc; 
        10'b0100001010: data <= 11'h7fc; 
        10'b0100001011: data <= 11'h7f7; 
        10'b0100001100: data <= 11'h7f6; 
        10'b0100001101: data <= 11'h7f1; 
        10'b0100001110: data <= 11'h7f0; 
        10'b0100001111: data <= 11'h7f3; 
        10'b0100010000: data <= 11'h7f6; 
        10'b0100010001: data <= 11'h7f8; 
        10'b0100010010: data <= 11'h7f6; 
        10'b0100010011: data <= 11'h7fa; 
        10'b0100010100: data <= 11'h7fb; 
        10'b0100010101: data <= 11'h7fc; 
        10'b0100010110: data <= 11'h7ff; 
        10'b0100010111: data <= 11'h001; 
        10'b0100011000: data <= 11'h7ff; 
        10'b0100011001: data <= 11'h001; 
        10'b0100011010: data <= 11'h001; 
        10'b0100011011: data <= 11'h7ff; 
        10'b0100011100: data <= 11'h7fe; 
        10'b0100011101: data <= 11'h000; 
        10'b0100011110: data <= 11'h001; 
        10'b0100011111: data <= 11'h001; 
        10'b0100100000: data <= 11'h005; 
        10'b0100100001: data <= 11'h000; 
        10'b0100100010: data <= 11'h001; 
        10'b0100100011: data <= 11'h000; 
        10'b0100100100: data <= 11'h7fd; 
        10'b0100100101: data <= 11'h7fe; 
        10'b0100100110: data <= 11'h7fc; 
        10'b0100100111: data <= 11'h7f7; 
        10'b0100101000: data <= 11'h7f7; 
        10'b0100101001: data <= 11'h7f5; 
        10'b0100101010: data <= 11'h7f5; 
        10'b0100101011: data <= 11'h7f7; 
        10'b0100101100: data <= 11'h7fa; 
        10'b0100101101: data <= 11'h7fc; 
        10'b0100101110: data <= 11'h7fa; 
        10'b0100101111: data <= 11'h7ff; 
        10'b0100110000: data <= 11'h7fc; 
        10'b0100110001: data <= 11'h7fd; 
        10'b0100110010: data <= 11'h7ff; 
        10'b0100110011: data <= 11'h000; 
        10'b0100110100: data <= 11'h7ff; 
        10'b0100110101: data <= 11'h000; 
        10'b0100110110: data <= 11'h7ff; 
        10'b0100110111: data <= 11'h000; 
        10'b0100111000: data <= 11'h7ff; 
        10'b0100111001: data <= 11'h000; 
        10'b0100111010: data <= 11'h000; 
        10'b0100111011: data <= 11'h004; 
        10'b0100111100: data <= 11'h003; 
        10'b0100111101: data <= 11'h001; 
        10'b0100111110: data <= 11'h002; 
        10'b0100111111: data <= 11'h001; 
        10'b0101000000: data <= 11'h001; 
        10'b0101000001: data <= 11'h000; 
        10'b0101000010: data <= 11'h7fe; 
        10'b0101000011: data <= 11'h7f9; 
        10'b0101000100: data <= 11'h7f9; 
        10'b0101000101: data <= 11'h7fa; 
        10'b0101000110: data <= 11'h7fa; 
        10'b0101000111: data <= 11'h7fc; 
        10'b0101001000: data <= 11'h7fe; 
        10'b0101001001: data <= 11'h001; 
        10'b0101001010: data <= 11'h003; 
        10'b0101001011: data <= 11'h004; 
        10'b0101001100: data <= 11'h000; 
        10'b0101001101: data <= 11'h7fe; 
        10'b0101001110: data <= 11'h7ff; 
        10'b0101001111: data <= 11'h000; 
        10'b0101010000: data <= 11'h7ff; 
        10'b0101010001: data <= 11'h000; 
        10'b0101010010: data <= 11'h7ff; 
        10'b0101010011: data <= 11'h000; 
        10'b0101010100: data <= 11'h001; 
        10'b0101010101: data <= 11'h002; 
        10'b0101010110: data <= 11'h003; 
        10'b0101010111: data <= 11'h004; 
        10'b0101011000: data <= 11'h002; 
        10'b0101011001: data <= 11'h002; 
        10'b0101011010: data <= 11'h002; 
        10'b0101011011: data <= 11'h004; 
        10'b0101011100: data <= 11'h004; 
        10'b0101011101: data <= 11'h003; 
        10'b0101011110: data <= 11'h7fd; 
        10'b0101011111: data <= 11'h7fb; 
        10'b0101100000: data <= 11'h000; 
        10'b0101100001: data <= 11'h000; 
        10'b0101100010: data <= 11'h7fb; 
        10'b0101100011: data <= 11'h7fc; 
        10'b0101100100: data <= 11'h7ff; 
        10'b0101100101: data <= 11'h003; 
        10'b0101100110: data <= 11'h006; 
        10'b0101100111: data <= 11'h00b; 
        10'b0101101000: data <= 11'h006; 
        10'b0101101001: data <= 11'h7fe; 
        10'b0101101010: data <= 11'h7fe; 
        10'b0101101011: data <= 11'h7ff; 
        10'b0101101100: data <= 11'h7ff; 
        10'b0101101101: data <= 11'h001; 
        10'b0101101110: data <= 11'h001; 
        10'b0101101111: data <= 11'h7ff; 
        10'b0101110000: data <= 11'h7fe; 
        10'b0101110001: data <= 11'h001; 
        10'b0101110010: data <= 11'h005; 
        10'b0101110011: data <= 11'h003; 
        10'b0101110100: data <= 11'h002; 
        10'b0101110101: data <= 11'h001; 
        10'b0101110110: data <= 11'h005; 
        10'b0101110111: data <= 11'h004; 
        10'b0101111000: data <= 11'h004; 
        10'b0101111001: data <= 11'h001; 
        10'b0101111010: data <= 11'h7ff; 
        10'b0101111011: data <= 11'h000; 
        10'b0101111100: data <= 11'h000; 
        10'b0101111101: data <= 11'h7ff; 
        10'b0101111110: data <= 11'h7fc; 
        10'b0101111111: data <= 11'h7ff; 
        10'b0110000000: data <= 11'h7fe; 
        10'b0110000001: data <= 11'h003; 
        10'b0110000010: data <= 11'h008; 
        10'b0110000011: data <= 11'h00d; 
        10'b0110000100: data <= 11'h007; 
        10'b0110000101: data <= 11'h7ff; 
        10'b0110000110: data <= 11'h000; 
        10'b0110000111: data <= 11'h001; 
        10'b0110001000: data <= 11'h000; 
        10'b0110001001: data <= 11'h000; 
        10'b0110001010: data <= 11'h001; 
        10'b0110001011: data <= 11'h000; 
        10'b0110001100: data <= 11'h7fe; 
        10'b0110001101: data <= 11'h002; 
        10'b0110001110: data <= 11'h004; 
        10'b0110001111: data <= 11'h004; 
        10'b0110010000: data <= 11'h005; 
        10'b0110010001: data <= 11'h005; 
        10'b0110010010: data <= 11'h005; 
        10'b0110010011: data <= 11'h006; 
        10'b0110010100: data <= 11'h002; 
        10'b0110010101: data <= 11'h7fd; 
        10'b0110010110: data <= 11'h000; 
        10'b0110010111: data <= 11'h002; 
        10'b0110011000: data <= 11'h001; 
        10'b0110011001: data <= 11'h7fe; 
        10'b0110011010: data <= 11'h7fe; 
        10'b0110011011: data <= 11'h000; 
        10'b0110011100: data <= 11'h004; 
        10'b0110011101: data <= 11'h004; 
        10'b0110011110: data <= 11'h00a; 
        10'b0110011111: data <= 11'h00b; 
        10'b0110100000: data <= 11'h007; 
        10'b0110100001: data <= 11'h000; 
        10'b0110100010: data <= 11'h7fe; 
        10'b0110100011: data <= 11'h7ff; 
        10'b0110100100: data <= 11'h001; 
        10'b0110100101: data <= 11'h000; 
        10'b0110100110: data <= 11'h000; 
        10'b0110100111: data <= 11'h7ff; 
        10'b0110101000: data <= 11'h7fd; 
        10'b0110101001: data <= 11'h000; 
        10'b0110101010: data <= 11'h005; 
        10'b0110101011: data <= 11'h006; 
        10'b0110101100: data <= 11'h004; 
        10'b0110101101: data <= 11'h006; 
        10'b0110101110: data <= 11'h008; 
        10'b0110101111: data <= 11'h009; 
        10'b0110110000: data <= 11'h002; 
        10'b0110110001: data <= 11'h7ff; 
        10'b0110110010: data <= 11'h004; 
        10'b0110110011: data <= 11'h003; 
        10'b0110110100: data <= 11'h001; 
        10'b0110110101: data <= 11'h7fe; 
        10'b0110110110: data <= 11'h000; 
        10'b0110110111: data <= 11'h002; 
        10'b0110111000: data <= 11'h004; 
        10'b0110111001: data <= 11'h006; 
        10'b0110111010: data <= 11'h005; 
        10'b0110111011: data <= 11'h007; 
        10'b0110111100: data <= 11'h004; 
        10'b0110111101: data <= 11'h7fe; 
        10'b0110111110: data <= 11'h7ff; 
        10'b0110111111: data <= 11'h7ff; 
        10'b0111000000: data <= 11'h000; 
        10'b0111000001: data <= 11'h7ff; 
        10'b0111000010: data <= 11'h7ff; 
        10'b0111000011: data <= 11'h7ff; 
        10'b0111000100: data <= 11'h7fc; 
        10'b0111000101: data <= 11'h7fe; 
        10'b0111000110: data <= 11'h007; 
        10'b0111000111: data <= 11'h007; 
        10'b0111001000: data <= 11'h005; 
        10'b0111001001: data <= 11'h007; 
        10'b0111001010: data <= 11'h00c; 
        10'b0111001011: data <= 11'h00c; 
        10'b0111001100: data <= 11'h004; 
        10'b0111001101: data <= 11'h002; 
        10'b0111001110: data <= 11'h005; 
        10'b0111001111: data <= 11'h003; 
        10'b0111010000: data <= 11'h7ff; 
        10'b0111010001: data <= 11'h7fd; 
        10'b0111010010: data <= 11'h001; 
        10'b0111010011: data <= 11'h003; 
        10'b0111010100: data <= 11'h001; 
        10'b0111010101: data <= 11'h000; 
        10'b0111010110: data <= 11'h003; 
        10'b0111010111: data <= 11'h002; 
        10'b0111011000: data <= 11'h7ff; 
        10'b0111011001: data <= 11'h7fe; 
        10'b0111011010: data <= 11'h7ff; 
        10'b0111011011: data <= 11'h000; 
        10'b0111011100: data <= 11'h000; 
        10'b0111011101: data <= 11'h001; 
        10'b0111011110: data <= 11'h001; 
        10'b0111011111: data <= 11'h000; 
        10'b0111100000: data <= 11'h7fa; 
        10'b0111100001: data <= 11'h7fd; 
        10'b0111100010: data <= 11'h003; 
        10'b0111100011: data <= 11'h005; 
        10'b0111100100: data <= 11'h006; 
        10'b0111100101: data <= 11'h008; 
        10'b0111100110: data <= 11'h00d; 
        10'b0111100111: data <= 11'h00d; 
        10'b0111101000: data <= 11'h007; 
        10'b0111101001: data <= 11'h004; 
        10'b0111101010: data <= 11'h004; 
        10'b0111101011: data <= 11'h002; 
        10'b0111101100: data <= 11'h000; 
        10'b0111101101: data <= 11'h001; 
        10'b0111101110: data <= 11'h005; 
        10'b0111101111: data <= 11'h002; 
        10'b0111110000: data <= 11'h001; 
        10'b0111110001: data <= 11'h7ff; 
        10'b0111110010: data <= 11'h001; 
        10'b0111110011: data <= 11'h000; 
        10'b0111110100: data <= 11'h7fe; 
        10'b0111110101: data <= 11'h7fd; 
        10'b0111110110: data <= 11'h000; 
        10'b0111110111: data <= 11'h000; 
        10'b0111111000: data <= 11'h000; 
        10'b0111111001: data <= 11'h7ff; 
        10'b0111111010: data <= 11'h000; 
        10'b0111111011: data <= 11'h7fe; 
        10'b0111111100: data <= 11'h7fb; 
        10'b0111111101: data <= 11'h7fb; 
        10'b0111111110: data <= 11'h7fd; 
        10'b0111111111: data <= 11'h004; 
        10'b1000000000: data <= 11'h006; 
        10'b1000000001: data <= 11'h005; 
        10'b1000000010: data <= 11'h009; 
        10'b1000000011: data <= 11'h00b; 
        10'b1000000100: data <= 11'h00d; 
        10'b1000000101: data <= 11'h006; 
        10'b1000000110: data <= 11'h002; 
        10'b1000000111: data <= 11'h003; 
        10'b1000001000: data <= 11'h006; 
        10'b1000001001: data <= 11'h004; 
        10'b1000001010: data <= 11'h005; 
        10'b1000001011: data <= 11'h003; 
        10'b1000001100: data <= 11'h000; 
        10'b1000001101: data <= 11'h001; 
        10'b1000001110: data <= 11'h001; 
        10'b1000001111: data <= 11'h7ff; 
        10'b1000010000: data <= 11'h7fe; 
        10'b1000010001: data <= 11'h7ff; 
        10'b1000010010: data <= 11'h7ff; 
        10'b1000010011: data <= 11'h7ff; 
        10'b1000010100: data <= 11'h000; 
        10'b1000010101: data <= 11'h7ff; 
        10'b1000010110: data <= 11'h001; 
        10'b1000010111: data <= 11'h7fe; 
        10'b1000011000: data <= 11'h7fd; 
        10'b1000011001: data <= 11'h7fa; 
        10'b1000011010: data <= 11'h7fc; 
        10'b1000011011: data <= 11'h000; 
        10'b1000011100: data <= 11'h004; 
        10'b1000011101: data <= 11'h006; 
        10'b1000011110: data <= 11'h008; 
        10'b1000011111: data <= 11'h00d; 
        10'b1000100000: data <= 11'h00e; 
        10'b1000100001: data <= 11'h007; 
        10'b1000100010: data <= 11'h007; 
        10'b1000100011: data <= 11'h007; 
        10'b1000100100: data <= 11'h005; 
        10'b1000100101: data <= 11'h004; 
        10'b1000100110: data <= 11'h006; 
        10'b1000100111: data <= 11'h004; 
        10'b1000101000: data <= 11'h003; 
        10'b1000101001: data <= 11'h001; 
        10'b1000101010: data <= 11'h7ff; 
        10'b1000101011: data <= 11'h7ff; 
        10'b1000101100: data <= 11'h7ff; 
        10'b1000101101: data <= 11'h000; 
        10'b1000101110: data <= 11'h7ff; 
        10'b1000101111: data <= 11'h001; 
        10'b1000110000: data <= 11'h7ff; 
        10'b1000110001: data <= 11'h7ff; 
        10'b1000110010: data <= 11'h000; 
        10'b1000110011: data <= 11'h7ff; 
        10'b1000110100: data <= 11'h7fc; 
        10'b1000110101: data <= 11'h7fb; 
        10'b1000110110: data <= 11'h7fb; 
        10'b1000110111: data <= 11'h7fe; 
        10'b1000111000: data <= 11'h001; 
        10'b1000111001: data <= 11'h004; 
        10'b1000111010: data <= 11'h007; 
        10'b1000111011: data <= 11'h004; 
        10'b1000111100: data <= 11'h009; 
        10'b1000111101: data <= 11'h00a; 
        10'b1000111110: data <= 11'h00c; 
        10'b1000111111: data <= 11'h00a; 
        10'b1001000000: data <= 11'h006; 
        10'b1001000001: data <= 11'h004; 
        10'b1001000010: data <= 11'h007; 
        10'b1001000011: data <= 11'h005; 
        10'b1001000100: data <= 11'h003; 
        10'b1001000101: data <= 11'h7ff; 
        10'b1001000110: data <= 11'h7fd; 
        10'b1001000111: data <= 11'h000; 
        10'b1001001000: data <= 11'h7ff; 
        10'b1001001001: data <= 11'h000; 
        10'b1001001010: data <= 11'h7ff; 
        10'b1001001011: data <= 11'h000; 
        10'b1001001100: data <= 11'h000; 
        10'b1001001101: data <= 11'h000; 
        10'b1001001110: data <= 11'h000; 
        10'b1001001111: data <= 11'h000; 
        10'b1001010000: data <= 11'h7fe; 
        10'b1001010001: data <= 11'h7fc; 
        10'b1001010010: data <= 11'h7fa; 
        10'b1001010011: data <= 11'h7fd; 
        10'b1001010100: data <= 11'h7fe; 
        10'b1001010101: data <= 11'h003; 
        10'b1001010110: data <= 11'h005; 
        10'b1001010111: data <= 11'h008; 
        10'b1001011000: data <= 11'h00a; 
        10'b1001011001: data <= 11'h00a; 
        10'b1001011010: data <= 11'h009; 
        10'b1001011011: data <= 11'h007; 
        10'b1001011100: data <= 11'h005; 
        10'b1001011101: data <= 11'h006; 
        10'b1001011110: data <= 11'h006; 
        10'b1001011111: data <= 11'h004; 
        10'b1001100000: data <= 11'h000; 
        10'b1001100001: data <= 11'h7fe; 
        10'b1001100010: data <= 11'h7fd; 
        10'b1001100011: data <= 11'h7fe; 
        10'b1001100100: data <= 11'h000; 
        10'b1001100101: data <= 11'h7ff; 
        10'b1001100110: data <= 11'h000; 
        10'b1001100111: data <= 11'h7ff; 
        10'b1001101000: data <= 11'h7ff; 
        10'b1001101001: data <= 11'h000; 
        10'b1001101010: data <= 11'h001; 
        10'b1001101011: data <= 11'h000; 
        10'b1001101100: data <= 11'h7ff; 
        10'b1001101101: data <= 11'h7fd; 
        10'b1001101110: data <= 11'h7fc; 
        10'b1001101111: data <= 11'h7fb; 
        10'b1001110000: data <= 11'h7fd; 
        10'b1001110001: data <= 11'h7fe; 
        10'b1001110010: data <= 11'h7ff; 
        10'b1001110011: data <= 11'h001; 
        10'b1001110100: data <= 11'h003; 
        10'b1001110101: data <= 11'h001; 
        10'b1001110110: data <= 11'h001; 
        10'b1001110111: data <= 11'h003; 
        10'b1001111000: data <= 11'h002; 
        10'b1001111001: data <= 11'h000; 
        10'b1001111010: data <= 11'h7ff; 
        10'b1001111011: data <= 11'h7fc; 
        10'b1001111100: data <= 11'h7fd; 
        10'b1001111101: data <= 11'h7fd; 
        10'b1001111110: data <= 11'h7fd; 
        10'b1001111111: data <= 11'h000; 
        10'b1010000000: data <= 11'h000; 
        10'b1010000001: data <= 11'h7ff; 
        10'b1010000010: data <= 11'h001; 
        10'b1010000011: data <= 11'h000; 
        10'b1010000100: data <= 11'h001; 
        10'b1010000101: data <= 11'h000; 
        10'b1010000110: data <= 11'h000; 
        10'b1010000111: data <= 11'h000; 
        10'b1010001000: data <= 11'h000; 
        10'b1010001001: data <= 11'h7ff; 
        10'b1010001010: data <= 11'h7fe; 
        10'b1010001011: data <= 11'h7fb; 
        10'b1010001100: data <= 11'h7fa; 
        10'b1010001101: data <= 11'h7f8; 
        10'b1010001110: data <= 11'h7f8; 
        10'b1010001111: data <= 11'h7f6; 
        10'b1010010000: data <= 11'h7fa; 
        10'b1010010001: data <= 11'h7fb; 
        10'b1010010010: data <= 11'h7fc; 
        10'b1010010011: data <= 11'h7fb; 
        10'b1010010100: data <= 11'h7f9; 
        10'b1010010101: data <= 11'h7f8; 
        10'b1010010110: data <= 11'h7fa; 
        10'b1010010111: data <= 11'h7fd; 
        10'b1010011000: data <= 11'h7fd; 
        10'b1010011001: data <= 11'h7fd; 
        10'b1010011010: data <= 11'h7ff; 
        10'b1010011011: data <= 11'h000; 
        10'b1010011100: data <= 11'h7ff; 
        10'b1010011101: data <= 11'h7ff; 
        10'b1010011110: data <= 11'h000; 
        10'b1010011111: data <= 11'h000; 
        10'b1010100000: data <= 11'h001; 
        10'b1010100001: data <= 11'h000; 
        10'b1010100010: data <= 11'h000; 
        10'b1010100011: data <= 11'h7ff; 
        10'b1010100100: data <= 11'h7ff; 
        10'b1010100101: data <= 11'h000; 
        10'b1010100110: data <= 11'h7ff; 
        10'b1010100111: data <= 11'h7fe; 
        10'b1010101000: data <= 11'h7ff; 
        10'b1010101001: data <= 11'h7fe; 
        10'b1010101010: data <= 11'h7fd; 
        10'b1010101011: data <= 11'h7fc; 
        10'b1010101100: data <= 11'h7fc; 
        10'b1010101101: data <= 11'h7fc; 
        10'b1010101110: data <= 11'h7fb; 
        10'b1010101111: data <= 11'h7fb; 
        10'b1010110000: data <= 11'h7fb; 
        10'b1010110001: data <= 11'h7fc; 
        10'b1010110010: data <= 11'h7ff; 
        10'b1010110011: data <= 11'h7ff; 
        10'b1010110100: data <= 11'h000; 
        10'b1010110101: data <= 11'h7ff; 
        10'b1010110110: data <= 11'h001; 
        10'b1010110111: data <= 11'h000; 
        10'b1010111000: data <= 11'h7ff; 
        10'b1010111001: data <= 11'h000; 
        10'b1010111010: data <= 11'h7ff; 
        10'b1010111011: data <= 11'h7ff; 
        10'b1010111100: data <= 11'h001; 
        10'b1010111101: data <= 11'h7ff; 
        10'b1010111110: data <= 11'h000; 
        10'b1010111111: data <= 11'h000; 
        10'b1011000000: data <= 11'h7ff; 
        10'b1011000001: data <= 11'h000; 
        10'b1011000010: data <= 11'h001; 
        10'b1011000011: data <= 11'h000; 
        10'b1011000100: data <= 11'h7ff; 
        10'b1011000101: data <= 11'h000; 
        10'b1011000110: data <= 11'h7ff; 
        10'b1011000111: data <= 11'h000; 
        10'b1011001000: data <= 11'h000; 
        10'b1011001001: data <= 11'h7ff; 
        10'b1011001010: data <= 11'h7ff; 
        10'b1011001011: data <= 11'h000; 
        10'b1011001100: data <= 11'h000; 
        10'b1011001101: data <= 11'h7ff; 
        10'b1011001110: data <= 11'h7ff; 
        10'b1011001111: data <= 11'h7ff; 
        10'b1011010000: data <= 11'h7ff; 
        10'b1011010001: data <= 11'h000; 
        10'b1011010010: data <= 11'h000; 
        10'b1011010011: data <= 11'h001; 
        10'b1011010100: data <= 11'h001; 
        10'b1011010101: data <= 11'h001; 
        10'b1011010110: data <= 11'h000; 
        10'b1011010111: data <= 11'h001; 
        10'b1011011000: data <= 11'h001; 
        10'b1011011001: data <= 11'h000; 
        10'b1011011010: data <= 11'h000; 
        10'b1011011011: data <= 11'h000; 
        10'b1011011100: data <= 11'h7ff; 
        10'b1011011101: data <= 11'h001; 
        10'b1011011110: data <= 11'h001; 
        10'b1011011111: data <= 11'h7ff; 
        10'b1011100000: data <= 11'h000; 
        10'b1011100001: data <= 11'h001; 
        10'b1011100010: data <= 11'h000; 
        10'b1011100011: data <= 11'h000; 
        10'b1011100100: data <= 11'h000; 
        10'b1011100101: data <= 11'h001; 
        10'b1011100110: data <= 11'h001; 
        10'b1011100111: data <= 11'h7ff; 
        10'b1011101000: data <= 11'h7ff; 
        10'b1011101001: data <= 11'h001; 
        10'b1011101010: data <= 11'h001; 
        10'b1011101011: data <= 11'h000; 
        10'b1011101100: data <= 11'h001; 
        10'b1011101101: data <= 11'h000; 
        10'b1011101110: data <= 11'h000; 
        10'b1011101111: data <= 11'h000; 
        10'b1011110000: data <= 11'h000; 
        10'b1011110001: data <= 11'h000; 
        10'b1011110010: data <= 11'h7ff; 
        10'b1011110011: data <= 11'h000; 
        10'b1011110100: data <= 11'h001; 
        10'b1011110101: data <= 11'h000; 
        10'b1011110110: data <= 11'h001; 
        10'b1011110111: data <= 11'h7ff; 
        10'b1011111000: data <= 11'h000; 
        10'b1011111001: data <= 11'h000; 
        10'b1011111010: data <= 11'h001; 
        10'b1011111011: data <= 11'h000; 
        10'b1011111100: data <= 11'h000; 
        10'b1011111101: data <= 11'h7ff; 
        10'b1011111110: data <= 11'h7ff; 
        10'b1011111111: data <= 11'h000; 
        10'b1100000000: data <= 11'h7ff; 
        10'b1100000001: data <= 11'h7ff; 
        10'b1100000010: data <= 11'h7ff; 
        10'b1100000011: data <= 11'h7ff; 
        10'b1100000100: data <= 11'h7ff; 
        10'b1100000101: data <= 11'h000; 
        10'b1100000110: data <= 11'h7ff; 
        10'b1100000111: data <= 11'h7ff; 
        10'b1100001000: data <= 11'h7ff; 
        10'b1100001001: data <= 11'h000; 
        10'b1100001010: data <= 11'h001; 
        10'b1100001011: data <= 11'h7ff; 
        10'b1100001100: data <= 11'h7ff; 
        10'b1100001101: data <= 11'h7ff; 
        10'b1100001110: data <= 11'h7ff; 
        10'b1100001111: data <= 11'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 6) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 12'hfff; 
        10'b0000000001: data <= 12'h001; 
        10'b0000000010: data <= 12'hffe; 
        10'b0000000011: data <= 12'h000; 
        10'b0000000100: data <= 12'h000; 
        10'b0000000101: data <= 12'h000; 
        10'b0000000110: data <= 12'h001; 
        10'b0000000111: data <= 12'h002; 
        10'b0000001000: data <= 12'hffe; 
        10'b0000001001: data <= 12'hfff; 
        10'b0000001010: data <= 12'hfff; 
        10'b0000001011: data <= 12'hfff; 
        10'b0000001100: data <= 12'h001; 
        10'b0000001101: data <= 12'h002; 
        10'b0000001110: data <= 12'h001; 
        10'b0000001111: data <= 12'hffe; 
        10'b0000010000: data <= 12'h000; 
        10'b0000010001: data <= 12'h002; 
        10'b0000010010: data <= 12'h000; 
        10'b0000010011: data <= 12'h000; 
        10'b0000010100: data <= 12'hffe; 
        10'b0000010101: data <= 12'hfff; 
        10'b0000010110: data <= 12'h001; 
        10'b0000010111: data <= 12'h002; 
        10'b0000011000: data <= 12'h001; 
        10'b0000011001: data <= 12'h001; 
        10'b0000011010: data <= 12'hffe; 
        10'b0000011011: data <= 12'hffe; 
        10'b0000011100: data <= 12'h001; 
        10'b0000011101: data <= 12'h001; 
        10'b0000011110: data <= 12'h001; 
        10'b0000011111: data <= 12'h000; 
        10'b0000100000: data <= 12'hffe; 
        10'b0000100001: data <= 12'hfff; 
        10'b0000100010: data <= 12'h001; 
        10'b0000100011: data <= 12'h003; 
        10'b0000100100: data <= 12'h002; 
        10'b0000100101: data <= 12'h001; 
        10'b0000100110: data <= 12'h003; 
        10'b0000100111: data <= 12'h003; 
        10'b0000101000: data <= 12'h003; 
        10'b0000101001: data <= 12'h003; 
        10'b0000101010: data <= 12'h002; 
        10'b0000101011: data <= 12'h002; 
        10'b0000101100: data <= 12'hffe; 
        10'b0000101101: data <= 12'h002; 
        10'b0000101110: data <= 12'h003; 
        10'b0000101111: data <= 12'h001; 
        10'b0000110000: data <= 12'h000; 
        10'b0000110001: data <= 12'hfff; 
        10'b0000110010: data <= 12'h003; 
        10'b0000110011: data <= 12'h002; 
        10'b0000110100: data <= 12'hfff; 
        10'b0000110101: data <= 12'h002; 
        10'b0000110110: data <= 12'h000; 
        10'b0000110111: data <= 12'h002; 
        10'b0000111000: data <= 12'hfff; 
        10'b0000111001: data <= 12'hffe; 
        10'b0000111010: data <= 12'hffe; 
        10'b0000111011: data <= 12'h000; 
        10'b0000111100: data <= 12'h001; 
        10'b0000111101: data <= 12'h001; 
        10'b0000111110: data <= 12'h001; 
        10'b0000111111: data <= 12'h003; 
        10'b0001000000: data <= 12'h002; 
        10'b0001000001: data <= 12'h005; 
        10'b0001000010: data <= 12'h006; 
        10'b0001000011: data <= 12'h007; 
        10'b0001000100: data <= 12'h007; 
        10'b0001000101: data <= 12'h007; 
        10'b0001000110: data <= 12'h004; 
        10'b0001000111: data <= 12'h003; 
        10'b0001001000: data <= 12'h006; 
        10'b0001001001: data <= 12'h003; 
        10'b0001001010: data <= 12'h003; 
        10'b0001001011: data <= 12'h003; 
        10'b0001001100: data <= 12'h003; 
        10'b0001001101: data <= 12'h001; 
        10'b0001001110: data <= 12'h002; 
        10'b0001001111: data <= 12'h000; 
        10'b0001010000: data <= 12'h001; 
        10'b0001010001: data <= 12'hfff; 
        10'b0001010010: data <= 12'hffe; 
        10'b0001010011: data <= 12'h001; 
        10'b0001010100: data <= 12'hffe; 
        10'b0001010101: data <= 12'h000; 
        10'b0001010110: data <= 12'h002; 
        10'b0001010111: data <= 12'h001; 
        10'b0001011000: data <= 12'h002; 
        10'b0001011001: data <= 12'hffe; 
        10'b0001011010: data <= 12'h002; 
        10'b0001011011: data <= 12'h003; 
        10'b0001011100: data <= 12'h003; 
        10'b0001011101: data <= 12'h006; 
        10'b0001011110: data <= 12'h006; 
        10'b0001011111: data <= 12'h007; 
        10'b0001100000: data <= 12'h007; 
        10'b0001100001: data <= 12'h007; 
        10'b0001100010: data <= 12'h00a; 
        10'b0001100011: data <= 12'h009; 
        10'b0001100100: data <= 12'h006; 
        10'b0001100101: data <= 12'h007; 
        10'b0001100110: data <= 12'h00c; 
        10'b0001100111: data <= 12'h00c; 
        10'b0001101000: data <= 12'h00c; 
        10'b0001101001: data <= 12'h00b; 
        10'b0001101010: data <= 12'h00b; 
        10'b0001101011: data <= 12'h006; 
        10'b0001101100: data <= 12'h006; 
        10'b0001101101: data <= 12'h001; 
        10'b0001101110: data <= 12'hfff; 
        10'b0001101111: data <= 12'h001; 
        10'b0001110000: data <= 12'h000; 
        10'b0001110001: data <= 12'h000; 
        10'b0001110010: data <= 12'h000; 
        10'b0001110011: data <= 12'h002; 
        10'b0001110100: data <= 12'h002; 
        10'b0001110101: data <= 12'h001; 
        10'b0001110110: data <= 12'h001; 
        10'b0001110111: data <= 12'h004; 
        10'b0001111000: data <= 12'h000; 
        10'b0001111001: data <= 12'hfff; 
        10'b0001111010: data <= 12'h004; 
        10'b0001111011: data <= 12'h001; 
        10'b0001111100: data <= 12'h002; 
        10'b0001111101: data <= 12'h001; 
        10'b0001111110: data <= 12'h001; 
        10'b0001111111: data <= 12'h002; 
        10'b0010000000: data <= 12'h008; 
        10'b0010000001: data <= 12'h008; 
        10'b0010000010: data <= 12'h00c; 
        10'b0010000011: data <= 12'h00c; 
        10'b0010000100: data <= 12'h00f; 
        10'b0010000101: data <= 12'h011; 
        10'b0010000110: data <= 12'h00f; 
        10'b0010000111: data <= 12'h00a; 
        10'b0010001000: data <= 12'h001; 
        10'b0010001001: data <= 12'h003; 
        10'b0010001010: data <= 12'h000; 
        10'b0010001011: data <= 12'h000; 
        10'b0010001100: data <= 12'h000; 
        10'b0010001101: data <= 12'h001; 
        10'b0010001110: data <= 12'h001; 
        10'b0010001111: data <= 12'hfff; 
        10'b0010010000: data <= 12'hffe; 
        10'b0010010001: data <= 12'h000; 
        10'b0010010010: data <= 12'hfff; 
        10'b0010010011: data <= 12'hffd; 
        10'b0010010100: data <= 12'h002; 
        10'b0010010101: data <= 12'hffd; 
        10'b0010010110: data <= 12'h001; 
        10'b0010010111: data <= 12'hff7; 
        10'b0010011000: data <= 12'hffb; 
        10'b0010011001: data <= 12'hffd; 
        10'b0010011010: data <= 12'hfff; 
        10'b0010011011: data <= 12'hffc; 
        10'b0010011100: data <= 12'hffc; 
        10'b0010011101: data <= 12'h001; 
        10'b0010011110: data <= 12'h006; 
        10'b0010011111: data <= 12'h00b; 
        10'b0010100000: data <= 12'h009; 
        10'b0010100001: data <= 12'h008; 
        10'b0010100010: data <= 12'h007; 
        10'b0010100011: data <= 12'h005; 
        10'b0010100100: data <= 12'hfff; 
        10'b0010100101: data <= 12'h000; 
        10'b0010100110: data <= 12'hffe; 
        10'b0010100111: data <= 12'h002; 
        10'b0010101000: data <= 12'h000; 
        10'b0010101001: data <= 12'h002; 
        10'b0010101010: data <= 12'h002; 
        10'b0010101011: data <= 12'hffe; 
        10'b0010101100: data <= 12'h001; 
        10'b0010101101: data <= 12'h000; 
        10'b0010101110: data <= 12'h001; 
        10'b0010101111: data <= 12'h000; 
        10'b0010110000: data <= 12'hffd; 
        10'b0010110001: data <= 12'hffc; 
        10'b0010110010: data <= 12'hff6; 
        10'b0010110011: data <= 12'hff3; 
        10'b0010110100: data <= 12'hff8; 
        10'b0010110101: data <= 12'hff1; 
        10'b0010110110: data <= 12'hff9; 
        10'b0010110111: data <= 12'hffb; 
        10'b0010111000: data <= 12'hff9; 
        10'b0010111001: data <= 12'hffa; 
        10'b0010111010: data <= 12'hffe; 
        10'b0010111011: data <= 12'hffc; 
        10'b0010111100: data <= 12'hff9; 
        10'b0010111101: data <= 12'hffa; 
        10'b0010111110: data <= 12'hff6; 
        10'b0010111111: data <= 12'hff9; 
        10'b0011000000: data <= 12'hffb; 
        10'b0011000001: data <= 12'hffa; 
        10'b0011000010: data <= 12'hfff; 
        10'b0011000011: data <= 12'h002; 
        10'b0011000100: data <= 12'h001; 
        10'b0011000101: data <= 12'h001; 
        10'b0011000110: data <= 12'h000; 
        10'b0011000111: data <= 12'h000; 
        10'b0011001000: data <= 12'h000; 
        10'b0011001001: data <= 12'hffe; 
        10'b0011001010: data <= 12'hffc; 
        10'b0011001011: data <= 12'hfff; 
        10'b0011001100: data <= 12'hffa; 
        10'b0011001101: data <= 12'hff9; 
        10'b0011001110: data <= 12'hff6; 
        10'b0011001111: data <= 12'hff8; 
        10'b0011010000: data <= 12'hff1; 
        10'b0011010001: data <= 12'hff0; 
        10'b0011010010: data <= 12'hff7; 
        10'b0011010011: data <= 12'hff8; 
        10'b0011010100: data <= 12'hff3; 
        10'b0011010101: data <= 12'hff4; 
        10'b0011010110: data <= 12'hff1; 
        10'b0011010111: data <= 12'hfec; 
        10'b0011011000: data <= 12'hfeb; 
        10'b0011011001: data <= 12'hfef; 
        10'b0011011010: data <= 12'hfee; 
        10'b0011011011: data <= 12'hff2; 
        10'b0011011100: data <= 12'hffb; 
        10'b0011011101: data <= 12'hffb; 
        10'b0011011110: data <= 12'hffe; 
        10'b0011011111: data <= 12'hfff; 
        10'b0011100000: data <= 12'hfff; 
        10'b0011100001: data <= 12'hfff; 
        10'b0011100010: data <= 12'h002; 
        10'b0011100011: data <= 12'hffd; 
        10'b0011100100: data <= 12'hffe; 
        10'b0011100101: data <= 12'hffd; 
        10'b0011100110: data <= 12'hff8; 
        10'b0011100111: data <= 12'hffe; 
        10'b0011101000: data <= 12'hffd; 
        10'b0011101001: data <= 12'hff8; 
        10'b0011101010: data <= 12'hff6; 
        10'b0011101011: data <= 12'hff5; 
        10'b0011101100: data <= 12'hff3; 
        10'b0011101101: data <= 12'hff1; 
        10'b0011101110: data <= 12'hff1; 
        10'b0011101111: data <= 12'hff0; 
        10'b0011110000: data <= 12'hfed; 
        10'b0011110001: data <= 12'hfea; 
        10'b0011110010: data <= 12'hfe1; 
        10'b0011110011: data <= 12'hfe4; 
        10'b0011110100: data <= 12'hfe7; 
        10'b0011110101: data <= 12'hfe7; 
        10'b0011110110: data <= 12'hfee; 
        10'b0011110111: data <= 12'hff0; 
        10'b0011111000: data <= 12'hff6; 
        10'b0011111001: data <= 12'hffa; 
        10'b0011111010: data <= 12'hffc; 
        10'b0011111011: data <= 12'h001; 
        10'b0011111100: data <= 12'h000; 
        10'b0011111101: data <= 12'hffe; 
        10'b0011111110: data <= 12'hfff; 
        10'b0011111111: data <= 12'hffe; 
        10'b0100000000: data <= 12'h000; 
        10'b0100000001: data <= 12'hffe; 
        10'b0100000010: data <= 12'hffd; 
        10'b0100000011: data <= 12'hffe; 
        10'b0100000100: data <= 12'h002; 
        10'b0100000101: data <= 12'hffb; 
        10'b0100000110: data <= 12'hff7; 
        10'b0100000111: data <= 12'hff9; 
        10'b0100001000: data <= 12'hffb; 
        10'b0100001001: data <= 12'hff7; 
        10'b0100001010: data <= 12'hff8; 
        10'b0100001011: data <= 12'hfef; 
        10'b0100001100: data <= 12'hfec; 
        10'b0100001101: data <= 12'hfe3; 
        10'b0100001110: data <= 12'hfe1; 
        10'b0100001111: data <= 12'hfe6; 
        10'b0100010000: data <= 12'hfeb; 
        10'b0100010001: data <= 12'hfef; 
        10'b0100010010: data <= 12'hfed; 
        10'b0100010011: data <= 12'hff4; 
        10'b0100010100: data <= 12'hff7; 
        10'b0100010101: data <= 12'hff9; 
        10'b0100010110: data <= 12'hffd; 
        10'b0100010111: data <= 12'h002; 
        10'b0100011000: data <= 12'hfff; 
        10'b0100011001: data <= 12'h002; 
        10'b0100011010: data <= 12'h001; 
        10'b0100011011: data <= 12'hffe; 
        10'b0100011100: data <= 12'hffd; 
        10'b0100011101: data <= 12'h001; 
        10'b0100011110: data <= 12'h003; 
        10'b0100011111: data <= 12'h003; 
        10'b0100100000: data <= 12'h009; 
        10'b0100100001: data <= 12'h000; 
        10'b0100100010: data <= 12'h002; 
        10'b0100100011: data <= 12'h001; 
        10'b0100100100: data <= 12'hffa; 
        10'b0100100101: data <= 12'hffc; 
        10'b0100100110: data <= 12'hff7; 
        10'b0100100111: data <= 12'hfee; 
        10'b0100101000: data <= 12'hfee; 
        10'b0100101001: data <= 12'hfeb; 
        10'b0100101010: data <= 12'hfea; 
        10'b0100101011: data <= 12'hfee; 
        10'b0100101100: data <= 12'hff4; 
        10'b0100101101: data <= 12'hff7; 
        10'b0100101110: data <= 12'hff5; 
        10'b0100101111: data <= 12'hfff; 
        10'b0100110000: data <= 12'hff9; 
        10'b0100110001: data <= 12'hffb; 
        10'b0100110010: data <= 12'hffe; 
        10'b0100110011: data <= 12'hfff; 
        10'b0100110100: data <= 12'hfff; 
        10'b0100110101: data <= 12'h001; 
        10'b0100110110: data <= 12'hfff; 
        10'b0100110111: data <= 12'h000; 
        10'b0100111000: data <= 12'hfff; 
        10'b0100111001: data <= 12'h000; 
        10'b0100111010: data <= 12'hfff; 
        10'b0100111011: data <= 12'h008; 
        10'b0100111100: data <= 12'h006; 
        10'b0100111101: data <= 12'h003; 
        10'b0100111110: data <= 12'h003; 
        10'b0100111111: data <= 12'h002; 
        10'b0101000000: data <= 12'h002; 
        10'b0101000001: data <= 12'h000; 
        10'b0101000010: data <= 12'hffc; 
        10'b0101000011: data <= 12'hff2; 
        10'b0101000100: data <= 12'hff3; 
        10'b0101000101: data <= 12'hff5; 
        10'b0101000110: data <= 12'hff5; 
        10'b0101000111: data <= 12'hff7; 
        10'b0101001000: data <= 12'hffc; 
        10'b0101001001: data <= 12'h002; 
        10'b0101001010: data <= 12'h005; 
        10'b0101001011: data <= 12'h008; 
        10'b0101001100: data <= 12'h000; 
        10'b0101001101: data <= 12'hffb; 
        10'b0101001110: data <= 12'hffe; 
        10'b0101001111: data <= 12'hfff; 
        10'b0101010000: data <= 12'hfff; 
        10'b0101010001: data <= 12'hfff; 
        10'b0101010010: data <= 12'hffe; 
        10'b0101010011: data <= 12'hfff; 
        10'b0101010100: data <= 12'h001; 
        10'b0101010101: data <= 12'h004; 
        10'b0101010110: data <= 12'h006; 
        10'b0101010111: data <= 12'h007; 
        10'b0101011000: data <= 12'h003; 
        10'b0101011001: data <= 12'h005; 
        10'b0101011010: data <= 12'h003; 
        10'b0101011011: data <= 12'h009; 
        10'b0101011100: data <= 12'h009; 
        10'b0101011101: data <= 12'h006; 
        10'b0101011110: data <= 12'hffb; 
        10'b0101011111: data <= 12'hff6; 
        10'b0101100000: data <= 12'h000; 
        10'b0101100001: data <= 12'hfff; 
        10'b0101100010: data <= 12'hff7; 
        10'b0101100011: data <= 12'hff7; 
        10'b0101100100: data <= 12'hfff; 
        10'b0101100101: data <= 12'h005; 
        10'b0101100110: data <= 12'h00c; 
        10'b0101100111: data <= 12'h016; 
        10'b0101101000: data <= 12'h00c; 
        10'b0101101001: data <= 12'hffd; 
        10'b0101101010: data <= 12'hffc; 
        10'b0101101011: data <= 12'hfff; 
        10'b0101101100: data <= 12'hfff; 
        10'b0101101101: data <= 12'h002; 
        10'b0101101110: data <= 12'h002; 
        10'b0101101111: data <= 12'hffe; 
        10'b0101110000: data <= 12'hffd; 
        10'b0101110001: data <= 12'h001; 
        10'b0101110010: data <= 12'h009; 
        10'b0101110011: data <= 12'h005; 
        10'b0101110100: data <= 12'h004; 
        10'b0101110101: data <= 12'h002; 
        10'b0101110110: data <= 12'h009; 
        10'b0101110111: data <= 12'h008; 
        10'b0101111000: data <= 12'h007; 
        10'b0101111001: data <= 12'h001; 
        10'b0101111010: data <= 12'hfff; 
        10'b0101111011: data <= 12'h000; 
        10'b0101111100: data <= 12'h001; 
        10'b0101111101: data <= 12'hffe; 
        10'b0101111110: data <= 12'hff8; 
        10'b0101111111: data <= 12'hfff; 
        10'b0110000000: data <= 12'hffc; 
        10'b0110000001: data <= 12'h007; 
        10'b0110000010: data <= 12'h011; 
        10'b0110000011: data <= 12'h01b; 
        10'b0110000100: data <= 12'h00f; 
        10'b0110000101: data <= 12'hfff; 
        10'b0110000110: data <= 12'h000; 
        10'b0110000111: data <= 12'h001; 
        10'b0110001000: data <= 12'hfff; 
        10'b0110001001: data <= 12'h000; 
        10'b0110001010: data <= 12'h002; 
        10'b0110001011: data <= 12'h000; 
        10'b0110001100: data <= 12'hffd; 
        10'b0110001101: data <= 12'h003; 
        10'b0110001110: data <= 12'h009; 
        10'b0110001111: data <= 12'h007; 
        10'b0110010000: data <= 12'h00a; 
        10'b0110010001: data <= 12'h00a; 
        10'b0110010010: data <= 12'h00a; 
        10'b0110010011: data <= 12'h00b; 
        10'b0110010100: data <= 12'h004; 
        10'b0110010101: data <= 12'hffb; 
        10'b0110010110: data <= 12'h000; 
        10'b0110010111: data <= 12'h005; 
        10'b0110011000: data <= 12'h002; 
        10'b0110011001: data <= 12'hffc; 
        10'b0110011010: data <= 12'hffd; 
        10'b0110011011: data <= 12'h000; 
        10'b0110011100: data <= 12'h007; 
        10'b0110011101: data <= 12'h007; 
        10'b0110011110: data <= 12'h013; 
        10'b0110011111: data <= 12'h016; 
        10'b0110100000: data <= 12'h00f; 
        10'b0110100001: data <= 12'h000; 
        10'b0110100010: data <= 12'hffc; 
        10'b0110100011: data <= 12'hffe; 
        10'b0110100100: data <= 12'h002; 
        10'b0110100101: data <= 12'hfff; 
        10'b0110100110: data <= 12'h000; 
        10'b0110100111: data <= 12'hffe; 
        10'b0110101000: data <= 12'hffa; 
        10'b0110101001: data <= 12'hfff; 
        10'b0110101010: data <= 12'h009; 
        10'b0110101011: data <= 12'h00c; 
        10'b0110101100: data <= 12'h008; 
        10'b0110101101: data <= 12'h00c; 
        10'b0110101110: data <= 12'h00f; 
        10'b0110101111: data <= 12'h013; 
        10'b0110110000: data <= 12'h005; 
        10'b0110110001: data <= 12'hfff; 
        10'b0110110010: data <= 12'h007; 
        10'b0110110011: data <= 12'h007; 
        10'b0110110100: data <= 12'h001; 
        10'b0110110101: data <= 12'hffd; 
        10'b0110110110: data <= 12'h001; 
        10'b0110110111: data <= 12'h004; 
        10'b0110111000: data <= 12'h009; 
        10'b0110111001: data <= 12'h00c; 
        10'b0110111010: data <= 12'h00b; 
        10'b0110111011: data <= 12'h00d; 
        10'b0110111100: data <= 12'h007; 
        10'b0110111101: data <= 12'hffc; 
        10'b0110111110: data <= 12'hffe; 
        10'b0110111111: data <= 12'hffe; 
        10'b0111000000: data <= 12'h000; 
        10'b0111000001: data <= 12'hffe; 
        10'b0111000010: data <= 12'hffe; 
        10'b0111000011: data <= 12'hffe; 
        10'b0111000100: data <= 12'hff8; 
        10'b0111000101: data <= 12'hffc; 
        10'b0111000110: data <= 12'h00d; 
        10'b0111000111: data <= 12'h00e; 
        10'b0111001000: data <= 12'h009; 
        10'b0111001001: data <= 12'h00e; 
        10'b0111001010: data <= 12'h018; 
        10'b0111001011: data <= 12'h017; 
        10'b0111001100: data <= 12'h007; 
        10'b0111001101: data <= 12'h004; 
        10'b0111001110: data <= 12'h00a; 
        10'b0111001111: data <= 12'h005; 
        10'b0111010000: data <= 12'hffd; 
        10'b0111010001: data <= 12'hffa; 
        10'b0111010010: data <= 12'h002; 
        10'b0111010011: data <= 12'h006; 
        10'b0111010100: data <= 12'h003; 
        10'b0111010101: data <= 12'h000; 
        10'b0111010110: data <= 12'h006; 
        10'b0111010111: data <= 12'h003; 
        10'b0111011000: data <= 12'hffe; 
        10'b0111011001: data <= 12'hffc; 
        10'b0111011010: data <= 12'hffd; 
        10'b0111011011: data <= 12'h000; 
        10'b0111011100: data <= 12'h000; 
        10'b0111011101: data <= 12'h001; 
        10'b0111011110: data <= 12'h002; 
        10'b0111011111: data <= 12'h000; 
        10'b0111100000: data <= 12'hff5; 
        10'b0111100001: data <= 12'hffa; 
        10'b0111100010: data <= 12'h006; 
        10'b0111100011: data <= 12'h00b; 
        10'b0111100100: data <= 12'h00c; 
        10'b0111100101: data <= 12'h00f; 
        10'b0111100110: data <= 12'h01a; 
        10'b0111100111: data <= 12'h01b; 
        10'b0111101000: data <= 12'h00e; 
        10'b0111101001: data <= 12'h008; 
        10'b0111101010: data <= 12'h008; 
        10'b0111101011: data <= 12'h005; 
        10'b0111101100: data <= 12'h000; 
        10'b0111101101: data <= 12'h001; 
        10'b0111101110: data <= 12'h00b; 
        10'b0111101111: data <= 12'h004; 
        10'b0111110000: data <= 12'h002; 
        10'b0111110001: data <= 12'hffd; 
        10'b0111110010: data <= 12'h003; 
        10'b0111110011: data <= 12'hfff; 
        10'b0111110100: data <= 12'hffd; 
        10'b0111110101: data <= 12'hffa; 
        10'b0111110110: data <= 12'hfff; 
        10'b0111110111: data <= 12'h001; 
        10'b0111111000: data <= 12'hfff; 
        10'b0111111001: data <= 12'hfff; 
        10'b0111111010: data <= 12'h000; 
        10'b0111111011: data <= 12'hffd; 
        10'b0111111100: data <= 12'hff5; 
        10'b0111111101: data <= 12'hff6; 
        10'b0111111110: data <= 12'hffb; 
        10'b0111111111: data <= 12'h007; 
        10'b1000000000: data <= 12'h00c; 
        10'b1000000001: data <= 12'h00b; 
        10'b1000000010: data <= 12'h012; 
        10'b1000000011: data <= 12'h017; 
        10'b1000000100: data <= 12'h01b; 
        10'b1000000101: data <= 12'h00c; 
        10'b1000000110: data <= 12'h003; 
        10'b1000000111: data <= 12'h007; 
        10'b1000001000: data <= 12'h00c; 
        10'b1000001001: data <= 12'h008; 
        10'b1000001010: data <= 12'h00a; 
        10'b1000001011: data <= 12'h005; 
        10'b1000001100: data <= 12'h001; 
        10'b1000001101: data <= 12'h002; 
        10'b1000001110: data <= 12'h002; 
        10'b1000001111: data <= 12'hfff; 
        10'b1000010000: data <= 12'hffc; 
        10'b1000010001: data <= 12'hffd; 
        10'b1000010010: data <= 12'hffe; 
        10'b1000010011: data <= 12'hffe; 
        10'b1000010100: data <= 12'h001; 
        10'b1000010101: data <= 12'hffe; 
        10'b1000010110: data <= 12'h001; 
        10'b1000010111: data <= 12'hffc; 
        10'b1000011000: data <= 12'hff9; 
        10'b1000011001: data <= 12'hff5; 
        10'b1000011010: data <= 12'hff7; 
        10'b1000011011: data <= 12'h001; 
        10'b1000011100: data <= 12'h008; 
        10'b1000011101: data <= 12'h00c; 
        10'b1000011110: data <= 12'h010; 
        10'b1000011111: data <= 12'h019; 
        10'b1000100000: data <= 12'h01c; 
        10'b1000100001: data <= 12'h00f; 
        10'b1000100010: data <= 12'h00d; 
        10'b1000100011: data <= 12'h00e; 
        10'b1000100100: data <= 12'h00a; 
        10'b1000100101: data <= 12'h008; 
        10'b1000100110: data <= 12'h00d; 
        10'b1000100111: data <= 12'h009; 
        10'b1000101000: data <= 12'h006; 
        10'b1000101001: data <= 12'h001; 
        10'b1000101010: data <= 12'hffe; 
        10'b1000101011: data <= 12'hffe; 
        10'b1000101100: data <= 12'hffd; 
        10'b1000101101: data <= 12'h000; 
        10'b1000101110: data <= 12'hfff; 
        10'b1000101111: data <= 12'h002; 
        10'b1000110000: data <= 12'hfff; 
        10'b1000110001: data <= 12'hffe; 
        10'b1000110010: data <= 12'hfff; 
        10'b1000110011: data <= 12'hffe; 
        10'b1000110100: data <= 12'hff7; 
        10'b1000110101: data <= 12'hff5; 
        10'b1000110110: data <= 12'hff7; 
        10'b1000110111: data <= 12'hffc; 
        10'b1000111000: data <= 12'h003; 
        10'b1000111001: data <= 12'h008; 
        10'b1000111010: data <= 12'h00d; 
        10'b1000111011: data <= 12'h009; 
        10'b1000111100: data <= 12'h011; 
        10'b1000111101: data <= 12'h015; 
        10'b1000111110: data <= 12'h019; 
        10'b1000111111: data <= 12'h015; 
        10'b1001000000: data <= 12'h00b; 
        10'b1001000001: data <= 12'h007; 
        10'b1001000010: data <= 12'h00e; 
        10'b1001000011: data <= 12'h00a; 
        10'b1001000100: data <= 12'h007; 
        10'b1001000101: data <= 12'hfff; 
        10'b1001000110: data <= 12'hffb; 
        10'b1001000111: data <= 12'h000; 
        10'b1001001000: data <= 12'hfff; 
        10'b1001001001: data <= 12'hfff; 
        10'b1001001010: data <= 12'hffe; 
        10'b1001001011: data <= 12'h000; 
        10'b1001001100: data <= 12'h000; 
        10'b1001001101: data <= 12'h000; 
        10'b1001001110: data <= 12'h001; 
        10'b1001001111: data <= 12'hfff; 
        10'b1001010000: data <= 12'hffd; 
        10'b1001010001: data <= 12'hff9; 
        10'b1001010010: data <= 12'hff4; 
        10'b1001010011: data <= 12'hffa; 
        10'b1001010100: data <= 12'hffd; 
        10'b1001010101: data <= 12'h006; 
        10'b1001010110: data <= 12'h00b; 
        10'b1001010111: data <= 12'h010; 
        10'b1001011000: data <= 12'h014; 
        10'b1001011001: data <= 12'h014; 
        10'b1001011010: data <= 12'h011; 
        10'b1001011011: data <= 12'h00f; 
        10'b1001011100: data <= 12'h009; 
        10'b1001011101: data <= 12'h00d; 
        10'b1001011110: data <= 12'h00c; 
        10'b1001011111: data <= 12'h007; 
        10'b1001100000: data <= 12'h001; 
        10'b1001100001: data <= 12'hffc; 
        10'b1001100010: data <= 12'hffa; 
        10'b1001100011: data <= 12'hffd; 
        10'b1001100100: data <= 12'h000; 
        10'b1001100101: data <= 12'hffe; 
        10'b1001100110: data <= 12'h000; 
        10'b1001100111: data <= 12'hfff; 
        10'b1001101000: data <= 12'hfff; 
        10'b1001101001: data <= 12'h000; 
        10'b1001101010: data <= 12'h002; 
        10'b1001101011: data <= 12'h001; 
        10'b1001101100: data <= 12'hfff; 
        10'b1001101101: data <= 12'hffa; 
        10'b1001101110: data <= 12'hff8; 
        10'b1001101111: data <= 12'hff6; 
        10'b1001110000: data <= 12'hff9; 
        10'b1001110001: data <= 12'hffd; 
        10'b1001110010: data <= 12'hffd; 
        10'b1001110011: data <= 12'h001; 
        10'b1001110100: data <= 12'h006; 
        10'b1001110101: data <= 12'h003; 
        10'b1001110110: data <= 12'h002; 
        10'b1001110111: data <= 12'h006; 
        10'b1001111000: data <= 12'h005; 
        10'b1001111001: data <= 12'h000; 
        10'b1001111010: data <= 12'hffe; 
        10'b1001111011: data <= 12'hff9; 
        10'b1001111100: data <= 12'hff9; 
        10'b1001111101: data <= 12'hffa; 
        10'b1001111110: data <= 12'hffb; 
        10'b1001111111: data <= 12'hfff; 
        10'b1010000000: data <= 12'hfff; 
        10'b1010000001: data <= 12'hffe; 
        10'b1010000010: data <= 12'h002; 
        10'b1010000011: data <= 12'h001; 
        10'b1010000100: data <= 12'h002; 
        10'b1010000101: data <= 12'hfff; 
        10'b1010000110: data <= 12'hfff; 
        10'b1010000111: data <= 12'h000; 
        10'b1010001000: data <= 12'h001; 
        10'b1010001001: data <= 12'hffd; 
        10'b1010001010: data <= 12'hffc; 
        10'b1010001011: data <= 12'hff7; 
        10'b1010001100: data <= 12'hff5; 
        10'b1010001101: data <= 12'hff0; 
        10'b1010001110: data <= 12'hff0; 
        10'b1010001111: data <= 12'hfed; 
        10'b1010010000: data <= 12'hff4; 
        10'b1010010001: data <= 12'hff7; 
        10'b1010010010: data <= 12'hff9; 
        10'b1010010011: data <= 12'hff5; 
        10'b1010010100: data <= 12'hff2; 
        10'b1010010101: data <= 12'hff0; 
        10'b1010010110: data <= 12'hff3; 
        10'b1010010111: data <= 12'hffa; 
        10'b1010011000: data <= 12'hffa; 
        10'b1010011001: data <= 12'hffb; 
        10'b1010011010: data <= 12'hffe; 
        10'b1010011011: data <= 12'h000; 
        10'b1010011100: data <= 12'hffe; 
        10'b1010011101: data <= 12'hffe; 
        10'b1010011110: data <= 12'hfff; 
        10'b1010011111: data <= 12'h000; 
        10'b1010100000: data <= 12'h001; 
        10'b1010100001: data <= 12'h001; 
        10'b1010100010: data <= 12'h001; 
        10'b1010100011: data <= 12'hffe; 
        10'b1010100100: data <= 12'hffe; 
        10'b1010100101: data <= 12'hfff; 
        10'b1010100110: data <= 12'hffe; 
        10'b1010100111: data <= 12'hffd; 
        10'b1010101000: data <= 12'hffe; 
        10'b1010101001: data <= 12'hffc; 
        10'b1010101010: data <= 12'hffa; 
        10'b1010101011: data <= 12'hff8; 
        10'b1010101100: data <= 12'hff7; 
        10'b1010101101: data <= 12'hff7; 
        10'b1010101110: data <= 12'hff6; 
        10'b1010101111: data <= 12'hff6; 
        10'b1010110000: data <= 12'hff6; 
        10'b1010110001: data <= 12'hff8; 
        10'b1010110010: data <= 12'hffd; 
        10'b1010110011: data <= 12'hffd; 
        10'b1010110100: data <= 12'hfff; 
        10'b1010110101: data <= 12'hfff; 
        10'b1010110110: data <= 12'h001; 
        10'b1010110111: data <= 12'h000; 
        10'b1010111000: data <= 12'hffe; 
        10'b1010111001: data <= 12'hfff; 
        10'b1010111010: data <= 12'hffe; 
        10'b1010111011: data <= 12'hffe; 
        10'b1010111100: data <= 12'h002; 
        10'b1010111101: data <= 12'hffe; 
        10'b1010111110: data <= 12'h001; 
        10'b1010111111: data <= 12'hfff; 
        10'b1011000000: data <= 12'hfff; 
        10'b1011000001: data <= 12'h000; 
        10'b1011000010: data <= 12'h001; 
        10'b1011000011: data <= 12'h000; 
        10'b1011000100: data <= 12'hffe; 
        10'b1011000101: data <= 12'h001; 
        10'b1011000110: data <= 12'hffe; 
        10'b1011000111: data <= 12'h000; 
        10'b1011001000: data <= 12'h000; 
        10'b1011001001: data <= 12'hffe; 
        10'b1011001010: data <= 12'hfff; 
        10'b1011001011: data <= 12'hfff; 
        10'b1011001100: data <= 12'h000; 
        10'b1011001101: data <= 12'hffe; 
        10'b1011001110: data <= 12'hfff; 
        10'b1011001111: data <= 12'hffe; 
        10'b1011010000: data <= 12'hffe; 
        10'b1011010001: data <= 12'h000; 
        10'b1011010010: data <= 12'hfff; 
        10'b1011010011: data <= 12'h002; 
        10'b1011010100: data <= 12'h002; 
        10'b1011010101: data <= 12'h002; 
        10'b1011010110: data <= 12'h000; 
        10'b1011010111: data <= 12'h001; 
        10'b1011011000: data <= 12'h002; 
        10'b1011011001: data <= 12'h000; 
        10'b1011011010: data <= 12'h000; 
        10'b1011011011: data <= 12'h000; 
        10'b1011011100: data <= 12'hfff; 
        10'b1011011101: data <= 12'h002; 
        10'b1011011110: data <= 12'h001; 
        10'b1011011111: data <= 12'hfff; 
        10'b1011100000: data <= 12'hfff; 
        10'b1011100001: data <= 12'h001; 
        10'b1011100010: data <= 12'hfff; 
        10'b1011100011: data <= 12'h000; 
        10'b1011100100: data <= 12'hfff; 
        10'b1011100101: data <= 12'h001; 
        10'b1011100110: data <= 12'h001; 
        10'b1011100111: data <= 12'hffe; 
        10'b1011101000: data <= 12'hfff; 
        10'b1011101001: data <= 12'h002; 
        10'b1011101010: data <= 12'h001; 
        10'b1011101011: data <= 12'hfff; 
        10'b1011101100: data <= 12'h001; 
        10'b1011101101: data <= 12'h000; 
        10'b1011101110: data <= 12'hfff; 
        10'b1011101111: data <= 12'h001; 
        10'b1011110000: data <= 12'h001; 
        10'b1011110001: data <= 12'h000; 
        10'b1011110010: data <= 12'hfff; 
        10'b1011110011: data <= 12'hfff; 
        10'b1011110100: data <= 12'h002; 
        10'b1011110101: data <= 12'h000; 
        10'b1011110110: data <= 12'h001; 
        10'b1011110111: data <= 12'hfff; 
        10'b1011111000: data <= 12'h001; 
        10'b1011111001: data <= 12'h000; 
        10'b1011111010: data <= 12'h002; 
        10'b1011111011: data <= 12'h000; 
        10'b1011111100: data <= 12'h000; 
        10'b1011111101: data <= 12'hffe; 
        10'b1011111110: data <= 12'hffe; 
        10'b1011111111: data <= 12'h001; 
        10'b1100000000: data <= 12'hffe; 
        10'b1100000001: data <= 12'hffe; 
        10'b1100000010: data <= 12'hfff; 
        10'b1100000011: data <= 12'hffe; 
        10'b1100000100: data <= 12'hfff; 
        10'b1100000101: data <= 12'hfff; 
        10'b1100000110: data <= 12'hffe; 
        10'b1100000111: data <= 12'hfff; 
        10'b1100001000: data <= 12'hfff; 
        10'b1100001001: data <= 12'hfff; 
        10'b1100001010: data <= 12'h002; 
        10'b1100001011: data <= 12'hffe; 
        10'b1100001100: data <= 12'hfff; 
        10'b1100001101: data <= 12'hffe; 
        10'b1100001110: data <= 12'hfff; 
        10'b1100001111: data <= 12'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 7) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 13'h1fff; 
        10'b0000000001: data <= 13'h0003; 
        10'b0000000010: data <= 13'h1ffd; 
        10'b0000000011: data <= 13'h0000; 
        10'b0000000100: data <= 13'h0000; 
        10'b0000000101: data <= 13'h0000; 
        10'b0000000110: data <= 13'h0002; 
        10'b0000000111: data <= 13'h0005; 
        10'b0000001000: data <= 13'h1ffd; 
        10'b0000001001: data <= 13'h1ffe; 
        10'b0000001010: data <= 13'h1ffe; 
        10'b0000001011: data <= 13'h1ffd; 
        10'b0000001100: data <= 13'h0001; 
        10'b0000001101: data <= 13'h0004; 
        10'b0000001110: data <= 13'h0002; 
        10'b0000001111: data <= 13'h1ffc; 
        10'b0000010000: data <= 13'h1fff; 
        10'b0000010001: data <= 13'h0005; 
        10'b0000010010: data <= 13'h0001; 
        10'b0000010011: data <= 13'h0000; 
        10'b0000010100: data <= 13'h1ffc; 
        10'b0000010101: data <= 13'h1ffe; 
        10'b0000010110: data <= 13'h0001; 
        10'b0000010111: data <= 13'h0004; 
        10'b0000011000: data <= 13'h0002; 
        10'b0000011001: data <= 13'h0003; 
        10'b0000011010: data <= 13'h1ffc; 
        10'b0000011011: data <= 13'h1ffd; 
        10'b0000011100: data <= 13'h0003; 
        10'b0000011101: data <= 13'h0002; 
        10'b0000011110: data <= 13'h0003; 
        10'b0000011111: data <= 13'h1fff; 
        10'b0000100000: data <= 13'h1ffc; 
        10'b0000100001: data <= 13'h1ffe; 
        10'b0000100010: data <= 13'h0002; 
        10'b0000100011: data <= 13'h0007; 
        10'b0000100100: data <= 13'h0005; 
        10'b0000100101: data <= 13'h0001; 
        10'b0000100110: data <= 13'h0006; 
        10'b0000100111: data <= 13'h0006; 
        10'b0000101000: data <= 13'h0006; 
        10'b0000101001: data <= 13'h0006; 
        10'b0000101010: data <= 13'h0004; 
        10'b0000101011: data <= 13'h0004; 
        10'b0000101100: data <= 13'h1ffc; 
        10'b0000101101: data <= 13'h0004; 
        10'b0000101110: data <= 13'h0005; 
        10'b0000101111: data <= 13'h0003; 
        10'b0000110000: data <= 13'h1fff; 
        10'b0000110001: data <= 13'h1ffd; 
        10'b0000110010: data <= 13'h0005; 
        10'b0000110011: data <= 13'h0004; 
        10'b0000110100: data <= 13'h1ffe; 
        10'b0000110101: data <= 13'h0005; 
        10'b0000110110: data <= 13'h1fff; 
        10'b0000110111: data <= 13'h0003; 
        10'b0000111000: data <= 13'h1ffd; 
        10'b0000111001: data <= 13'h1ffd; 
        10'b0000111010: data <= 13'h1ffc; 
        10'b0000111011: data <= 13'h0000; 
        10'b0000111100: data <= 13'h0002; 
        10'b0000111101: data <= 13'h0001; 
        10'b0000111110: data <= 13'h0002; 
        10'b0000111111: data <= 13'h0007; 
        10'b0001000000: data <= 13'h0005; 
        10'b0001000001: data <= 13'h000a; 
        10'b0001000010: data <= 13'h000d; 
        10'b0001000011: data <= 13'h000e; 
        10'b0001000100: data <= 13'h000e; 
        10'b0001000101: data <= 13'h000f; 
        10'b0001000110: data <= 13'h0008; 
        10'b0001000111: data <= 13'h0005; 
        10'b0001001000: data <= 13'h000c; 
        10'b0001001001: data <= 13'h0005; 
        10'b0001001010: data <= 13'h0005; 
        10'b0001001011: data <= 13'h0006; 
        10'b0001001100: data <= 13'h0006; 
        10'b0001001101: data <= 13'h0003; 
        10'b0001001110: data <= 13'h0004; 
        10'b0001001111: data <= 13'h0001; 
        10'b0001010000: data <= 13'h0002; 
        10'b0001010001: data <= 13'h1fff; 
        10'b0001010010: data <= 13'h1ffc; 
        10'b0001010011: data <= 13'h0001; 
        10'b0001010100: data <= 13'h1ffc; 
        10'b0001010101: data <= 13'h0000; 
        10'b0001010110: data <= 13'h0003; 
        10'b0001010111: data <= 13'h0002; 
        10'b0001011000: data <= 13'h0004; 
        10'b0001011001: data <= 13'h1ffc; 
        10'b0001011010: data <= 13'h0005; 
        10'b0001011011: data <= 13'h0005; 
        10'b0001011100: data <= 13'h0006; 
        10'b0001011101: data <= 13'h000d; 
        10'b0001011110: data <= 13'h000b; 
        10'b0001011111: data <= 13'h000e; 
        10'b0001100000: data <= 13'h000e; 
        10'b0001100001: data <= 13'h000d; 
        10'b0001100010: data <= 13'h0013; 
        10'b0001100011: data <= 13'h0012; 
        10'b0001100100: data <= 13'h000b; 
        10'b0001100101: data <= 13'h000e; 
        10'b0001100110: data <= 13'h0017; 
        10'b0001100111: data <= 13'h0017; 
        10'b0001101000: data <= 13'h0019; 
        10'b0001101001: data <= 13'h0016; 
        10'b0001101010: data <= 13'h0016; 
        10'b0001101011: data <= 13'h000d; 
        10'b0001101100: data <= 13'h000b; 
        10'b0001101101: data <= 13'h0003; 
        10'b0001101110: data <= 13'h1ffe; 
        10'b0001101111: data <= 13'h0003; 
        10'b0001110000: data <= 13'h0001; 
        10'b0001110001: data <= 13'h1fff; 
        10'b0001110010: data <= 13'h0000; 
        10'b0001110011: data <= 13'h0004; 
        10'b0001110100: data <= 13'h0003; 
        10'b0001110101: data <= 13'h0001; 
        10'b0001110110: data <= 13'h0001; 
        10'b0001110111: data <= 13'h0008; 
        10'b0001111000: data <= 13'h1fff; 
        10'b0001111001: data <= 13'h1ffe; 
        10'b0001111010: data <= 13'h0008; 
        10'b0001111011: data <= 13'h0003; 
        10'b0001111100: data <= 13'h0004; 
        10'b0001111101: data <= 13'h0001; 
        10'b0001111110: data <= 13'h0003; 
        10'b0001111111: data <= 13'h0004; 
        10'b0010000000: data <= 13'h000f; 
        10'b0010000001: data <= 13'h000f; 
        10'b0010000010: data <= 13'h0018; 
        10'b0010000011: data <= 13'h0018; 
        10'b0010000100: data <= 13'h001f; 
        10'b0010000101: data <= 13'h0022; 
        10'b0010000110: data <= 13'h001d; 
        10'b0010000111: data <= 13'h0014; 
        10'b0010001000: data <= 13'h0003; 
        10'b0010001001: data <= 13'h0005; 
        10'b0010001010: data <= 13'h0001; 
        10'b0010001011: data <= 13'h0000; 
        10'b0010001100: data <= 13'h0001; 
        10'b0010001101: data <= 13'h0002; 
        10'b0010001110: data <= 13'h0001; 
        10'b0010001111: data <= 13'h1ffe; 
        10'b0010010000: data <= 13'h1ffd; 
        10'b0010010001: data <= 13'h0000; 
        10'b0010010010: data <= 13'h1ffd; 
        10'b0010010011: data <= 13'h1ffb; 
        10'b0010010100: data <= 13'h0004; 
        10'b0010010101: data <= 13'h1ffb; 
        10'b0010010110: data <= 13'h0002; 
        10'b0010010111: data <= 13'h1fee; 
        10'b0010011000: data <= 13'h1ff7; 
        10'b0010011001: data <= 13'h1ff9; 
        10'b0010011010: data <= 13'h1ffe; 
        10'b0010011011: data <= 13'h1ff8; 
        10'b0010011100: data <= 13'h1ff8; 
        10'b0010011101: data <= 13'h0002; 
        10'b0010011110: data <= 13'h000b; 
        10'b0010011111: data <= 13'h0015; 
        10'b0010100000: data <= 13'h0013; 
        10'b0010100001: data <= 13'h0011; 
        10'b0010100010: data <= 13'h000d; 
        10'b0010100011: data <= 13'h0009; 
        10'b0010100100: data <= 13'h1fff; 
        10'b0010100101: data <= 13'h0000; 
        10'b0010100110: data <= 13'h1ffb; 
        10'b0010100111: data <= 13'h0004; 
        10'b0010101000: data <= 13'h1fff; 
        10'b0010101001: data <= 13'h0004; 
        10'b0010101010: data <= 13'h0004; 
        10'b0010101011: data <= 13'h1ffb; 
        10'b0010101100: data <= 13'h0002; 
        10'b0010101101: data <= 13'h1fff; 
        10'b0010101110: data <= 13'h0001; 
        10'b0010101111: data <= 13'h0000; 
        10'b0010110000: data <= 13'h1ff9; 
        10'b0010110001: data <= 13'h1ff8; 
        10'b0010110010: data <= 13'h1feb; 
        10'b0010110011: data <= 13'h1fe5; 
        10'b0010110100: data <= 13'h1ff0; 
        10'b0010110101: data <= 13'h1fe1; 
        10'b0010110110: data <= 13'h1ff2; 
        10'b0010110111: data <= 13'h1ff6; 
        10'b0010111000: data <= 13'h1ff2; 
        10'b0010111001: data <= 13'h1ff4; 
        10'b0010111010: data <= 13'h1ffd; 
        10'b0010111011: data <= 13'h1ff8; 
        10'b0010111100: data <= 13'h1ff2; 
        10'b0010111101: data <= 13'h1ff3; 
        10'b0010111110: data <= 13'h1fec; 
        10'b0010111111: data <= 13'h1ff3; 
        10'b0011000000: data <= 13'h1ff5; 
        10'b0011000001: data <= 13'h1ff5; 
        10'b0011000010: data <= 13'h1ffe; 
        10'b0011000011: data <= 13'h0004; 
        10'b0011000100: data <= 13'h0001; 
        10'b0011000101: data <= 13'h0002; 
        10'b0011000110: data <= 13'h0000; 
        10'b0011000111: data <= 13'h1fff; 
        10'b0011001000: data <= 13'h0000; 
        10'b0011001001: data <= 13'h1ffc; 
        10'b0011001010: data <= 13'h1ff8; 
        10'b0011001011: data <= 13'h1fff; 
        10'b0011001100: data <= 13'h1ff5; 
        10'b0011001101: data <= 13'h1ff2; 
        10'b0011001110: data <= 13'h1feb; 
        10'b0011001111: data <= 13'h1ff0; 
        10'b0011010000: data <= 13'h1fe3; 
        10'b0011010001: data <= 13'h1fdf; 
        10'b0011010010: data <= 13'h1fef; 
        10'b0011010011: data <= 13'h1ff0; 
        10'b0011010100: data <= 13'h1fe6; 
        10'b0011010101: data <= 13'h1fe8; 
        10'b0011010110: data <= 13'h1fe2; 
        10'b0011010111: data <= 13'h1fd7; 
        10'b0011011000: data <= 13'h1fd6; 
        10'b0011011001: data <= 13'h1fdd; 
        10'b0011011010: data <= 13'h1fdc; 
        10'b0011011011: data <= 13'h1fe3; 
        10'b0011011100: data <= 13'h1ff5; 
        10'b0011011101: data <= 13'h1ff6; 
        10'b0011011110: data <= 13'h1ffc; 
        10'b0011011111: data <= 13'h1ffd; 
        10'b0011100000: data <= 13'h1fff; 
        10'b0011100001: data <= 13'h1fff; 
        10'b0011100010: data <= 13'h0004; 
        10'b0011100011: data <= 13'h1ffa; 
        10'b0011100100: data <= 13'h1ffb; 
        10'b0011100101: data <= 13'h1ffa; 
        10'b0011100110: data <= 13'h1ff0; 
        10'b0011100111: data <= 13'h1ffd; 
        10'b0011101000: data <= 13'h1ffa; 
        10'b0011101001: data <= 13'h1ff0; 
        10'b0011101010: data <= 13'h1fed; 
        10'b0011101011: data <= 13'h1fea; 
        10'b0011101100: data <= 13'h1fe6; 
        10'b0011101101: data <= 13'h1fe2; 
        10'b0011101110: data <= 13'h1fe2; 
        10'b0011101111: data <= 13'h1fe0; 
        10'b0011110000: data <= 13'h1fda; 
        10'b0011110001: data <= 13'h1fd5; 
        10'b0011110010: data <= 13'h1fc3; 
        10'b0011110011: data <= 13'h1fc7; 
        10'b0011110100: data <= 13'h1fcd; 
        10'b0011110101: data <= 13'h1fce; 
        10'b0011110110: data <= 13'h1fdd; 
        10'b0011110111: data <= 13'h1fe1; 
        10'b0011111000: data <= 13'h1fed; 
        10'b0011111001: data <= 13'h1ff4; 
        10'b0011111010: data <= 13'h1ff7; 
        10'b0011111011: data <= 13'h0001; 
        10'b0011111100: data <= 13'h1fff; 
        10'b0011111101: data <= 13'h1ffd; 
        10'b0011111110: data <= 13'h1ffe; 
        10'b0011111111: data <= 13'h1ffc; 
        10'b0100000000: data <= 13'h0000; 
        10'b0100000001: data <= 13'h1ffc; 
        10'b0100000010: data <= 13'h1ffb; 
        10'b0100000011: data <= 13'h1ffd; 
        10'b0100000100: data <= 13'h0004; 
        10'b0100000101: data <= 13'h1ff6; 
        10'b0100000110: data <= 13'h1fed; 
        10'b0100000111: data <= 13'h1ff2; 
        10'b0100001000: data <= 13'h1ff7; 
        10'b0100001001: data <= 13'h1fef; 
        10'b0100001010: data <= 13'h1ff0; 
        10'b0100001011: data <= 13'h1fdd; 
        10'b0100001100: data <= 13'h1fd8; 
        10'b0100001101: data <= 13'h1fc5; 
        10'b0100001110: data <= 13'h1fc1; 
        10'b0100001111: data <= 13'h1fcd; 
        10'b0100010000: data <= 13'h1fd6; 
        10'b0100010001: data <= 13'h1fdf; 
        10'b0100010010: data <= 13'h1fd9; 
        10'b0100010011: data <= 13'h1fe7; 
        10'b0100010100: data <= 13'h1fed; 
        10'b0100010101: data <= 13'h1ff2; 
        10'b0100010110: data <= 13'h1ffa; 
        10'b0100010111: data <= 13'h0003; 
        10'b0100011000: data <= 13'h1ffd; 
        10'b0100011001: data <= 13'h0004; 
        10'b0100011010: data <= 13'h0003; 
        10'b0100011011: data <= 13'h1ffb; 
        10'b0100011100: data <= 13'h1ff9; 
        10'b0100011101: data <= 13'h0002; 
        10'b0100011110: data <= 13'h0005; 
        10'b0100011111: data <= 13'h0005; 
        10'b0100100000: data <= 13'h0013; 
        10'b0100100001: data <= 13'h0000; 
        10'b0100100010: data <= 13'h0004; 
        10'b0100100011: data <= 13'h0002; 
        10'b0100100100: data <= 13'h1ff5; 
        10'b0100100101: data <= 13'h1ff8; 
        10'b0100100110: data <= 13'h1fef; 
        10'b0100100111: data <= 13'h1fdc; 
        10'b0100101000: data <= 13'h1fdb; 
        10'b0100101001: data <= 13'h1fd5; 
        10'b0100101010: data <= 13'h1fd3; 
        10'b0100101011: data <= 13'h1fdc; 
        10'b0100101100: data <= 13'h1fe8; 
        10'b0100101101: data <= 13'h1fef; 
        10'b0100101110: data <= 13'h1fe9; 
        10'b0100101111: data <= 13'h1ffe; 
        10'b0100110000: data <= 13'h1ff1; 
        10'b0100110001: data <= 13'h1ff6; 
        10'b0100110010: data <= 13'h1ffd; 
        10'b0100110011: data <= 13'h1fff; 
        10'b0100110100: data <= 13'h1ffe; 
        10'b0100110101: data <= 13'h0002; 
        10'b0100110110: data <= 13'h1ffd; 
        10'b0100110111: data <= 13'h0000; 
        10'b0100111000: data <= 13'h1ffd; 
        10'b0100111001: data <= 13'h0001; 
        10'b0100111010: data <= 13'h1fff; 
        10'b0100111011: data <= 13'h0010; 
        10'b0100111100: data <= 13'h000b; 
        10'b0100111101: data <= 13'h0005; 
        10'b0100111110: data <= 13'h0007; 
        10'b0100111111: data <= 13'h0005; 
        10'b0101000000: data <= 13'h0005; 
        10'b0101000001: data <= 13'h0001; 
        10'b0101000010: data <= 13'h1ff8; 
        10'b0101000011: data <= 13'h1fe3; 
        10'b0101000100: data <= 13'h1fe5; 
        10'b0101000101: data <= 13'h1fe9; 
        10'b0101000110: data <= 13'h1fe9; 
        10'b0101000111: data <= 13'h1fee; 
        10'b0101001000: data <= 13'h1ff8; 
        10'b0101001001: data <= 13'h0003; 
        10'b0101001010: data <= 13'h000b; 
        10'b0101001011: data <= 13'h0011; 
        10'b0101001100: data <= 13'h0000; 
        10'b0101001101: data <= 13'h1ff7; 
        10'b0101001110: data <= 13'h1ffc; 
        10'b0101001111: data <= 13'h1fff; 
        10'b0101010000: data <= 13'h1ffe; 
        10'b0101010001: data <= 13'h1fff; 
        10'b0101010010: data <= 13'h1ffc; 
        10'b0101010011: data <= 13'h1ffe; 
        10'b0101010100: data <= 13'h0002; 
        10'b0101010101: data <= 13'h0007; 
        10'b0101010110: data <= 13'h000b; 
        10'b0101010111: data <= 13'h000f; 
        10'b0101011000: data <= 13'h0007; 
        10'b0101011001: data <= 13'h000a; 
        10'b0101011010: data <= 13'h0007; 
        10'b0101011011: data <= 13'h0012; 
        10'b0101011100: data <= 13'h0011; 
        10'b0101011101: data <= 13'h000c; 
        10'b0101011110: data <= 13'h1ff5; 
        10'b0101011111: data <= 13'h1fed; 
        10'b0101100000: data <= 13'h1fff; 
        10'b0101100001: data <= 13'h1ffe; 
        10'b0101100010: data <= 13'h1fed; 
        10'b0101100011: data <= 13'h1fee; 
        10'b0101100100: data <= 13'h1ffe; 
        10'b0101100101: data <= 13'h000a; 
        10'b0101100110: data <= 13'h0019; 
        10'b0101100111: data <= 13'h002b; 
        10'b0101101000: data <= 13'h0017; 
        10'b0101101001: data <= 13'h1ff9; 
        10'b0101101010: data <= 13'h1ff8; 
        10'b0101101011: data <= 13'h1ffe; 
        10'b0101101100: data <= 13'h1ffe; 
        10'b0101101101: data <= 13'h0004; 
        10'b0101101110: data <= 13'h0003; 
        10'b0101101111: data <= 13'h1ffc; 
        10'b0101110000: data <= 13'h1ffa; 
        10'b0101110001: data <= 13'h0002; 
        10'b0101110010: data <= 13'h0013; 
        10'b0101110011: data <= 13'h000a; 
        10'b0101110100: data <= 13'h0009; 
        10'b0101110101: data <= 13'h0004; 
        10'b0101110110: data <= 13'h0012; 
        10'b0101110111: data <= 13'h000f; 
        10'b0101111000: data <= 13'h000e; 
        10'b0101111001: data <= 13'h0002; 
        10'b0101111010: data <= 13'h1ffd; 
        10'b0101111011: data <= 13'h0000; 
        10'b0101111100: data <= 13'h0001; 
        10'b0101111101: data <= 13'h1ffc; 
        10'b0101111110: data <= 13'h1ff0; 
        10'b0101111111: data <= 13'h1ffe; 
        10'b0110000000: data <= 13'h1ff8; 
        10'b0110000001: data <= 13'h000d; 
        10'b0110000010: data <= 13'h0022; 
        10'b0110000011: data <= 13'h0036; 
        10'b0110000100: data <= 13'h001d; 
        10'b0110000101: data <= 13'h1ffe; 
        10'b0110000110: data <= 13'h0000; 
        10'b0110000111: data <= 13'h0003; 
        10'b0110001000: data <= 13'h1ffe; 
        10'b0110001001: data <= 13'h0000; 
        10'b0110001010: data <= 13'h0003; 
        10'b0110001011: data <= 13'h0000; 
        10'b0110001100: data <= 13'h1ffa; 
        10'b0110001101: data <= 13'h0007; 
        10'b0110001110: data <= 13'h0011; 
        10'b0110001111: data <= 13'h000f; 
        10'b0110010000: data <= 13'h0015; 
        10'b0110010001: data <= 13'h0013; 
        10'b0110010010: data <= 13'h0015; 
        10'b0110010011: data <= 13'h0017; 
        10'b0110010100: data <= 13'h0008; 
        10'b0110010101: data <= 13'h1ff5; 
        10'b0110010110: data <= 13'h0001; 
        10'b0110010111: data <= 13'h0009; 
        10'b0110011000: data <= 13'h0004; 
        10'b0110011001: data <= 13'h1ff9; 
        10'b0110011010: data <= 13'h1ff9; 
        10'b0110011011: data <= 13'h1fff; 
        10'b0110011100: data <= 13'h000f; 
        10'b0110011101: data <= 13'h000f; 
        10'b0110011110: data <= 13'h0026; 
        10'b0110011111: data <= 13'h002d; 
        10'b0110100000: data <= 13'h001d; 
        10'b0110100001: data <= 13'h0000; 
        10'b0110100010: data <= 13'h1ff8; 
        10'b0110100011: data <= 13'h1ffc; 
        10'b0110100100: data <= 13'h0003; 
        10'b0110100101: data <= 13'h1ffe; 
        10'b0110100110: data <= 13'h0001; 
        10'b0110100111: data <= 13'h1ffd; 
        10'b0110101000: data <= 13'h1ff4; 
        10'b0110101001: data <= 13'h1ffe; 
        10'b0110101010: data <= 13'h0012; 
        10'b0110101011: data <= 13'h0018; 
        10'b0110101100: data <= 13'h000f; 
        10'b0110101101: data <= 13'h0018; 
        10'b0110101110: data <= 13'h001f; 
        10'b0110101111: data <= 13'h0025; 
        10'b0110110000: data <= 13'h000a; 
        10'b0110110001: data <= 13'h1ffd; 
        10'b0110110010: data <= 13'h000e; 
        10'b0110110011: data <= 13'h000d; 
        10'b0110110100: data <= 13'h0002; 
        10'b0110110101: data <= 13'h1ff9; 
        10'b0110110110: data <= 13'h0001; 
        10'b0110110111: data <= 13'h0007; 
        10'b0110111000: data <= 13'h0011; 
        10'b0110111001: data <= 13'h0018; 
        10'b0110111010: data <= 13'h0016; 
        10'b0110111011: data <= 13'h001b; 
        10'b0110111100: data <= 13'h000e; 
        10'b0110111101: data <= 13'h1ff9; 
        10'b0110111110: data <= 13'h1ffb; 
        10'b0110111111: data <= 13'h1ffb; 
        10'b0111000000: data <= 13'h0001; 
        10'b0111000001: data <= 13'h1ffd; 
        10'b0111000010: data <= 13'h1ffc; 
        10'b0111000011: data <= 13'h1ffc; 
        10'b0111000100: data <= 13'h1ff0; 
        10'b0111000101: data <= 13'h1ff7; 
        10'b0111000110: data <= 13'h001b; 
        10'b0111000111: data <= 13'h001b; 
        10'b0111001000: data <= 13'h0012; 
        10'b0111001001: data <= 13'h001c; 
        10'b0111001010: data <= 13'h002f; 
        10'b0111001011: data <= 13'h002f; 
        10'b0111001100: data <= 13'h000e; 
        10'b0111001101: data <= 13'h0009; 
        10'b0111001110: data <= 13'h0014; 
        10'b0111001111: data <= 13'h000b; 
        10'b0111010000: data <= 13'h1ffa; 
        10'b0111010001: data <= 13'h1ff5; 
        10'b0111010010: data <= 13'h0004; 
        10'b0111010011: data <= 13'h000c; 
        10'b0111010100: data <= 13'h0006; 
        10'b0111010101: data <= 13'h0000; 
        10'b0111010110: data <= 13'h000b; 
        10'b0111010111: data <= 13'h0007; 
        10'b0111011000: data <= 13'h1ffd; 
        10'b0111011001: data <= 13'h1ff7; 
        10'b0111011010: data <= 13'h1ffb; 
        10'b0111011011: data <= 13'h1fff; 
        10'b0111011100: data <= 13'h0001; 
        10'b0111011101: data <= 13'h0003; 
        10'b0111011110: data <= 13'h0004; 
        10'b0111011111: data <= 13'h1fff; 
        10'b0111100000: data <= 13'h1fe9; 
        10'b0111100001: data <= 13'h1ff4; 
        10'b0111100010: data <= 13'h000b; 
        10'b0111100011: data <= 13'h0015; 
        10'b0111100100: data <= 13'h0018; 
        10'b0111100101: data <= 13'h001e; 
        10'b0111100110: data <= 13'h0035; 
        10'b0111100111: data <= 13'h0035; 
        10'b0111101000: data <= 13'h001c; 
        10'b0111101001: data <= 13'h0010; 
        10'b0111101010: data <= 13'h0010; 
        10'b0111101011: data <= 13'h000a; 
        10'b0111101100: data <= 13'h0000; 
        10'b0111101101: data <= 13'h0003; 
        10'b0111101110: data <= 13'h0016; 
        10'b0111101111: data <= 13'h0008; 
        10'b0111110000: data <= 13'h0003; 
        10'b0111110001: data <= 13'h1ffa; 
        10'b0111110010: data <= 13'h0005; 
        10'b0111110011: data <= 13'h1fff; 
        10'b0111110100: data <= 13'h1ffa; 
        10'b0111110101: data <= 13'h1ff4; 
        10'b0111110110: data <= 13'h1ffe; 
        10'b0111110111: data <= 13'h0002; 
        10'b0111111000: data <= 13'h1ffe; 
        10'b0111111001: data <= 13'h1ffe; 
        10'b0111111010: data <= 13'h0000; 
        10'b0111111011: data <= 13'h1ff9; 
        10'b0111111100: data <= 13'h1feb; 
        10'b0111111101: data <= 13'h1feb; 
        10'b0111111110: data <= 13'h1ff6; 
        10'b0111111111: data <= 13'h000f; 
        10'b1000000000: data <= 13'h0017; 
        10'b1000000001: data <= 13'h0015; 
        10'b1000000010: data <= 13'h0025; 
        10'b1000000011: data <= 13'h002d; 
        10'b1000000100: data <= 13'h0036; 
        10'b1000000101: data <= 13'h0019; 
        10'b1000000110: data <= 13'h0007; 
        10'b1000000111: data <= 13'h000e; 
        10'b1000001000: data <= 13'h0018; 
        10'b1000001001: data <= 13'h000f; 
        10'b1000001010: data <= 13'h0013; 
        10'b1000001011: data <= 13'h000a; 
        10'b1000001100: data <= 13'h0001; 
        10'b1000001101: data <= 13'h0003; 
        10'b1000001110: data <= 13'h0004; 
        10'b1000001111: data <= 13'h1ffe; 
        10'b1000010000: data <= 13'h1ff8; 
        10'b1000010001: data <= 13'h1ffa; 
        10'b1000010010: data <= 13'h1ffc; 
        10'b1000010011: data <= 13'h1ffb; 
        10'b1000010100: data <= 13'h0001; 
        10'b1000010101: data <= 13'h1ffd; 
        10'b1000010110: data <= 13'h0002; 
        10'b1000010111: data <= 13'h1ff8; 
        10'b1000011000: data <= 13'h1ff2; 
        10'b1000011001: data <= 13'h1fea; 
        10'b1000011010: data <= 13'h1fef; 
        10'b1000011011: data <= 13'h0001; 
        10'b1000011100: data <= 13'h000f; 
        10'b1000011101: data <= 13'h0018; 
        10'b1000011110: data <= 13'h0020; 
        10'b1000011111: data <= 13'h0033; 
        10'b1000100000: data <= 13'h0039; 
        10'b1000100001: data <= 13'h001d; 
        10'b1000100010: data <= 13'h001a; 
        10'b1000100011: data <= 13'h001b; 
        10'b1000100100: data <= 13'h0014; 
        10'b1000100101: data <= 13'h0010; 
        10'b1000100110: data <= 13'h0019; 
        10'b1000100111: data <= 13'h0011; 
        10'b1000101000: data <= 13'h000b; 
        10'b1000101001: data <= 13'h0002; 
        10'b1000101010: data <= 13'h1ffc; 
        10'b1000101011: data <= 13'h1ffb; 
        10'b1000101100: data <= 13'h1ffb; 
        10'b1000101101: data <= 13'h1fff; 
        10'b1000101110: data <= 13'h1ffe; 
        10'b1000101111: data <= 13'h0004; 
        10'b1000110000: data <= 13'h1ffe; 
        10'b1000110001: data <= 13'h1ffd; 
        10'b1000110010: data <= 13'h1fff; 
        10'b1000110011: data <= 13'h1ffc; 
        10'b1000110100: data <= 13'h1fee; 
        10'b1000110101: data <= 13'h1feb; 
        10'b1000110110: data <= 13'h1fee; 
        10'b1000110111: data <= 13'h1ff8; 
        10'b1000111000: data <= 13'h0005; 
        10'b1000111001: data <= 13'h0010; 
        10'b1000111010: data <= 13'h001a; 
        10'b1000111011: data <= 13'h0012; 
        10'b1000111100: data <= 13'h0023; 
        10'b1000111101: data <= 13'h0029; 
        10'b1000111110: data <= 13'h0031; 
        10'b1000111111: data <= 13'h002a; 
        10'b1001000000: data <= 13'h0017; 
        10'b1001000001: data <= 13'h000f; 
        10'b1001000010: data <= 13'h001c; 
        10'b1001000011: data <= 13'h0014; 
        10'b1001000100: data <= 13'h000d; 
        10'b1001000101: data <= 13'h1ffd; 
        10'b1001000110: data <= 13'h1ff6; 
        10'b1001000111: data <= 13'h0001; 
        10'b1001001000: data <= 13'h1ffd; 
        10'b1001001001: data <= 13'h1fff; 
        10'b1001001010: data <= 13'h1ffd; 
        10'b1001001011: data <= 13'h0001; 
        10'b1001001100: data <= 13'h0000; 
        10'b1001001101: data <= 13'h0000; 
        10'b1001001110: data <= 13'h0001; 
        10'b1001001111: data <= 13'h1fff; 
        10'b1001010000: data <= 13'h1ff9; 
        10'b1001010001: data <= 13'h1ff1; 
        10'b1001010010: data <= 13'h1fe7; 
        10'b1001010011: data <= 13'h1ff5; 
        10'b1001010100: data <= 13'h1ff9; 
        10'b1001010101: data <= 13'h000c; 
        10'b1001010110: data <= 13'h0016; 
        10'b1001010111: data <= 13'h001f; 
        10'b1001011000: data <= 13'h0028; 
        10'b1001011001: data <= 13'h0029; 
        10'b1001011010: data <= 13'h0022; 
        10'b1001011011: data <= 13'h001d; 
        10'b1001011100: data <= 13'h0012; 
        10'b1001011101: data <= 13'h0019; 
        10'b1001011110: data <= 13'h0017; 
        10'b1001011111: data <= 13'h000f; 
        10'b1001100000: data <= 13'h0002; 
        10'b1001100001: data <= 13'h1ff8; 
        10'b1001100010: data <= 13'h1ff5; 
        10'b1001100011: data <= 13'h1ffa; 
        10'b1001100100: data <= 13'h0000; 
        10'b1001100101: data <= 13'h1ffc; 
        10'b1001100110: data <= 13'h1fff; 
        10'b1001100111: data <= 13'h1ffe; 
        10'b1001101000: data <= 13'h1ffe; 
        10'b1001101001: data <= 13'h0000; 
        10'b1001101010: data <= 13'h0004; 
        10'b1001101011: data <= 13'h0001; 
        10'b1001101100: data <= 13'h1ffe; 
        10'b1001101101: data <= 13'h1ff3; 
        10'b1001101110: data <= 13'h1ff1; 
        10'b1001101111: data <= 13'h1fec; 
        10'b1001110000: data <= 13'h1ff2; 
        10'b1001110001: data <= 13'h1ffa; 
        10'b1001110010: data <= 13'h1ffb; 
        10'b1001110011: data <= 13'h0002; 
        10'b1001110100: data <= 13'h000c; 
        10'b1001110101: data <= 13'h0005; 
        10'b1001110110: data <= 13'h0004; 
        10'b1001110111: data <= 13'h000d; 
        10'b1001111000: data <= 13'h0009; 
        10'b1001111001: data <= 13'h0000; 
        10'b1001111010: data <= 13'h1ffd; 
        10'b1001111011: data <= 13'h1ff2; 
        10'b1001111100: data <= 13'h1ff2; 
        10'b1001111101: data <= 13'h1ff5; 
        10'b1001111110: data <= 13'h1ff5; 
        10'b1001111111: data <= 13'h1fff; 
        10'b1010000000: data <= 13'h1ffe; 
        10'b1010000001: data <= 13'h1ffc; 
        10'b1010000010: data <= 13'h0004; 
        10'b1010000011: data <= 13'h0002; 
        10'b1010000100: data <= 13'h0003; 
        10'b1010000101: data <= 13'h1fff; 
        10'b1010000110: data <= 13'h1ffe; 
        10'b1010000111: data <= 13'h0000; 
        10'b1010001000: data <= 13'h0001; 
        10'b1010001001: data <= 13'h1ffb; 
        10'b1010001010: data <= 13'h1ff8; 
        10'b1010001011: data <= 13'h1fee; 
        10'b1010001100: data <= 13'h1fe9; 
        10'b1010001101: data <= 13'h1fdf; 
        10'b1010001110: data <= 13'h1fdf; 
        10'b1010001111: data <= 13'h1fda; 
        10'b1010010000: data <= 13'h1fe8; 
        10'b1010010001: data <= 13'h1fed; 
        10'b1010010010: data <= 13'h1ff2; 
        10'b1010010011: data <= 13'h1feb; 
        10'b1010010100: data <= 13'h1fe4; 
        10'b1010010101: data <= 13'h1fe0; 
        10'b1010010110: data <= 13'h1fe7; 
        10'b1010010111: data <= 13'h1ff4; 
        10'b1010011000: data <= 13'h1ff4; 
        10'b1010011001: data <= 13'h1ff6; 
        10'b1010011010: data <= 13'h1ffc; 
        10'b1010011011: data <= 13'h0001; 
        10'b1010011100: data <= 13'h1ffc; 
        10'b1010011101: data <= 13'h1ffc; 
        10'b1010011110: data <= 13'h1ffe; 
        10'b1010011111: data <= 13'h0000; 
        10'b1010100000: data <= 13'h0002; 
        10'b1010100001: data <= 13'h0002; 
        10'b1010100010: data <= 13'h0001; 
        10'b1010100011: data <= 13'h1ffc; 
        10'b1010100100: data <= 13'h1ffd; 
        10'b1010100101: data <= 13'h1ffe; 
        10'b1010100110: data <= 13'h1ffc; 
        10'b1010100111: data <= 13'h1ffa; 
        10'b1010101000: data <= 13'h1ffb; 
        10'b1010101001: data <= 13'h1ff8; 
        10'b1010101010: data <= 13'h1ff4; 
        10'b1010101011: data <= 13'h1ff1; 
        10'b1010101100: data <= 13'h1fee; 
        10'b1010101101: data <= 13'h1fef; 
        10'b1010101110: data <= 13'h1fec; 
        10'b1010101111: data <= 13'h1fec; 
        10'b1010110000: data <= 13'h1feb; 
        10'b1010110001: data <= 13'h1ff0; 
        10'b1010110010: data <= 13'h1ffa; 
        10'b1010110011: data <= 13'h1ffb; 
        10'b1010110100: data <= 13'h1ffe; 
        10'b1010110101: data <= 13'h1ffd; 
        10'b1010110110: data <= 13'h0002; 
        10'b1010110111: data <= 13'h1fff; 
        10'b1010111000: data <= 13'h1ffc; 
        10'b1010111001: data <= 13'h1fff; 
        10'b1010111010: data <= 13'h1ffd; 
        10'b1010111011: data <= 13'h1ffd; 
        10'b1010111100: data <= 13'h0004; 
        10'b1010111101: data <= 13'h1ffc; 
        10'b1010111110: data <= 13'h0001; 
        10'b1010111111: data <= 13'h1ffe; 
        10'b1011000000: data <= 13'h1ffd; 
        10'b1011000001: data <= 13'h1fff; 
        10'b1011000010: data <= 13'h0003; 
        10'b1011000011: data <= 13'h0000; 
        10'b1011000100: data <= 13'h1ffc; 
        10'b1011000101: data <= 13'h0002; 
        10'b1011000110: data <= 13'h1ffc; 
        10'b1011000111: data <= 13'h1fff; 
        10'b1011001000: data <= 13'h0000; 
        10'b1011001001: data <= 13'h1ffb; 
        10'b1011001010: data <= 13'h1ffd; 
        10'b1011001011: data <= 13'h1ffe; 
        10'b1011001100: data <= 13'h0000; 
        10'b1011001101: data <= 13'h1ffc; 
        10'b1011001110: data <= 13'h1ffe; 
        10'b1011001111: data <= 13'h1ffc; 
        10'b1011010000: data <= 13'h1ffd; 
        10'b1011010001: data <= 13'h0001; 
        10'b1011010010: data <= 13'h1ffe; 
        10'b1011010011: data <= 13'h0003; 
        10'b1011010100: data <= 13'h0004; 
        10'b1011010101: data <= 13'h0004; 
        10'b1011010110: data <= 13'h0000; 
        10'b1011010111: data <= 13'h0003; 
        10'b1011011000: data <= 13'h0004; 
        10'b1011011001: data <= 13'h0000; 
        10'b1011011010: data <= 13'h0001; 
        10'b1011011011: data <= 13'h1fff; 
        10'b1011011100: data <= 13'h1ffe; 
        10'b1011011101: data <= 13'h0004; 
        10'b1011011110: data <= 13'h0003; 
        10'b1011011111: data <= 13'h1ffe; 
        10'b1011100000: data <= 13'h1fff; 
        10'b1011100001: data <= 13'h0002; 
        10'b1011100010: data <= 13'h1ffe; 
        10'b1011100011: data <= 13'h0001; 
        10'b1011100100: data <= 13'h1ffe; 
        10'b1011100101: data <= 13'h0003; 
        10'b1011100110: data <= 13'h0003; 
        10'b1011100111: data <= 13'h1ffc; 
        10'b1011101000: data <= 13'h1ffd; 
        10'b1011101001: data <= 13'h0004; 
        10'b1011101010: data <= 13'h0003; 
        10'b1011101011: data <= 13'h1fff; 
        10'b1011101100: data <= 13'h0003; 
        10'b1011101101: data <= 13'h1fff; 
        10'b1011101110: data <= 13'h1fff; 
        10'b1011101111: data <= 13'h0002; 
        10'b1011110000: data <= 13'h0002; 
        10'b1011110001: data <= 13'h1fff; 
        10'b1011110010: data <= 13'h1ffe; 
        10'b1011110011: data <= 13'h1fff; 
        10'b1011110100: data <= 13'h0004; 
        10'b1011110101: data <= 13'h0000; 
        10'b1011110110: data <= 13'h0002; 
        10'b1011110111: data <= 13'h1ffe; 
        10'b1011111000: data <= 13'h0001; 
        10'b1011111001: data <= 13'h0000; 
        10'b1011111010: data <= 13'h0004; 
        10'b1011111011: data <= 13'h0001; 
        10'b1011111100: data <= 13'h1fff; 
        10'b1011111101: data <= 13'h1ffb; 
        10'b1011111110: data <= 13'h1ffd; 
        10'b1011111111: data <= 13'h0001; 
        10'b1100000000: data <= 13'h1ffc; 
        10'b1100000001: data <= 13'h1ffd; 
        10'b1100000010: data <= 13'h1ffd; 
        10'b1100000011: data <= 13'h1ffc; 
        10'b1100000100: data <= 13'h1ffd; 
        10'b1100000101: data <= 13'h1fff; 
        10'b1100000110: data <= 13'h1ffc; 
        10'b1100000111: data <= 13'h1ffd; 
        10'b1100001000: data <= 13'h1ffe; 
        10'b1100001001: data <= 13'h1ffe; 
        10'b1100001010: data <= 13'h0004; 
        10'b1100001011: data <= 13'h1ffc; 
        10'b1100001100: data <= 13'h1ffe; 
        10'b1100001101: data <= 13'h1ffc; 
        10'b1100001110: data <= 13'h1ffd; 
        10'b1100001111: data <= 13'h0001; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 8) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 14'h3ffd; 
        10'b0000000001: data <= 14'h0006; 
        10'b0000000010: data <= 14'h3ff9; 
        10'b0000000011: data <= 14'h3fff; 
        10'b0000000100: data <= 14'h0000; 
        10'b0000000101: data <= 14'h3fff; 
        10'b0000000110: data <= 14'h0003; 
        10'b0000000111: data <= 14'h0009; 
        10'b0000001000: data <= 14'h3ffa; 
        10'b0000001001: data <= 14'h3ffc; 
        10'b0000001010: data <= 14'h3ffc; 
        10'b0000001011: data <= 14'h3ffa; 
        10'b0000001100: data <= 14'h0003; 
        10'b0000001101: data <= 14'h0008; 
        10'b0000001110: data <= 14'h0005; 
        10'b0000001111: data <= 14'h3ff8; 
        10'b0000010000: data <= 14'h3fff; 
        10'b0000010001: data <= 14'h0009; 
        10'b0000010010: data <= 14'h0002; 
        10'b0000010011: data <= 14'h3fff; 
        10'b0000010100: data <= 14'h3ff9; 
        10'b0000010101: data <= 14'h3ffb; 
        10'b0000010110: data <= 14'h0002; 
        10'b0000010111: data <= 14'h0008; 
        10'b0000011000: data <= 14'h0004; 
        10'b0000011001: data <= 14'h0005; 
        10'b0000011010: data <= 14'h3ff9; 
        10'b0000011011: data <= 14'h3ff9; 
        10'b0000011100: data <= 14'h0006; 
        10'b0000011101: data <= 14'h0005; 
        10'b0000011110: data <= 14'h0006; 
        10'b0000011111: data <= 14'h3ffe; 
        10'b0000100000: data <= 14'h3ff8; 
        10'b0000100001: data <= 14'h3ffb; 
        10'b0000100010: data <= 14'h0004; 
        10'b0000100011: data <= 14'h000d; 
        10'b0000100100: data <= 14'h0009; 
        10'b0000100101: data <= 14'h0003; 
        10'b0000100110: data <= 14'h000b; 
        10'b0000100111: data <= 14'h000c; 
        10'b0000101000: data <= 14'h000d; 
        10'b0000101001: data <= 14'h000c; 
        10'b0000101010: data <= 14'h0007; 
        10'b0000101011: data <= 14'h0008; 
        10'b0000101100: data <= 14'h3ff8; 
        10'b0000101101: data <= 14'h0008; 
        10'b0000101110: data <= 14'h000a; 
        10'b0000101111: data <= 14'h0006; 
        10'b0000110000: data <= 14'h3ffe; 
        10'b0000110001: data <= 14'h3ffb; 
        10'b0000110010: data <= 14'h000b; 
        10'b0000110011: data <= 14'h0008; 
        10'b0000110100: data <= 14'h3ffd; 
        10'b0000110101: data <= 14'h0009; 
        10'b0000110110: data <= 14'h3ffe; 
        10'b0000110111: data <= 14'h0007; 
        10'b0000111000: data <= 14'h3ffb; 
        10'b0000111001: data <= 14'h3ffa; 
        10'b0000111010: data <= 14'h3ff8; 
        10'b0000111011: data <= 14'h3fff; 
        10'b0000111100: data <= 14'h0005; 
        10'b0000111101: data <= 14'h0003; 
        10'b0000111110: data <= 14'h0005; 
        10'b0000111111: data <= 14'h000d; 
        10'b0001000000: data <= 14'h0009; 
        10'b0001000001: data <= 14'h0014; 
        10'b0001000010: data <= 14'h0019; 
        10'b0001000011: data <= 14'h001c; 
        10'b0001000100: data <= 14'h001c; 
        10'b0001000101: data <= 14'h001e; 
        10'b0001000110: data <= 14'h000f; 
        10'b0001000111: data <= 14'h000b; 
        10'b0001001000: data <= 14'h0019; 
        10'b0001001001: data <= 14'h000b; 
        10'b0001001010: data <= 14'h000b; 
        10'b0001001011: data <= 14'h000c; 
        10'b0001001100: data <= 14'h000b; 
        10'b0001001101: data <= 14'h0006; 
        10'b0001001110: data <= 14'h0008; 
        10'b0001001111: data <= 14'h0001; 
        10'b0001010000: data <= 14'h0004; 
        10'b0001010001: data <= 14'h3ffe; 
        10'b0001010010: data <= 14'h3ff8; 
        10'b0001010011: data <= 14'h0003; 
        10'b0001010100: data <= 14'h3ff9; 
        10'b0001010101: data <= 14'h0001; 
        10'b0001010110: data <= 14'h0007; 
        10'b0001010111: data <= 14'h0004; 
        10'b0001011000: data <= 14'h0009; 
        10'b0001011001: data <= 14'h3ff8; 
        10'b0001011010: data <= 14'h000a; 
        10'b0001011011: data <= 14'h000b; 
        10'b0001011100: data <= 14'h000d; 
        10'b0001011101: data <= 14'h0019; 
        10'b0001011110: data <= 14'h0016; 
        10'b0001011111: data <= 14'h001c; 
        10'b0001100000: data <= 14'h001b; 
        10'b0001100001: data <= 14'h001a; 
        10'b0001100010: data <= 14'h0027; 
        10'b0001100011: data <= 14'h0025; 
        10'b0001100100: data <= 14'h0017; 
        10'b0001100101: data <= 14'h001d; 
        10'b0001100110: data <= 14'h002e; 
        10'b0001100111: data <= 14'h002e; 
        10'b0001101000: data <= 14'h0031; 
        10'b0001101001: data <= 14'h002c; 
        10'b0001101010: data <= 14'h002c; 
        10'b0001101011: data <= 14'h001a; 
        10'b0001101100: data <= 14'h0017; 
        10'b0001101101: data <= 14'h0006; 
        10'b0001101110: data <= 14'h3ffc; 
        10'b0001101111: data <= 14'h0005; 
        10'b0001110000: data <= 14'h0001; 
        10'b0001110001: data <= 14'h3ffe; 
        10'b0001110010: data <= 14'h3fff; 
        10'b0001110011: data <= 14'h0008; 
        10'b0001110100: data <= 14'h0007; 
        10'b0001110101: data <= 14'h0002; 
        10'b0001110110: data <= 14'h0002; 
        10'b0001110111: data <= 14'h0010; 
        10'b0001111000: data <= 14'h3ffe; 
        10'b0001111001: data <= 14'h3ffd; 
        10'b0001111010: data <= 14'h000f; 
        10'b0001111011: data <= 14'h0006; 
        10'b0001111100: data <= 14'h0007; 
        10'b0001111101: data <= 14'h0003; 
        10'b0001111110: data <= 14'h0006; 
        10'b0001111111: data <= 14'h0009; 
        10'b0010000000: data <= 14'h001f; 
        10'b0010000001: data <= 14'h001f; 
        10'b0010000010: data <= 14'h0030; 
        10'b0010000011: data <= 14'h0031; 
        10'b0010000100: data <= 14'h003d; 
        10'b0010000101: data <= 14'h0044; 
        10'b0010000110: data <= 14'h003a; 
        10'b0010000111: data <= 14'h0027; 
        10'b0010001000: data <= 14'h0006; 
        10'b0010001001: data <= 14'h000a; 
        10'b0010001010: data <= 14'h0001; 
        10'b0010001011: data <= 14'h0000; 
        10'b0010001100: data <= 14'h0002; 
        10'b0010001101: data <= 14'h0005; 
        10'b0010001110: data <= 14'h0003; 
        10'b0010001111: data <= 14'h3ffc; 
        10'b0010010000: data <= 14'h3ffa; 
        10'b0010010001: data <= 14'h3fff; 
        10'b0010010010: data <= 14'h3ffb; 
        10'b0010010011: data <= 14'h3ff5; 
        10'b0010010100: data <= 14'h0008; 
        10'b0010010101: data <= 14'h3ff6; 
        10'b0010010110: data <= 14'h0004; 
        10'b0010010111: data <= 14'h3fdc; 
        10'b0010011000: data <= 14'h3fed; 
        10'b0010011001: data <= 14'h3ff3; 
        10'b0010011010: data <= 14'h3ffb; 
        10'b0010011011: data <= 14'h3fef; 
        10'b0010011100: data <= 14'h3fef; 
        10'b0010011101: data <= 14'h0003; 
        10'b0010011110: data <= 14'h0017; 
        10'b0010011111: data <= 14'h002b; 
        10'b0010100000: data <= 14'h0025; 
        10'b0010100001: data <= 14'h0021; 
        10'b0010100010: data <= 14'h001a; 
        10'b0010100011: data <= 14'h0012; 
        10'b0010100100: data <= 14'h3ffe; 
        10'b0010100101: data <= 14'h0001; 
        10'b0010100110: data <= 14'h3ff7; 
        10'b0010100111: data <= 14'h0009; 
        10'b0010101000: data <= 14'h3fff; 
        10'b0010101001: data <= 14'h0008; 
        10'b0010101010: data <= 14'h0007; 
        10'b0010101011: data <= 14'h3ff7; 
        10'b0010101100: data <= 14'h0003; 
        10'b0010101101: data <= 14'h3fff; 
        10'b0010101110: data <= 14'h0003; 
        10'b0010101111: data <= 14'h0000; 
        10'b0010110000: data <= 14'h3ff3; 
        10'b0010110001: data <= 14'h3ff0; 
        10'b0010110010: data <= 14'h3fd7; 
        10'b0010110011: data <= 14'h3fca; 
        10'b0010110100: data <= 14'h3fe1; 
        10'b0010110101: data <= 14'h3fc3; 
        10'b0010110110: data <= 14'h3fe5; 
        10'b0010110111: data <= 14'h3fec; 
        10'b0010111000: data <= 14'h3fe4; 
        10'b0010111001: data <= 14'h3fe7; 
        10'b0010111010: data <= 14'h3ff9; 
        10'b0010111011: data <= 14'h3fef; 
        10'b0010111100: data <= 14'h3fe5; 
        10'b0010111101: data <= 14'h3fe6; 
        10'b0010111110: data <= 14'h3fd8; 
        10'b0010111111: data <= 14'h3fe6; 
        10'b0011000000: data <= 14'h3fea; 
        10'b0011000001: data <= 14'h3fe9; 
        10'b0011000010: data <= 14'h3ffd; 
        10'b0011000011: data <= 14'h0007; 
        10'b0011000100: data <= 14'h0003; 
        10'b0011000101: data <= 14'h0004; 
        10'b0011000110: data <= 14'h0000; 
        10'b0011000111: data <= 14'h3fff; 
        10'b0011001000: data <= 14'h0001; 
        10'b0011001001: data <= 14'h3ff8; 
        10'b0011001010: data <= 14'h3ff0; 
        10'b0011001011: data <= 14'h3ffd; 
        10'b0011001100: data <= 14'h3fe9; 
        10'b0011001101: data <= 14'h3fe4; 
        10'b0011001110: data <= 14'h3fd7; 
        10'b0011001111: data <= 14'h3fdf; 
        10'b0011010000: data <= 14'h3fc6; 
        10'b0011010001: data <= 14'h3fbe; 
        10'b0011010010: data <= 14'h3fde; 
        10'b0011010011: data <= 14'h3fdf; 
        10'b0011010100: data <= 14'h3fcd; 
        10'b0011010101: data <= 14'h3fd0; 
        10'b0011010110: data <= 14'h3fc4; 
        10'b0011010111: data <= 14'h3faf; 
        10'b0011011000: data <= 14'h3fad; 
        10'b0011011001: data <= 14'h3fbb; 
        10'b0011011010: data <= 14'h3fb7; 
        10'b0011011011: data <= 14'h3fc7; 
        10'b0011011100: data <= 14'h3fea; 
        10'b0011011101: data <= 14'h3fec; 
        10'b0011011110: data <= 14'h3ff8; 
        10'b0011011111: data <= 14'h3ffa; 
        10'b0011100000: data <= 14'h3ffd; 
        10'b0011100001: data <= 14'h3ffe; 
        10'b0011100010: data <= 14'h0009; 
        10'b0011100011: data <= 14'h3ff5; 
        10'b0011100100: data <= 14'h3ff7; 
        10'b0011100101: data <= 14'h3ff4; 
        10'b0011100110: data <= 14'h3fe1; 
        10'b0011100111: data <= 14'h3ff9; 
        10'b0011101000: data <= 14'h3ff4; 
        10'b0011101001: data <= 14'h3fdf; 
        10'b0011101010: data <= 14'h3fda; 
        10'b0011101011: data <= 14'h3fd4; 
        10'b0011101100: data <= 14'h3fcb; 
        10'b0011101101: data <= 14'h3fc3; 
        10'b0011101110: data <= 14'h3fc5; 
        10'b0011101111: data <= 14'h3fc1; 
        10'b0011110000: data <= 14'h3fb5; 
        10'b0011110001: data <= 14'h3fa9; 
        10'b0011110010: data <= 14'h3f86; 
        10'b0011110011: data <= 14'h3f8e; 
        10'b0011110100: data <= 14'h3f9a; 
        10'b0011110101: data <= 14'h3f9b; 
        10'b0011110110: data <= 14'h3fb9; 
        10'b0011110111: data <= 14'h3fc2; 
        10'b0011111000: data <= 14'h3fd9; 
        10'b0011111001: data <= 14'h3fe8; 
        10'b0011111010: data <= 14'h3fee; 
        10'b0011111011: data <= 14'h0003; 
        10'b0011111100: data <= 14'h3fff; 
        10'b0011111101: data <= 14'h3ff9; 
        10'b0011111110: data <= 14'h3ffc; 
        10'b0011111111: data <= 14'h3ff8; 
        10'b0100000000: data <= 14'h0000; 
        10'b0100000001: data <= 14'h3ff9; 
        10'b0100000010: data <= 14'h3ff5; 
        10'b0100000011: data <= 14'h3ffa; 
        10'b0100000100: data <= 14'h0007; 
        10'b0100000101: data <= 14'h3fec; 
        10'b0100000110: data <= 14'h3fdb; 
        10'b0100000111: data <= 14'h3fe3; 
        10'b0100001000: data <= 14'h3fee; 
        10'b0100001001: data <= 14'h3fdd; 
        10'b0100001010: data <= 14'h3fe0; 
        10'b0100001011: data <= 14'h3fba; 
        10'b0100001100: data <= 14'h3faf; 
        10'b0100001101: data <= 14'h3f8b; 
        10'b0100001110: data <= 14'h3f83; 
        10'b0100001111: data <= 14'h3f9a; 
        10'b0100010000: data <= 14'h3fac; 
        10'b0100010001: data <= 14'h3fbd; 
        10'b0100010010: data <= 14'h3fb3; 
        10'b0100010011: data <= 14'h3fce; 
        10'b0100010100: data <= 14'h3fda; 
        10'b0100010101: data <= 14'h3fe4; 
        10'b0100010110: data <= 14'h3ff4; 
        10'b0100010111: data <= 14'h0006; 
        10'b0100011000: data <= 14'h3ffa; 
        10'b0100011001: data <= 14'h0008; 
        10'b0100011010: data <= 14'h0005; 
        10'b0100011011: data <= 14'h3ff7; 
        10'b0100011100: data <= 14'h3ff3; 
        10'b0100011101: data <= 14'h0003; 
        10'b0100011110: data <= 14'h000b; 
        10'b0100011111: data <= 14'h000a; 
        10'b0100100000: data <= 14'h0026; 
        10'b0100100001: data <= 14'h3fff; 
        10'b0100100010: data <= 14'h0008; 
        10'b0100100011: data <= 14'h0003; 
        10'b0100100100: data <= 14'h3fe9; 
        10'b0100100101: data <= 14'h3ff0; 
        10'b0100100110: data <= 14'h3fde; 
        10'b0100100111: data <= 14'h3fb8; 
        10'b0100101000: data <= 14'h3fb7; 
        10'b0100101001: data <= 14'h3faa; 
        10'b0100101010: data <= 14'h3fa7; 
        10'b0100101011: data <= 14'h3fb9; 
        10'b0100101100: data <= 14'h3fd0; 
        10'b0100101101: data <= 14'h3fdd; 
        10'b0100101110: data <= 14'h3fd2; 
        10'b0100101111: data <= 14'h3ffb; 
        10'b0100110000: data <= 14'h3fe2; 
        10'b0100110001: data <= 14'h3feb; 
        10'b0100110010: data <= 14'h3ffa; 
        10'b0100110011: data <= 14'h3ffd; 
        10'b0100110100: data <= 14'h3ffb; 
        10'b0100110101: data <= 14'h0003; 
        10'b0100110110: data <= 14'h3ffb; 
        10'b0100110111: data <= 14'h3fff; 
        10'b0100111000: data <= 14'h3ffb; 
        10'b0100111001: data <= 14'h0001; 
        10'b0100111010: data <= 14'h3ffd; 
        10'b0100111011: data <= 14'h0020; 
        10'b0100111100: data <= 14'h0017; 
        10'b0100111101: data <= 14'h000b; 
        10'b0100111110: data <= 14'h000e; 
        10'b0100111111: data <= 14'h000a; 
        10'b0101000000: data <= 14'h000a; 
        10'b0101000001: data <= 14'h0002; 
        10'b0101000010: data <= 14'h3fef; 
        10'b0101000011: data <= 14'h3fc7; 
        10'b0101000100: data <= 14'h3fca; 
        10'b0101000101: data <= 14'h3fd2; 
        10'b0101000110: data <= 14'h3fd2; 
        10'b0101000111: data <= 14'h3fdc; 
        10'b0101001000: data <= 14'h3fef; 
        10'b0101001001: data <= 14'h0006; 
        10'b0101001010: data <= 14'h0016; 
        10'b0101001011: data <= 14'h0022; 
        10'b0101001100: data <= 14'h0000; 
        10'b0101001101: data <= 14'h3fee; 
        10'b0101001110: data <= 14'h3ff8; 
        10'b0101001111: data <= 14'h3ffd; 
        10'b0101010000: data <= 14'h3ffb; 
        10'b0101010001: data <= 14'h3ffd; 
        10'b0101010010: data <= 14'h3ff8; 
        10'b0101010011: data <= 14'h3ffc; 
        10'b0101010100: data <= 14'h0005; 
        10'b0101010101: data <= 14'h000f; 
        10'b0101010110: data <= 14'h0017; 
        10'b0101010111: data <= 14'h001e; 
        10'b0101011000: data <= 14'h000e; 
        10'b0101011001: data <= 14'h0013; 
        10'b0101011010: data <= 14'h000e; 
        10'b0101011011: data <= 14'h0024; 
        10'b0101011100: data <= 14'h0023; 
        10'b0101011101: data <= 14'h0019; 
        10'b0101011110: data <= 14'h3feb; 
        10'b0101011111: data <= 14'h3fda; 
        10'b0101100000: data <= 14'h3ffe; 
        10'b0101100001: data <= 14'h3ffc; 
        10'b0101100010: data <= 14'h3fdb; 
        10'b0101100011: data <= 14'h3fdc; 
        10'b0101100100: data <= 14'h3ffc; 
        10'b0101100101: data <= 14'h0014; 
        10'b0101100110: data <= 14'h0031; 
        10'b0101100111: data <= 14'h0057; 
        10'b0101101000: data <= 14'h002f; 
        10'b0101101001: data <= 14'h3ff3; 
        10'b0101101010: data <= 14'h3ff1; 
        10'b0101101011: data <= 14'h3ffb; 
        10'b0101101100: data <= 14'h3ffb; 
        10'b0101101101: data <= 14'h0008; 
        10'b0101101110: data <= 14'h0006; 
        10'b0101101111: data <= 14'h3ff7; 
        10'b0101110000: data <= 14'h3ff4; 
        10'b0101110001: data <= 14'h0005; 
        10'b0101110010: data <= 14'h0026; 
        10'b0101110011: data <= 14'h0014; 
        10'b0101110100: data <= 14'h0011; 
        10'b0101110101: data <= 14'h0009; 
        10'b0101110110: data <= 14'h0025; 
        10'b0101110111: data <= 14'h001f; 
        10'b0101111000: data <= 14'h001c; 
        10'b0101111001: data <= 14'h0005; 
        10'b0101111010: data <= 14'h3ffb; 
        10'b0101111011: data <= 14'h3fff; 
        10'b0101111100: data <= 14'h0003; 
        10'b0101111101: data <= 14'h3ff8; 
        10'b0101111110: data <= 14'h3fdf; 
        10'b0101111111: data <= 14'h3ffc; 
        10'b0110000000: data <= 14'h3ff0; 
        10'b0110000001: data <= 14'h001a; 
        10'b0110000010: data <= 14'h0044; 
        10'b0110000011: data <= 14'h006b; 
        10'b0110000100: data <= 14'h003a; 
        10'b0110000101: data <= 14'h3ffb; 
        10'b0110000110: data <= 14'h0000; 
        10'b0110000111: data <= 14'h0005; 
        10'b0110001000: data <= 14'h3ffc; 
        10'b0110001001: data <= 14'h0001; 
        10'b0110001010: data <= 14'h0006; 
        10'b0110001011: data <= 14'h0000; 
        10'b0110001100: data <= 14'h3ff3; 
        10'b0110001101: data <= 14'h000e; 
        10'b0110001110: data <= 14'h0023; 
        10'b0110001111: data <= 14'h001e; 
        10'b0110010000: data <= 14'h0029; 
        10'b0110010001: data <= 14'h0026; 
        10'b0110010010: data <= 14'h002a; 
        10'b0110010011: data <= 14'h002d; 
        10'b0110010100: data <= 14'h000f; 
        10'b0110010101: data <= 14'h3fea; 
        10'b0110010110: data <= 14'h0001; 
        10'b0110010111: data <= 14'h0012; 
        10'b0110011000: data <= 14'h0009; 
        10'b0110011001: data <= 14'h3ff2; 
        10'b0110011010: data <= 14'h3ff2; 
        10'b0110011011: data <= 14'h3ffe; 
        10'b0110011100: data <= 14'h001d; 
        10'b0110011101: data <= 14'h001d; 
        10'b0110011110: data <= 14'h004d; 
        10'b0110011111: data <= 14'h0059; 
        10'b0110100000: data <= 14'h003b; 
        10'b0110100001: data <= 14'h3fff; 
        10'b0110100010: data <= 14'h3fef; 
        10'b0110100011: data <= 14'h3ff8; 
        10'b0110100100: data <= 14'h0006; 
        10'b0110100101: data <= 14'h3ffd; 
        10'b0110100110: data <= 14'h0001; 
        10'b0110100111: data <= 14'h3ff9; 
        10'b0110101000: data <= 14'h3fe8; 
        10'b0110101001: data <= 14'h3ffd; 
        10'b0110101010: data <= 14'h0024; 
        10'b0110101011: data <= 14'h0030; 
        10'b0110101100: data <= 14'h001f; 
        10'b0110101101: data <= 14'h0030; 
        10'b0110101110: data <= 14'h003d; 
        10'b0110101111: data <= 14'h004b; 
        10'b0110110000: data <= 14'h0013; 
        10'b0110110001: data <= 14'h3ffb; 
        10'b0110110010: data <= 14'h001d; 
        10'b0110110011: data <= 14'h001a; 
        10'b0110110100: data <= 14'h0004; 
        10'b0110110101: data <= 14'h3ff2; 
        10'b0110110110: data <= 14'h0003; 
        10'b0110110111: data <= 14'h000f; 
        10'b0110111000: data <= 14'h0022; 
        10'b0110111001: data <= 14'h002f; 
        10'b0110111010: data <= 14'h002b; 
        10'b0110111011: data <= 14'h0036; 
        10'b0110111100: data <= 14'h001d; 
        10'b0110111101: data <= 14'h3ff1; 
        10'b0110111110: data <= 14'h3ff7; 
        10'b0110111111: data <= 14'h3ff7; 
        10'b0111000000: data <= 14'h0002; 
        10'b0111000001: data <= 14'h3ff9; 
        10'b0111000010: data <= 14'h3ff9; 
        10'b0111000011: data <= 14'h3ff8; 
        10'b0111000100: data <= 14'h3fe0; 
        10'b0111000101: data <= 14'h3fef; 
        10'b0111000110: data <= 14'h0035; 
        10'b0111000111: data <= 14'h0037; 
        10'b0111001000: data <= 14'h0024; 
        10'b0111001001: data <= 14'h0038; 
        10'b0111001010: data <= 14'h005f; 
        10'b0111001011: data <= 14'h005e; 
        10'b0111001100: data <= 14'h001d; 
        10'b0111001101: data <= 14'h0011; 
        10'b0111001110: data <= 14'h0029; 
        10'b0111001111: data <= 14'h0016; 
        10'b0111010000: data <= 14'h3ff5; 
        10'b0111010001: data <= 14'h3fea; 
        10'b0111010010: data <= 14'h0008; 
        10'b0111010011: data <= 14'h0018; 
        10'b0111010100: data <= 14'h000b; 
        10'b0111010101: data <= 14'h0000; 
        10'b0111010110: data <= 14'h0016; 
        10'b0111010111: data <= 14'h000d; 
        10'b0111011000: data <= 14'h3ffa; 
        10'b0111011001: data <= 14'h3fef; 
        10'b0111011010: data <= 14'h3ff5; 
        10'b0111011011: data <= 14'h3fff; 
        10'b0111011100: data <= 14'h0002; 
        10'b0111011101: data <= 14'h0005; 
        10'b0111011110: data <= 14'h0007; 
        10'b0111011111: data <= 14'h3fff; 
        10'b0111100000: data <= 14'h3fd2; 
        10'b0111100001: data <= 14'h3fe8; 
        10'b0111100010: data <= 14'h0016; 
        10'b0111100011: data <= 14'h002a; 
        10'b0111100100: data <= 14'h0030; 
        10'b0111100101: data <= 14'h003d; 
        10'b0111100110: data <= 14'h0069; 
        10'b0111100111: data <= 14'h006b; 
        10'b0111101000: data <= 14'h0037; 
        10'b0111101001: data <= 14'h001f; 
        10'b0111101010: data <= 14'h001f; 
        10'b0111101011: data <= 14'h0014; 
        10'b0111101100: data <= 14'h0000; 
        10'b0111101101: data <= 14'h0006; 
        10'b0111101110: data <= 14'h002c; 
        10'b0111101111: data <= 14'h000f; 
        10'b0111110000: data <= 14'h0006; 
        10'b0111110001: data <= 14'h3ff5; 
        10'b0111110010: data <= 14'h000a; 
        10'b0111110011: data <= 14'h3ffe; 
        10'b0111110100: data <= 14'h3ff4; 
        10'b0111110101: data <= 14'h3fe8; 
        10'b0111110110: data <= 14'h3ffd; 
        10'b0111110111: data <= 14'h0004; 
        10'b0111111000: data <= 14'h3ffc; 
        10'b0111111001: data <= 14'h3ffb; 
        10'b0111111010: data <= 14'h0000; 
        10'b0111111011: data <= 14'h3ff3; 
        10'b0111111100: data <= 14'h3fd5; 
        10'b0111111101: data <= 14'h3fd6; 
        10'b0111111110: data <= 14'h3fec; 
        10'b0111111111: data <= 14'h001d; 
        10'b1000000000: data <= 14'h002f; 
        10'b1000000001: data <= 14'h002b; 
        10'b1000000010: data <= 14'h004a; 
        10'b1000000011: data <= 14'h005b; 
        10'b1000000100: data <= 14'h006b; 
        10'b1000000101: data <= 14'h0032; 
        10'b1000000110: data <= 14'h000d; 
        10'b1000000111: data <= 14'h001c; 
        10'b1000001000: data <= 14'h0030; 
        10'b1000001001: data <= 14'h001f; 
        10'b1000001010: data <= 14'h0027; 
        10'b1000001011: data <= 14'h0014; 
        10'b1000001100: data <= 14'h0003; 
        10'b1000001101: data <= 14'h0007; 
        10'b1000001110: data <= 14'h0007; 
        10'b1000001111: data <= 14'h3ffc; 
        10'b1000010000: data <= 14'h3ff1; 
        10'b1000010001: data <= 14'h3ff5; 
        10'b1000010010: data <= 14'h3ff7; 
        10'b1000010011: data <= 14'h3ff7; 
        10'b1000010100: data <= 14'h0002; 
        10'b1000010101: data <= 14'h3ffa; 
        10'b1000010110: data <= 14'h0004; 
        10'b1000010111: data <= 14'h3fef; 
        10'b1000011000: data <= 14'h3fe4; 
        10'b1000011001: data <= 14'h3fd3; 
        10'b1000011010: data <= 14'h3fdd; 
        10'b1000011011: data <= 14'h0002; 
        10'b1000011100: data <= 14'h001e; 
        10'b1000011101: data <= 14'h0030; 
        10'b1000011110: data <= 14'h0040; 
        10'b1000011111: data <= 14'h0065; 
        10'b1000100000: data <= 14'h0072; 
        10'b1000100001: data <= 14'h003b; 
        10'b1000100010: data <= 14'h0034; 
        10'b1000100011: data <= 14'h0037; 
        10'b1000100100: data <= 14'h0027; 
        10'b1000100101: data <= 14'h0020; 
        10'b1000100110: data <= 14'h0032; 
        10'b1000100111: data <= 14'h0022; 
        10'b1000101000: data <= 14'h0016; 
        10'b1000101001: data <= 14'h0005; 
        10'b1000101010: data <= 14'h3ff8; 
        10'b1000101011: data <= 14'h3ff6; 
        10'b1000101100: data <= 14'h3ff6; 
        10'b1000101101: data <= 14'h3ffe; 
        10'b1000101110: data <= 14'h3ffb; 
        10'b1000101111: data <= 14'h0007; 
        10'b1000110000: data <= 14'h3ffc; 
        10'b1000110001: data <= 14'h3ff9; 
        10'b1000110010: data <= 14'h3ffe; 
        10'b1000110011: data <= 14'h3ff8; 
        10'b1000110100: data <= 14'h3fdc; 
        10'b1000110101: data <= 14'h3fd6; 
        10'b1000110110: data <= 14'h3fdb; 
        10'b1000110111: data <= 14'h3ff1; 
        10'b1000111000: data <= 14'h000a; 
        10'b1000111001: data <= 14'h0020; 
        10'b1000111010: data <= 14'h0035; 
        10'b1000111011: data <= 14'h0023; 
        10'b1000111100: data <= 14'h0045; 
        10'b1000111101: data <= 14'h0053; 
        10'b1000111110: data <= 14'h0062; 
        10'b1000111111: data <= 14'h0054; 
        10'b1001000000: data <= 14'h002d; 
        10'b1001000001: data <= 14'h001d; 
        10'b1001000010: data <= 14'h0038; 
        10'b1001000011: data <= 14'h0028; 
        10'b1001000100: data <= 14'h001b; 
        10'b1001000101: data <= 14'h3ffa; 
        10'b1001000110: data <= 14'h3feb; 
        10'b1001000111: data <= 14'h0001; 
        10'b1001001000: data <= 14'h3ffb; 
        10'b1001001001: data <= 14'h3ffd; 
        10'b1001001010: data <= 14'h3ffa; 
        10'b1001001011: data <= 14'h0001; 
        10'b1001001100: data <= 14'h3fff; 
        10'b1001001101: data <= 14'h0001; 
        10'b1001001110: data <= 14'h0003; 
        10'b1001001111: data <= 14'h3ffd; 
        10'b1001010000: data <= 14'h3ff3; 
        10'b1001010001: data <= 14'h3fe3; 
        10'b1001010010: data <= 14'h3fce; 
        10'b1001010011: data <= 14'h3fea; 
        10'b1001010100: data <= 14'h3ff3; 
        10'b1001010101: data <= 14'h0018; 
        10'b1001010110: data <= 14'h002c; 
        10'b1001010111: data <= 14'h003e; 
        10'b1001011000: data <= 14'h0050; 
        10'b1001011001: data <= 14'h0051; 
        10'b1001011010: data <= 14'h0044; 
        10'b1001011011: data <= 14'h003b; 
        10'b1001011100: data <= 14'h0025; 
        10'b1001011101: data <= 14'h0032; 
        10'b1001011110: data <= 14'h002f; 
        10'b1001011111: data <= 14'h001e; 
        10'b1001100000: data <= 14'h0004; 
        10'b1001100001: data <= 14'h3ff0; 
        10'b1001100010: data <= 14'h3fea; 
        10'b1001100011: data <= 14'h3ff3; 
        10'b1001100100: data <= 14'h0001; 
        10'b1001100101: data <= 14'h3ff8; 
        10'b1001100110: data <= 14'h3ffe; 
        10'b1001100111: data <= 14'h3ffb; 
        10'b1001101000: data <= 14'h3ffb; 
        10'b1001101001: data <= 14'h3fff; 
        10'b1001101010: data <= 14'h0008; 
        10'b1001101011: data <= 14'h0002; 
        10'b1001101100: data <= 14'h3ffb; 
        10'b1001101101: data <= 14'h3fe7; 
        10'b1001101110: data <= 14'h3fe2; 
        10'b1001101111: data <= 14'h3fd7; 
        10'b1001110000: data <= 14'h3fe5; 
        10'b1001110001: data <= 14'h3ff4; 
        10'b1001110010: data <= 14'h3ff6; 
        10'b1001110011: data <= 14'h0005; 
        10'b1001110100: data <= 14'h0017; 
        10'b1001110101: data <= 14'h000a; 
        10'b1001110110: data <= 14'h0009; 
        10'b1001110111: data <= 14'h0019; 
        10'b1001111000: data <= 14'h0013; 
        10'b1001111001: data <= 14'h0000; 
        10'b1001111010: data <= 14'h3ffa; 
        10'b1001111011: data <= 14'h3fe4; 
        10'b1001111100: data <= 14'h3fe5; 
        10'b1001111101: data <= 14'h3fe9; 
        10'b1001111110: data <= 14'h3feb; 
        10'b1001111111: data <= 14'h3ffe; 
        10'b1010000000: data <= 14'h3ffc; 
        10'b1010000001: data <= 14'h3ff8; 
        10'b1010000010: data <= 14'h0009; 
        10'b1010000011: data <= 14'h0003; 
        10'b1010000100: data <= 14'h0007; 
        10'b1010000101: data <= 14'h3ffd; 
        10'b1010000110: data <= 14'h3ffc; 
        10'b1010000111: data <= 14'h0001; 
        10'b1010001000: data <= 14'h0002; 
        10'b1010001001: data <= 14'h3ff5; 
        10'b1010001010: data <= 14'h3ff0; 
        10'b1010001011: data <= 14'h3fdc; 
        10'b1010001100: data <= 14'h3fd2; 
        10'b1010001101: data <= 14'h3fbe; 
        10'b1010001110: data <= 14'h3fbf; 
        10'b1010001111: data <= 14'h3fb4; 
        10'b1010010000: data <= 14'h3fd1; 
        10'b1010010001: data <= 14'h3fdb; 
        10'b1010010010: data <= 14'h3fe3; 
        10'b1010010011: data <= 14'h3fd5; 
        10'b1010010100: data <= 14'h3fc8; 
        10'b1010010101: data <= 14'h3fc0; 
        10'b1010010110: data <= 14'h3fce; 
        10'b1010010111: data <= 14'h3fe9; 
        10'b1010011000: data <= 14'h3fe9; 
        10'b1010011001: data <= 14'h3fec; 
        10'b1010011010: data <= 14'h3ff9; 
        10'b1010011011: data <= 14'h0001; 
        10'b1010011100: data <= 14'h3ff7; 
        10'b1010011101: data <= 14'h3ff9; 
        10'b1010011110: data <= 14'h3ffd; 
        10'b1010011111: data <= 14'h3fff; 
        10'b1010100000: data <= 14'h0005; 
        10'b1010100001: data <= 14'h0004; 
        10'b1010100010: data <= 14'h0003; 
        10'b1010100011: data <= 14'h3ff8; 
        10'b1010100100: data <= 14'h3ffa; 
        10'b1010100101: data <= 14'h3ffd; 
        10'b1010100110: data <= 14'h3ff8; 
        10'b1010100111: data <= 14'h3ff3; 
        10'b1010101000: data <= 14'h3ff6; 
        10'b1010101001: data <= 14'h3ff0; 
        10'b1010101010: data <= 14'h3fe8; 
        10'b1010101011: data <= 14'h3fe2; 
        10'b1010101100: data <= 14'h3fdd; 
        10'b1010101101: data <= 14'h3fde; 
        10'b1010101110: data <= 14'h3fd8; 
        10'b1010101111: data <= 14'h3fd8; 
        10'b1010110000: data <= 14'h3fd6; 
        10'b1010110001: data <= 14'h3fe0; 
        10'b1010110010: data <= 14'h3ff5; 
        10'b1010110011: data <= 14'h3ff6; 
        10'b1010110100: data <= 14'h3ffc; 
        10'b1010110101: data <= 14'h3ffa; 
        10'b1010110110: data <= 14'h0004; 
        10'b1010110111: data <= 14'h3ffe; 
        10'b1010111000: data <= 14'h3ff8; 
        10'b1010111001: data <= 14'h3ffd; 
        10'b1010111010: data <= 14'h3ffa; 
        10'b1010111011: data <= 14'h3ffa; 
        10'b1010111100: data <= 14'h0008; 
        10'b1010111101: data <= 14'h3ff9; 
        10'b1010111110: data <= 14'h0002; 
        10'b1010111111: data <= 14'h3ffc; 
        10'b1011000000: data <= 14'h3ffa; 
        10'b1011000001: data <= 14'h3fff; 
        10'b1011000010: data <= 14'h0005; 
        10'b1011000011: data <= 14'h0000; 
        10'b1011000100: data <= 14'h3ff7; 
        10'b1011000101: data <= 14'h0003; 
        10'b1011000110: data <= 14'h3ff7; 
        10'b1011000111: data <= 14'h3fff; 
        10'b1011001000: data <= 14'h0000; 
        10'b1011001001: data <= 14'h3ff7; 
        10'b1011001010: data <= 14'h3ffb; 
        10'b1011001011: data <= 14'h3ffd; 
        10'b1011001100: data <= 14'h3fff; 
        10'b1011001101: data <= 14'h3ff8; 
        10'b1011001110: data <= 14'h3ffb; 
        10'b1011001111: data <= 14'h3ff7; 
        10'b1011010000: data <= 14'h3ff9; 
        10'b1011010001: data <= 14'h0001; 
        10'b1011010010: data <= 14'h3ffd; 
        10'b1011010011: data <= 14'h0006; 
        10'b1011010100: data <= 14'h0009; 
        10'b1011010101: data <= 14'h0008; 
        10'b1011010110: data <= 14'h0000; 
        10'b1011010111: data <= 14'h0006; 
        10'b1011011000: data <= 14'h0008; 
        10'b1011011001: data <= 14'h0000; 
        10'b1011011010: data <= 14'h0002; 
        10'b1011011011: data <= 14'h3ffe; 
        10'b1011011100: data <= 14'h3ffb; 
        10'b1011011101: data <= 14'h0007; 
        10'b1011011110: data <= 14'h0005; 
        10'b1011011111: data <= 14'h3ffb; 
        10'b1011100000: data <= 14'h3ffd; 
        10'b1011100001: data <= 14'h0004; 
        10'b1011100010: data <= 14'h3ffd; 
        10'b1011100011: data <= 14'h0002; 
        10'b1011100100: data <= 14'h3ffc; 
        10'b1011100101: data <= 14'h0005; 
        10'b1011100110: data <= 14'h0006; 
        10'b1011100111: data <= 14'h3ff9; 
        10'b1011101000: data <= 14'h3ffb; 
        10'b1011101001: data <= 14'h0007; 
        10'b1011101010: data <= 14'h0006; 
        10'b1011101011: data <= 14'h3ffd; 
        10'b1011101100: data <= 14'h0005; 
        10'b1011101101: data <= 14'h3ffe; 
        10'b1011101110: data <= 14'h3ffe; 
        10'b1011101111: data <= 14'h0003; 
        10'b1011110000: data <= 14'h0004; 
        10'b1011110001: data <= 14'h3ffe; 
        10'b1011110010: data <= 14'h3ffc; 
        10'b1011110011: data <= 14'h3ffe; 
        10'b1011110100: data <= 14'h0008; 
        10'b1011110101: data <= 14'h0000; 
        10'b1011110110: data <= 14'h0005; 
        10'b1011110111: data <= 14'h3ffb; 
        10'b1011111000: data <= 14'h0003; 
        10'b1011111001: data <= 14'h0000; 
        10'b1011111010: data <= 14'h0008; 
        10'b1011111011: data <= 14'h0001; 
        10'b1011111100: data <= 14'h3fff; 
        10'b1011111101: data <= 14'h3ff7; 
        10'b1011111110: data <= 14'h3ffa; 
        10'b1011111111: data <= 14'h0003; 
        10'b1100000000: data <= 14'h3ff8; 
        10'b1100000001: data <= 14'h3ff9; 
        10'b1100000010: data <= 14'h3ffb; 
        10'b1100000011: data <= 14'h3ff8; 
        10'b1100000100: data <= 14'h3ffa; 
        10'b1100000101: data <= 14'h3ffd; 
        10'b1100000110: data <= 14'h3ff9; 
        10'b1100000111: data <= 14'h3ffa; 
        10'b1100001000: data <= 14'h3ffb; 
        10'b1100001001: data <= 14'h3ffc; 
        10'b1100001010: data <= 14'h0008; 
        10'b1100001011: data <= 14'h3ff9; 
        10'b1100001100: data <= 14'h3ffb; 
        10'b1100001101: data <= 14'h3ff9; 
        10'b1100001110: data <= 14'h3ffb; 
        10'b1100001111: data <= 14'h0001; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 9) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 15'h7ffa; 
        10'b0000000001: data <= 15'h000c; 
        10'b0000000010: data <= 15'h7ff3; 
        10'b0000000011: data <= 15'h7fff; 
        10'b0000000100: data <= 15'h0000; 
        10'b0000000101: data <= 15'h7ffe; 
        10'b0000000110: data <= 15'h0006; 
        10'b0000000111: data <= 15'h0012; 
        10'b0000001000: data <= 15'h7ff4; 
        10'b0000001001: data <= 15'h7ff8; 
        10'b0000001010: data <= 15'h7ff8; 
        10'b0000001011: data <= 15'h7ff4; 
        10'b0000001100: data <= 15'h0006; 
        10'b0000001101: data <= 15'h0011; 
        10'b0000001110: data <= 15'h0009; 
        10'b0000001111: data <= 15'h7ff1; 
        10'b0000010000: data <= 15'h7ffe; 
        10'b0000010001: data <= 15'h0012; 
        10'b0000010010: data <= 15'h0003; 
        10'b0000010011: data <= 15'h7ffe; 
        10'b0000010100: data <= 15'h7ff2; 
        10'b0000010101: data <= 15'h7ff7; 
        10'b0000010110: data <= 15'h0004; 
        10'b0000010111: data <= 15'h0010; 
        10'b0000011000: data <= 15'h0009; 
        10'b0000011001: data <= 15'h000b; 
        10'b0000011010: data <= 15'h7ff2; 
        10'b0000011011: data <= 15'h7ff2; 
        10'b0000011100: data <= 15'h000c; 
        10'b0000011101: data <= 15'h0009; 
        10'b0000011110: data <= 15'h000c; 
        10'b0000011111: data <= 15'h7ffd; 
        10'b0000100000: data <= 15'h7ff0; 
        10'b0000100001: data <= 15'h7ff6; 
        10'b0000100010: data <= 15'h0008; 
        10'b0000100011: data <= 15'h001b; 
        10'b0000100100: data <= 15'h0012; 
        10'b0000100101: data <= 15'h0005; 
        10'b0000100110: data <= 15'h0016; 
        10'b0000100111: data <= 15'h0018; 
        10'b0000101000: data <= 15'h0019; 
        10'b0000101001: data <= 15'h0018; 
        10'b0000101010: data <= 15'h000f; 
        10'b0000101011: data <= 15'h0010; 
        10'b0000101100: data <= 15'h7fef; 
        10'b0000101101: data <= 15'h000f; 
        10'b0000101110: data <= 15'h0015; 
        10'b0000101111: data <= 15'h000c; 
        10'b0000110000: data <= 15'h7ffd; 
        10'b0000110001: data <= 15'h7ff6; 
        10'b0000110010: data <= 15'h0016; 
        10'b0000110011: data <= 15'h0010; 
        10'b0000110100: data <= 15'h7ff9; 
        10'b0000110101: data <= 15'h0012; 
        10'b0000110110: data <= 15'h7ffd; 
        10'b0000110111: data <= 15'h000e; 
        10'b0000111000: data <= 15'h7ff5; 
        10'b0000111001: data <= 15'h7ff3; 
        10'b0000111010: data <= 15'h7ff0; 
        10'b0000111011: data <= 15'h7ffe; 
        10'b0000111100: data <= 15'h0009; 
        10'b0000111101: data <= 15'h0006; 
        10'b0000111110: data <= 15'h0009; 
        10'b0000111111: data <= 15'h001a; 
        10'b0001000000: data <= 15'h0013; 
        10'b0001000001: data <= 15'h0028; 
        10'b0001000010: data <= 15'h0032; 
        10'b0001000011: data <= 15'h0039; 
        10'b0001000100: data <= 15'h0039; 
        10'b0001000101: data <= 15'h003c; 
        10'b0001000110: data <= 15'h001e; 
        10'b0001000111: data <= 15'h0015; 
        10'b0001001000: data <= 15'h0032; 
        10'b0001001001: data <= 15'h0016; 
        10'b0001001010: data <= 15'h0015; 
        10'b0001001011: data <= 15'h0017; 
        10'b0001001100: data <= 15'h0017; 
        10'b0001001101: data <= 15'h000c; 
        10'b0001001110: data <= 15'h000f; 
        10'b0001001111: data <= 15'h0003; 
        10'b0001010000: data <= 15'h0008; 
        10'b0001010001: data <= 15'h7ffb; 
        10'b0001010010: data <= 15'h7fef; 
        10'b0001010011: data <= 15'h0005; 
        10'b0001010100: data <= 15'h7ff2; 
        10'b0001010101: data <= 15'h0002; 
        10'b0001010110: data <= 15'h000d; 
        10'b0001010111: data <= 15'h0008; 
        10'b0001011000: data <= 15'h0012; 
        10'b0001011001: data <= 15'h7ff1; 
        10'b0001011010: data <= 15'h0013; 
        10'b0001011011: data <= 15'h0015; 
        10'b0001011100: data <= 15'h0019; 
        10'b0001011101: data <= 15'h0033; 
        10'b0001011110: data <= 15'h002d; 
        10'b0001011111: data <= 15'h0038; 
        10'b0001100000: data <= 15'h0037; 
        10'b0001100001: data <= 15'h0035; 
        10'b0001100010: data <= 15'h004e; 
        10'b0001100011: data <= 15'h0049; 
        10'b0001100100: data <= 15'h002e; 
        10'b0001100101: data <= 15'h003a; 
        10'b0001100110: data <= 15'h005c; 
        10'b0001100111: data <= 15'h005c; 
        10'b0001101000: data <= 15'h0062; 
        10'b0001101001: data <= 15'h0057; 
        10'b0001101010: data <= 15'h0058; 
        10'b0001101011: data <= 15'h0033; 
        10'b0001101100: data <= 15'h002d; 
        10'b0001101101: data <= 15'h000b; 
        10'b0001101110: data <= 15'h7ff8; 
        10'b0001101111: data <= 15'h000a; 
        10'b0001110000: data <= 15'h0003; 
        10'b0001110001: data <= 15'h7ffd; 
        10'b0001110010: data <= 15'h7fff; 
        10'b0001110011: data <= 15'h0010; 
        10'b0001110100: data <= 15'h000d; 
        10'b0001110101: data <= 15'h0005; 
        10'b0001110110: data <= 15'h0005; 
        10'b0001110111: data <= 15'h001f; 
        10'b0001111000: data <= 15'h7ffc; 
        10'b0001111001: data <= 15'h7ff9; 
        10'b0001111010: data <= 15'h001e; 
        10'b0001111011: data <= 15'h000b; 
        10'b0001111100: data <= 15'h000e; 
        10'b0001111101: data <= 15'h0005; 
        10'b0001111110: data <= 15'h000c; 
        10'b0001111111: data <= 15'h0012; 
        10'b0010000000: data <= 15'h003e; 
        10'b0010000001: data <= 15'h003d; 
        10'b0010000010: data <= 15'h0060; 
        10'b0010000011: data <= 15'h0061; 
        10'b0010000100: data <= 15'h007b; 
        10'b0010000101: data <= 15'h0088; 
        10'b0010000110: data <= 15'h0075; 
        10'b0010000111: data <= 15'h004f; 
        10'b0010001000: data <= 15'h000b; 
        10'b0010001001: data <= 15'h0015; 
        10'b0010001010: data <= 15'h0003; 
        10'b0010001011: data <= 15'h0000; 
        10'b0010001100: data <= 15'h0003; 
        10'b0010001101: data <= 15'h000a; 
        10'b0010001110: data <= 15'h0005; 
        10'b0010001111: data <= 15'h7ff9; 
        10'b0010010000: data <= 15'h7ff3; 
        10'b0010010001: data <= 15'h7fff; 
        10'b0010010010: data <= 15'h7ff5; 
        10'b0010010011: data <= 15'h7fea; 
        10'b0010010100: data <= 15'h0010; 
        10'b0010010101: data <= 15'h7feb; 
        10'b0010010110: data <= 15'h0007; 
        10'b0010010111: data <= 15'h7fb9; 
        10'b0010011000: data <= 15'h7fda; 
        10'b0010011001: data <= 15'h7fe6; 
        10'b0010011010: data <= 15'h7ff6; 
        10'b0010011011: data <= 15'h7fde; 
        10'b0010011100: data <= 15'h7fde; 
        10'b0010011101: data <= 15'h0006; 
        10'b0010011110: data <= 15'h002e; 
        10'b0010011111: data <= 15'h0056; 
        10'b0010100000: data <= 15'h004b; 
        10'b0010100001: data <= 15'h0043; 
        10'b0010100010: data <= 15'h0035; 
        10'b0010100011: data <= 15'h0024; 
        10'b0010100100: data <= 15'h7ffc; 
        10'b0010100101: data <= 15'h0002; 
        10'b0010100110: data <= 15'h7fee; 
        10'b0010100111: data <= 15'h0011; 
        10'b0010101000: data <= 15'h7ffe; 
        10'b0010101001: data <= 15'h000f; 
        10'b0010101010: data <= 15'h000e; 
        10'b0010101011: data <= 15'h7fed; 
        10'b0010101100: data <= 15'h0007; 
        10'b0010101101: data <= 15'h7ffd; 
        10'b0010101110: data <= 15'h0006; 
        10'b0010101111: data <= 15'h0000; 
        10'b0010110000: data <= 15'h7fe5; 
        10'b0010110001: data <= 15'h7fe0; 
        10'b0010110010: data <= 15'h7fae; 
        10'b0010110011: data <= 15'h7f95; 
        10'b0010110100: data <= 15'h7fc2; 
        10'b0010110101: data <= 15'h7f86; 
        10'b0010110110: data <= 15'h7fca; 
        10'b0010110111: data <= 15'h7fd8; 
        10'b0010111000: data <= 15'h7fc7; 
        10'b0010111001: data <= 15'h7fce; 
        10'b0010111010: data <= 15'h7ff2; 
        10'b0010111011: data <= 15'h7fde; 
        10'b0010111100: data <= 15'h7fca; 
        10'b0010111101: data <= 15'h7fcc; 
        10'b0010111110: data <= 15'h7fb0; 
        10'b0010111111: data <= 15'h7fcc; 
        10'b0011000000: data <= 15'h7fd4; 
        10'b0011000001: data <= 15'h7fd2; 
        10'b0011000010: data <= 15'h7ff9; 
        10'b0011000011: data <= 15'h000f; 
        10'b0011000100: data <= 15'h0006; 
        10'b0011000101: data <= 15'h0009; 
        10'b0011000110: data <= 15'h0001; 
        10'b0011000111: data <= 15'h7ffd; 
        10'b0011001000: data <= 15'h0001; 
        10'b0011001001: data <= 15'h7ff0; 
        10'b0011001010: data <= 15'h7fe0; 
        10'b0011001011: data <= 15'h7ffb; 
        10'b0011001100: data <= 15'h7fd2; 
        10'b0011001101: data <= 15'h7fc7; 
        10'b0011001110: data <= 15'h7fad; 
        10'b0011001111: data <= 15'h7fbf; 
        10'b0011010000: data <= 15'h7f8b; 
        10'b0011010001: data <= 15'h7f7d; 
        10'b0011010010: data <= 15'h7fbb; 
        10'b0011010011: data <= 15'h7fbf; 
        10'b0011010100: data <= 15'h7f9a; 
        10'b0011010101: data <= 15'h7f9f; 
        10'b0011010110: data <= 15'h7f88; 
        10'b0011010111: data <= 15'h7f5d; 
        10'b0011011000: data <= 15'h7f5a; 
        10'b0011011001: data <= 15'h7f75; 
        10'b0011011010: data <= 15'h7f6f; 
        10'b0011011011: data <= 15'h7f8d; 
        10'b0011011100: data <= 15'h7fd4; 
        10'b0011011101: data <= 15'h7fd8; 
        10'b0011011110: data <= 15'h7ff0; 
        10'b0011011111: data <= 15'h7ff4; 
        10'b0011100000: data <= 15'h7ffa; 
        10'b0011100001: data <= 15'h7ffb; 
        10'b0011100010: data <= 15'h0012; 
        10'b0011100011: data <= 15'h7fea; 
        10'b0011100100: data <= 15'h7fed; 
        10'b0011100101: data <= 15'h7fe7; 
        10'b0011100110: data <= 15'h7fc2; 
        10'b0011100111: data <= 15'h7ff2; 
        10'b0011101000: data <= 15'h7fe9; 
        10'b0011101001: data <= 15'h7fbf; 
        10'b0011101010: data <= 15'h7fb4; 
        10'b0011101011: data <= 15'h7fa9; 
        10'b0011101100: data <= 15'h7f97; 
        10'b0011101101: data <= 15'h7f86; 
        10'b0011101110: data <= 15'h7f89; 
        10'b0011101111: data <= 15'h7f81; 
        10'b0011110000: data <= 15'h7f6a; 
        10'b0011110001: data <= 15'h7f53; 
        10'b0011110010: data <= 15'h7f0b; 
        10'b0011110011: data <= 15'h7f1c; 
        10'b0011110100: data <= 15'h7f34; 
        10'b0011110101: data <= 15'h7f36; 
        10'b0011110110: data <= 15'h7f73; 
        10'b0011110111: data <= 15'h7f84; 
        10'b0011111000: data <= 15'h7fb2; 
        10'b0011111001: data <= 15'h7fcf; 
        10'b0011111010: data <= 15'h7fdd; 
        10'b0011111011: data <= 15'h0005; 
        10'b0011111100: data <= 15'h7ffd; 
        10'b0011111101: data <= 15'h7ff2; 
        10'b0011111110: data <= 15'h7ff8; 
        10'b0011111111: data <= 15'h7ff0; 
        10'b0100000000: data <= 15'h0000; 
        10'b0100000001: data <= 15'h7ff2; 
        10'b0100000010: data <= 15'h7fea; 
        10'b0100000011: data <= 15'h7ff3; 
        10'b0100000100: data <= 15'h000f; 
        10'b0100000101: data <= 15'h7fd9; 
        10'b0100000110: data <= 15'h7fb6; 
        10'b0100000111: data <= 15'h7fc7; 
        10'b0100001000: data <= 15'h7fdb; 
        10'b0100001001: data <= 15'h7fbb; 
        10'b0100001010: data <= 15'h7fc0; 
        10'b0100001011: data <= 15'h7f75; 
        10'b0100001100: data <= 15'h7f5e; 
        10'b0100001101: data <= 15'h7f15; 
        10'b0100001110: data <= 15'h7f06; 
        10'b0100001111: data <= 15'h7f34; 
        10'b0100010000: data <= 15'h7f58; 
        10'b0100010001: data <= 15'h7f7b; 
        10'b0100010010: data <= 15'h7f66; 
        10'b0100010011: data <= 15'h7f9d; 
        10'b0100010100: data <= 15'h7fb4; 
        10'b0100010101: data <= 15'h7fc8; 
        10'b0100010110: data <= 15'h7fe9; 
        10'b0100010111: data <= 15'h000c; 
        10'b0100011000: data <= 15'h7ff4; 
        10'b0100011001: data <= 15'h000f; 
        10'b0100011010: data <= 15'h000a; 
        10'b0100011011: data <= 15'h7fee; 
        10'b0100011100: data <= 15'h7fe6; 
        10'b0100011101: data <= 15'h0007; 
        10'b0100011110: data <= 15'h0016; 
        10'b0100011111: data <= 15'h0015; 
        10'b0100100000: data <= 15'h004c; 
        10'b0100100001: data <= 15'h7ffe; 
        10'b0100100010: data <= 15'h000f; 
        10'b0100100011: data <= 15'h0006; 
        10'b0100100100: data <= 15'h7fd2; 
        10'b0100100101: data <= 15'h7fe1; 
        10'b0100100110: data <= 15'h7fbb; 
        10'b0100100111: data <= 15'h7f70; 
        10'b0100101000: data <= 15'h7f6e; 
        10'b0100101001: data <= 15'h7f54; 
        10'b0100101010: data <= 15'h7f4d; 
        10'b0100101011: data <= 15'h7f71; 
        10'b0100101100: data <= 15'h7f9f; 
        10'b0100101101: data <= 15'h7fbb; 
        10'b0100101110: data <= 15'h7fa5; 
        10'b0100101111: data <= 15'h7ff6; 
        10'b0100110000: data <= 15'h7fc5; 
        10'b0100110001: data <= 15'h7fd7; 
        10'b0100110010: data <= 15'h7ff4; 
        10'b0100110011: data <= 15'h7ffa; 
        10'b0100110100: data <= 15'h7ff6; 
        10'b0100110101: data <= 15'h0006; 
        10'b0100110110: data <= 15'h7ff6; 
        10'b0100110111: data <= 15'h7fff; 
        10'b0100111000: data <= 15'h7ff6; 
        10'b0100111001: data <= 15'h0003; 
        10'b0100111010: data <= 15'h7ffa; 
        10'b0100111011: data <= 15'h0040; 
        10'b0100111100: data <= 15'h002d; 
        10'b0100111101: data <= 15'h0016; 
        10'b0100111110: data <= 15'h001c; 
        10'b0100111111: data <= 15'h0013; 
        10'b0101000000: data <= 15'h0013; 
        10'b0101000001: data <= 15'h0003; 
        10'b0101000010: data <= 15'h7fdf; 
        10'b0101000011: data <= 15'h7f8e; 
        10'b0101000100: data <= 15'h7f95; 
        10'b0101000101: data <= 15'h7fa5; 
        10'b0101000110: data <= 15'h7fa5; 
        10'b0101000111: data <= 15'h7fb9; 
        10'b0101001000: data <= 15'h7fdf; 
        10'b0101001001: data <= 15'h000d; 
        10'b0101001010: data <= 15'h002c; 
        10'b0101001011: data <= 15'h0044; 
        10'b0101001100: data <= 15'h0000; 
        10'b0101001101: data <= 15'h7fdc; 
        10'b0101001110: data <= 15'h7ff1; 
        10'b0101001111: data <= 15'h7ffa; 
        10'b0101010000: data <= 15'h7ff6; 
        10'b0101010001: data <= 15'h7ffb; 
        10'b0101010010: data <= 15'h7ff0; 
        10'b0101010011: data <= 15'h7ff9; 
        10'b0101010100: data <= 15'h0009; 
        10'b0101010101: data <= 15'h001e; 
        10'b0101010110: data <= 15'h002d; 
        10'b0101010111: data <= 15'h003c; 
        10'b0101011000: data <= 15'h001c; 
        10'b0101011001: data <= 15'h0027; 
        10'b0101011010: data <= 15'h001b; 
        10'b0101011011: data <= 15'h0048; 
        10'b0101011100: data <= 15'h0045; 
        10'b0101011101: data <= 15'h0031; 
        10'b0101011110: data <= 15'h7fd6; 
        10'b0101011111: data <= 15'h7fb3; 
        10'b0101100000: data <= 15'h7ffd; 
        10'b0101100001: data <= 15'h7ff9; 
        10'b0101100010: data <= 15'h7fb5; 
        10'b0101100011: data <= 15'h7fb8; 
        10'b0101100100: data <= 15'h7ff7; 
        10'b0101100101: data <= 15'h0029; 
        10'b0101100110: data <= 15'h0062; 
        10'b0101100111: data <= 15'h00ae; 
        10'b0101101000: data <= 15'h005e; 
        10'b0101101001: data <= 15'h7fe5; 
        10'b0101101010: data <= 15'h7fe1; 
        10'b0101101011: data <= 15'h7ff7; 
        10'b0101101100: data <= 15'h7ff7; 
        10'b0101101101: data <= 15'h0010; 
        10'b0101101110: data <= 15'h000c; 
        10'b0101101111: data <= 15'h7fee; 
        10'b0101110000: data <= 15'h7fe8; 
        10'b0101110001: data <= 15'h000a; 
        10'b0101110010: data <= 15'h004b; 
        10'b0101110011: data <= 15'h0029; 
        10'b0101110100: data <= 15'h0023; 
        10'b0101110101: data <= 15'h0011; 
        10'b0101110110: data <= 15'h0049; 
        10'b0101110111: data <= 15'h003d; 
        10'b0101111000: data <= 15'h0038; 
        10'b0101111001: data <= 15'h000a; 
        10'b0101111010: data <= 15'h7ff6; 
        10'b0101111011: data <= 15'h7ffe; 
        10'b0101111100: data <= 15'h0006; 
        10'b0101111101: data <= 15'h7ff0; 
        10'b0101111110: data <= 15'h7fbf; 
        10'b0101111111: data <= 15'h7ff7; 
        10'b0110000000: data <= 15'h7fe1; 
        10'b0110000001: data <= 15'h0034; 
        10'b0110000010: data <= 15'h0088; 
        10'b0110000011: data <= 15'h00d7; 
        10'b0110000100: data <= 15'h0074; 
        10'b0110000101: data <= 15'h7ff7; 
        10'b0110000110: data <= 15'h0000; 
        10'b0110000111: data <= 15'h000b; 
        10'b0110001000: data <= 15'h7ff8; 
        10'b0110001001: data <= 15'h0002; 
        10'b0110001010: data <= 15'h000c; 
        10'b0110001011: data <= 15'h0001; 
        10'b0110001100: data <= 15'h7fe7; 
        10'b0110001101: data <= 15'h001b; 
        10'b0110001110: data <= 15'h0045; 
        10'b0110001111: data <= 15'h003c; 
        10'b0110010000: data <= 15'h0052; 
        10'b0110010001: data <= 15'h004d; 
        10'b0110010010: data <= 15'h0053; 
        10'b0110010011: data <= 15'h005a; 
        10'b0110010100: data <= 15'h001e; 
        10'b0110010101: data <= 15'h7fd4; 
        10'b0110010110: data <= 15'h0003; 
        10'b0110010111: data <= 15'h0025; 
        10'b0110011000: data <= 15'h0011; 
        10'b0110011001: data <= 15'h7fe3; 
        10'b0110011010: data <= 15'h7fe4; 
        10'b0110011011: data <= 15'h7ffc; 
        10'b0110011100: data <= 15'h003b; 
        10'b0110011101: data <= 15'h003a; 
        10'b0110011110: data <= 15'h009a; 
        10'b0110011111: data <= 15'h00b3; 
        10'b0110100000: data <= 15'h0075; 
        10'b0110100001: data <= 15'h7ffe; 
        10'b0110100010: data <= 15'h7fde; 
        10'b0110100011: data <= 15'h7fef; 
        10'b0110100100: data <= 15'h000d; 
        10'b0110100101: data <= 15'h7ffa; 
        10'b0110100110: data <= 15'h0002; 
        10'b0110100111: data <= 15'h7ff2; 
        10'b0110101000: data <= 15'h7fcf; 
        10'b0110101001: data <= 15'h7ffa; 
        10'b0110101010: data <= 15'h0048; 
        10'b0110101011: data <= 15'h0060; 
        10'b0110101100: data <= 15'h003e; 
        10'b0110101101: data <= 15'h0061; 
        10'b0110101110: data <= 15'h007a; 
        10'b0110101111: data <= 15'h0095; 
        10'b0110110000: data <= 15'h0027; 
        10'b0110110001: data <= 15'h7ff5; 
        10'b0110110010: data <= 15'h003a; 
        10'b0110110011: data <= 15'h0035; 
        10'b0110110100: data <= 15'h0008; 
        10'b0110110101: data <= 15'h7fe5; 
        10'b0110110110: data <= 15'h0005; 
        10'b0110110111: data <= 15'h001e; 
        10'b0110111000: data <= 15'h0045; 
        10'b0110111001: data <= 15'h005f; 
        10'b0110111010: data <= 15'h0057; 
        10'b0110111011: data <= 15'h006c; 
        10'b0110111100: data <= 15'h0039; 
        10'b0110111101: data <= 15'h7fe3; 
        10'b0110111110: data <= 15'h7fee; 
        10'b0110111111: data <= 15'h7fed; 
        10'b0111000000: data <= 15'h0003; 
        10'b0111000001: data <= 15'h7ff2; 
        10'b0111000010: data <= 15'h7ff2; 
        10'b0111000011: data <= 15'h7ff0; 
        10'b0111000100: data <= 15'h7fc0; 
        10'b0111000101: data <= 15'h7fdd; 
        10'b0111000110: data <= 15'h006b; 
        10'b0111000111: data <= 15'h006d; 
        10'b0111001000: data <= 15'h0048; 
        10'b0111001001: data <= 15'h006f; 
        10'b0111001010: data <= 15'h00bd; 
        10'b0111001011: data <= 15'h00bc; 
        10'b0111001100: data <= 15'h0039; 
        10'b0111001101: data <= 15'h0022; 
        10'b0111001110: data <= 15'h0052; 
        10'b0111001111: data <= 15'h002b; 
        10'b0111010000: data <= 15'h7fea; 
        10'b0111010001: data <= 15'h7fd3; 
        10'b0111010010: data <= 15'h000f; 
        10'b0111010011: data <= 15'h0030; 
        10'b0111010100: data <= 15'h0016; 
        10'b0111010101: data <= 15'h0001; 
        10'b0111010110: data <= 15'h002c; 
        10'b0111010111: data <= 15'h001b; 
        10'b0111011000: data <= 15'h7ff3; 
        10'b0111011001: data <= 15'h7fdd; 
        10'b0111011010: data <= 15'h7feb; 
        10'b0111011011: data <= 15'h7ffd; 
        10'b0111011100: data <= 15'h0003; 
        10'b0111011101: data <= 15'h000b; 
        10'b0111011110: data <= 15'h000f; 
        10'b0111011111: data <= 15'h7ffd; 
        10'b0111100000: data <= 15'h7fa5; 
        10'b0111100001: data <= 15'h7fd0; 
        10'b0111100010: data <= 15'h002d; 
        10'b0111100011: data <= 15'h0055; 
        10'b0111100100: data <= 15'h0061; 
        10'b0111100101: data <= 15'h007a; 
        10'b0111100110: data <= 15'h00d2; 
        10'b0111100111: data <= 15'h00d6; 
        10'b0111101000: data <= 15'h006e; 
        10'b0111101001: data <= 15'h003e; 
        10'b0111101010: data <= 15'h003f; 
        10'b0111101011: data <= 15'h0028; 
        10'b0111101100: data <= 15'h0000; 
        10'b0111101101: data <= 15'h000b; 
        10'b0111101110: data <= 15'h0058; 
        10'b0111101111: data <= 15'h001e; 
        10'b0111110000: data <= 15'h000d; 
        10'b0111110001: data <= 15'h7fea; 
        10'b0111110010: data <= 15'h0014; 
        10'b0111110011: data <= 15'h7ffc; 
        10'b0111110100: data <= 15'h7fe7; 
        10'b0111110101: data <= 15'h7fd0; 
        10'b0111110110: data <= 15'h7ff9; 
        10'b0111110111: data <= 15'h0008; 
        10'b0111111000: data <= 15'h7ff9; 
        10'b0111111001: data <= 15'h7ff6; 
        10'b0111111010: data <= 15'h0000; 
        10'b0111111011: data <= 15'h7fe5; 
        10'b0111111100: data <= 15'h7faa; 
        10'b0111111101: data <= 15'h7fac; 
        10'b0111111110: data <= 15'h7fd7; 
        10'b0111111111: data <= 15'h003a; 
        10'b1000000000: data <= 15'h005e; 
        10'b1000000001: data <= 15'h0055; 
        10'b1000000010: data <= 15'h0093; 
        10'b1000000011: data <= 15'h00b6; 
        10'b1000000100: data <= 15'h00d6; 
        10'b1000000101: data <= 15'h0063; 
        10'b1000000110: data <= 15'h001b; 
        10'b1000000111: data <= 15'h0037; 
        10'b1000001000: data <= 15'h0060; 
        10'b1000001001: data <= 15'h003e; 
        10'b1000001010: data <= 15'h004d; 
        10'b1000001011: data <= 15'h0029; 
        10'b1000001100: data <= 15'h0005; 
        10'b1000001101: data <= 15'h000e; 
        10'b1000001110: data <= 15'h000f; 
        10'b1000001111: data <= 15'h7ff8; 
        10'b1000010000: data <= 15'h7fe1; 
        10'b1000010001: data <= 15'h7fe9; 
        10'b1000010010: data <= 15'h7fef; 
        10'b1000010011: data <= 15'h7fed; 
        10'b1000010100: data <= 15'h0005; 
        10'b1000010101: data <= 15'h7ff3; 
        10'b1000010110: data <= 15'h0008; 
        10'b1000010111: data <= 15'h7fde; 
        10'b1000011000: data <= 15'h7fc8; 
        10'b1000011001: data <= 15'h7fa7; 
        10'b1000011010: data <= 15'h7fbb; 
        10'b1000011011: data <= 15'h0005; 
        10'b1000011100: data <= 15'h003d; 
        10'b1000011101: data <= 15'h005f; 
        10'b1000011110: data <= 15'h007f; 
        10'b1000011111: data <= 15'h00cb; 
        10'b1000100000: data <= 15'h00e4; 
        10'b1000100001: data <= 15'h0075; 
        10'b1000100010: data <= 15'h0069; 
        10'b1000100011: data <= 15'h006e; 
        10'b1000100100: data <= 15'h004e; 
        10'b1000100101: data <= 15'h0040; 
        10'b1000100110: data <= 15'h0064; 
        10'b1000100111: data <= 15'h0044; 
        10'b1000101000: data <= 15'h002c; 
        10'b1000101001: data <= 15'h0009; 
        10'b1000101010: data <= 15'h7ff0; 
        10'b1000101011: data <= 15'h7fec; 
        10'b1000101100: data <= 15'h7feb; 
        10'b1000101101: data <= 15'h7ffd; 
        10'b1000101110: data <= 15'h7ff6; 
        10'b1000101111: data <= 15'h000f; 
        10'b1000110000: data <= 15'h7ff7; 
        10'b1000110001: data <= 15'h7ff3; 
        10'b1000110010: data <= 15'h7ffb; 
        10'b1000110011: data <= 15'h7ff1; 
        10'b1000110100: data <= 15'h7fb9; 
        10'b1000110101: data <= 15'h7fab; 
        10'b1000110110: data <= 15'h7fb6; 
        10'b1000110111: data <= 15'h7fe2; 
        10'b1000111000: data <= 15'h0014; 
        10'b1000111001: data <= 15'h0040; 
        10'b1000111010: data <= 15'h0069; 
        10'b1000111011: data <= 15'h0046; 
        10'b1000111100: data <= 15'h008a; 
        10'b1000111101: data <= 15'h00a6; 
        10'b1000111110: data <= 15'h00c4; 
        10'b1000111111: data <= 15'h00a7; 
        10'b1001000000: data <= 15'h005b; 
        10'b1001000001: data <= 15'h003a; 
        10'b1001000010: data <= 15'h0071; 
        10'b1001000011: data <= 15'h004f; 
        10'b1001000100: data <= 15'h0036; 
        10'b1001000101: data <= 15'h7ff5; 
        10'b1001000110: data <= 15'h7fd6; 
        10'b1001000111: data <= 15'h0003; 
        10'b1001001000: data <= 15'h7ff6; 
        10'b1001001001: data <= 15'h7ffb; 
        10'b1001001010: data <= 15'h7ff3; 
        10'b1001001011: data <= 15'h0003; 
        10'b1001001100: data <= 15'h7ffe; 
        10'b1001001101: data <= 15'h0002; 
        10'b1001001110: data <= 15'h0005; 
        10'b1001001111: data <= 15'h7ffb; 
        10'b1001010000: data <= 15'h7fe5; 
        10'b1001010001: data <= 15'h7fc5; 
        10'b1001010010: data <= 15'h7f9d; 
        10'b1001010011: data <= 15'h7fd3; 
        10'b1001010100: data <= 15'h7fe5; 
        10'b1001010101: data <= 15'h0030; 
        10'b1001010110: data <= 15'h0057; 
        10'b1001010111: data <= 15'h007c; 
        10'b1001011000: data <= 15'h00a0; 
        10'b1001011001: data <= 15'h00a2; 
        10'b1001011010: data <= 15'h0088; 
        10'b1001011011: data <= 15'h0075; 
        10'b1001011100: data <= 15'h0049; 
        10'b1001011101: data <= 15'h0064; 
        10'b1001011110: data <= 15'h005d; 
        10'b1001011111: data <= 15'h003c; 
        10'b1001100000: data <= 15'h0008; 
        10'b1001100001: data <= 15'h7fe0; 
        10'b1001100010: data <= 15'h7fd4; 
        10'b1001100011: data <= 15'h7fe6; 
        10'b1001100100: data <= 15'h0001; 
        10'b1001100101: data <= 15'h7fef; 
        10'b1001100110: data <= 15'h7ffc; 
        10'b1001100111: data <= 15'h7ff7; 
        10'b1001101000: data <= 15'h7ff7; 
        10'b1001101001: data <= 15'h7ffe; 
        10'b1001101010: data <= 15'h0010; 
        10'b1001101011: data <= 15'h0004; 
        10'b1001101100: data <= 15'h7ff7; 
        10'b1001101101: data <= 15'h7fcd; 
        10'b1001101110: data <= 15'h7fc3; 
        10'b1001101111: data <= 15'h7faf; 
        10'b1001110000: data <= 15'h7fca; 
        10'b1001110001: data <= 15'h7fe7; 
        10'b1001110010: data <= 15'h7fec; 
        10'b1001110011: data <= 15'h000a; 
        10'b1001110100: data <= 15'h002f; 
        10'b1001110101: data <= 15'h0014; 
        10'b1001110110: data <= 15'h0011; 
        10'b1001110111: data <= 15'h0032; 
        10'b1001111000: data <= 15'h0026; 
        10'b1001111001: data <= 15'h0000; 
        10'b1001111010: data <= 15'h7ff3; 
        10'b1001111011: data <= 15'h7fc8; 
        10'b1001111100: data <= 15'h7fca; 
        10'b1001111101: data <= 15'h7fd3; 
        10'b1001111110: data <= 15'h7fd6; 
        10'b1001111111: data <= 15'h7ffc; 
        10'b1010000000: data <= 15'h7ff9; 
        10'b1010000001: data <= 15'h7ff0; 
        10'b1010000010: data <= 15'h0011; 
        10'b1010000011: data <= 15'h0007; 
        10'b1010000100: data <= 15'h000e; 
        10'b1010000101: data <= 15'h7ffb; 
        10'b1010000110: data <= 15'h7ff8; 
        10'b1010000111: data <= 15'h0002; 
        10'b1010001000: data <= 15'h0005; 
        10'b1010001001: data <= 15'h7feb; 
        10'b1010001010: data <= 15'h7fdf; 
        10'b1010001011: data <= 15'h7fb8; 
        10'b1010001100: data <= 15'h7fa5; 
        10'b1010001101: data <= 15'h7f7c; 
        10'b1010001110: data <= 15'h7f7d; 
        10'b1010001111: data <= 15'h7f67; 
        10'b1010010000: data <= 15'h7fa2; 
        10'b1010010001: data <= 15'h7fb6; 
        10'b1010010010: data <= 15'h7fc6; 
        10'b1010010011: data <= 15'h7faa; 
        10'b1010010100: data <= 15'h7f8f; 
        10'b1010010101: data <= 15'h7f80; 
        10'b1010010110: data <= 15'h7f9b; 
        10'b1010010111: data <= 15'h7fd2; 
        10'b1010011000: data <= 15'h7fd1; 
        10'b1010011001: data <= 15'h7fd7; 
        10'b1010011010: data <= 15'h7ff1; 
        10'b1010011011: data <= 15'h0002; 
        10'b1010011100: data <= 15'h7fef; 
        10'b1010011101: data <= 15'h7ff2; 
        10'b1010011110: data <= 15'h7ffa; 
        10'b1010011111: data <= 15'h7ffe; 
        10'b1010100000: data <= 15'h000a; 
        10'b1010100001: data <= 15'h0008; 
        10'b1010100010: data <= 15'h0005; 
        10'b1010100011: data <= 15'h7ff0; 
        10'b1010100100: data <= 15'h7ff3; 
        10'b1010100101: data <= 15'h7ffa; 
        10'b1010100110: data <= 15'h7ff0; 
        10'b1010100111: data <= 15'h7fe7; 
        10'b1010101000: data <= 15'h7fec; 
        10'b1010101001: data <= 15'h7fe0; 
        10'b1010101010: data <= 15'h7fd0; 
        10'b1010101011: data <= 15'h7fc4; 
        10'b1010101100: data <= 15'h7fba; 
        10'b1010101101: data <= 15'h7fbb; 
        10'b1010101110: data <= 15'h7fb0; 
        10'b1010101111: data <= 15'h7fb0; 
        10'b1010110000: data <= 15'h7fac; 
        10'b1010110001: data <= 15'h7fc0; 
        10'b1010110010: data <= 15'h7fea; 
        10'b1010110011: data <= 15'h7feb; 
        10'b1010110100: data <= 15'h7ff9; 
        10'b1010110101: data <= 15'h7ff5; 
        10'b1010110110: data <= 15'h0008; 
        10'b1010110111: data <= 15'h7ffc; 
        10'b1010111000: data <= 15'h7fef; 
        10'b1010111001: data <= 15'h7ffb; 
        10'b1010111010: data <= 15'h7ff4; 
        10'b1010111011: data <= 15'h7ff4; 
        10'b1010111100: data <= 15'h0010; 
        10'b1010111101: data <= 15'h7ff1; 
        10'b1010111110: data <= 15'h0004; 
        10'b1010111111: data <= 15'h7ff9; 
        10'b1011000000: data <= 15'h7ff5; 
        10'b1011000001: data <= 15'h7ffe; 
        10'b1011000010: data <= 15'h000a; 
        10'b1011000011: data <= 15'h7fff; 
        10'b1011000100: data <= 15'h7fee; 
        10'b1011000101: data <= 15'h0006; 
        10'b1011000110: data <= 15'h7fef; 
        10'b1011000111: data <= 15'h7ffd; 
        10'b1011001000: data <= 15'h0001; 
        10'b1011001001: data <= 15'h7fee; 
        10'b1011001010: data <= 15'h7ff6; 
        10'b1011001011: data <= 15'h7ffa; 
        10'b1011001100: data <= 15'h7ffe; 
        10'b1011001101: data <= 15'h7ff0; 
        10'b1011001110: data <= 15'h7ff7; 
        10'b1011001111: data <= 15'h7fee; 
        10'b1011010000: data <= 15'h7ff2; 
        10'b1011010001: data <= 15'h0002; 
        10'b1011010010: data <= 15'h7ff9; 
        10'b1011010011: data <= 15'h000d; 
        10'b1011010100: data <= 15'h0012; 
        10'b1011010101: data <= 15'h0010; 
        10'b1011010110: data <= 15'h0001; 
        10'b1011010111: data <= 15'h000c; 
        10'b1011011000: data <= 15'h0011; 
        10'b1011011001: data <= 15'h7fff; 
        10'b1011011010: data <= 15'h0003; 
        10'b1011011011: data <= 15'h7ffd; 
        10'b1011011100: data <= 15'h7ff7; 
        10'b1011011101: data <= 15'h000e; 
        10'b1011011110: data <= 15'h000b; 
        10'b1011011111: data <= 15'h7ff7; 
        10'b1011100000: data <= 15'h7ffa; 
        10'b1011100001: data <= 15'h0008; 
        10'b1011100010: data <= 15'h7ff9; 
        10'b1011100011: data <= 15'h0004; 
        10'b1011100100: data <= 15'h7ff9; 
        10'b1011100101: data <= 15'h000a; 
        10'b1011100110: data <= 15'h000b; 
        10'b1011100111: data <= 15'h7ff2; 
        10'b1011101000: data <= 15'h7ff5; 
        10'b1011101001: data <= 15'h000e; 
        10'b1011101010: data <= 15'h000b; 
        10'b1011101011: data <= 15'h7ffa; 
        10'b1011101100: data <= 15'h000a; 
        10'b1011101101: data <= 15'h7ffc; 
        10'b1011101110: data <= 15'h7ffc; 
        10'b1011101111: data <= 15'h0006; 
        10'b1011110000: data <= 15'h0007; 
        10'b1011110001: data <= 15'h7ffc; 
        10'b1011110010: data <= 15'h7ff8; 
        10'b1011110011: data <= 15'h7ffb; 
        10'b1011110100: data <= 15'h0010; 
        10'b1011110101: data <= 15'h7fff; 
        10'b1011110110: data <= 15'h0009; 
        10'b1011110111: data <= 15'h7ff7; 
        10'b1011111000: data <= 15'h0006; 
        10'b1011111001: data <= 15'h0000; 
        10'b1011111010: data <= 15'h000f; 
        10'b1011111011: data <= 15'h0002; 
        10'b1011111100: data <= 15'h7ffe; 
        10'b1011111101: data <= 15'h7fee; 
        10'b1011111110: data <= 15'h7ff4; 
        10'b1011111111: data <= 15'h0006; 
        10'b1100000000: data <= 15'h7ff0; 
        10'b1100000001: data <= 15'h7ff2; 
        10'b1100000010: data <= 15'h7ff6; 
        10'b1100000011: data <= 15'h7fef; 
        10'b1100000100: data <= 15'h7ff5; 
        10'b1100000101: data <= 15'h7ffa; 
        10'b1100000110: data <= 15'h7ff1; 
        10'b1100000111: data <= 15'h7ff5; 
        10'b1100001000: data <= 15'h7ff6; 
        10'b1100001001: data <= 15'h7ff8; 
        10'b1100001010: data <= 15'h000f; 
        10'b1100001011: data <= 15'h7ff1; 
        10'b1100001100: data <= 15'h7ff6; 
        10'b1100001101: data <= 15'h7ff2; 
        10'b1100001110: data <= 15'h7ff6; 
        10'b1100001111: data <= 15'h0003; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 10) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 16'hfff5; 
        10'b0000000001: data <= 16'h0017; 
        10'b0000000010: data <= 16'hffe6; 
        10'b0000000011: data <= 16'hfffe; 
        10'b0000000100: data <= 16'hffff; 
        10'b0000000101: data <= 16'hfffc; 
        10'b0000000110: data <= 16'h000c; 
        10'b0000000111: data <= 16'h0025; 
        10'b0000001000: data <= 16'hffe8; 
        10'b0000001001: data <= 16'hfff0; 
        10'b0000001010: data <= 16'hfff1; 
        10'b0000001011: data <= 16'hffe9; 
        10'b0000001100: data <= 16'h000c; 
        10'b0000001101: data <= 16'h0022; 
        10'b0000001110: data <= 16'h0013; 
        10'b0000001111: data <= 16'hffe1; 
        10'b0000010000: data <= 16'hfffc; 
        10'b0000010001: data <= 16'h0025; 
        10'b0000010010: data <= 16'h0006; 
        10'b0000010011: data <= 16'hfffd; 
        10'b0000010100: data <= 16'hffe4; 
        10'b0000010101: data <= 16'hffed; 
        10'b0000010110: data <= 16'h0009; 
        10'b0000010111: data <= 16'h0020; 
        10'b0000011000: data <= 16'h0011; 
        10'b0000011001: data <= 16'h0015; 
        10'b0000011010: data <= 16'hffe3; 
        10'b0000011011: data <= 16'hffe4; 
        10'b0000011100: data <= 16'h0018; 
        10'b0000011101: data <= 16'h0013; 
        10'b0000011110: data <= 16'h0018; 
        10'b0000011111: data <= 16'hfffa; 
        10'b0000100000: data <= 16'hffe0; 
        10'b0000100001: data <= 16'hffed; 
        10'b0000100010: data <= 16'h0010; 
        10'b0000100011: data <= 16'h0036; 
        10'b0000100100: data <= 16'h0024; 
        10'b0000100101: data <= 16'h000b; 
        10'b0000100110: data <= 16'h002c; 
        10'b0000100111: data <= 16'h002f; 
        10'b0000101000: data <= 16'h0032; 
        10'b0000101001: data <= 16'h002f; 
        10'b0000101010: data <= 16'h001e; 
        10'b0000101011: data <= 16'h0020; 
        10'b0000101100: data <= 16'hffde; 
        10'b0000101101: data <= 16'h001e; 
        10'b0000101110: data <= 16'h0029; 
        10'b0000101111: data <= 16'h0017; 
        10'b0000110000: data <= 16'hfff9; 
        10'b0000110001: data <= 16'hffeb; 
        10'b0000110010: data <= 16'h002c; 
        10'b0000110011: data <= 16'h0021; 
        10'b0000110100: data <= 16'hfff2; 
        10'b0000110101: data <= 16'h0025; 
        10'b0000110110: data <= 16'hfffa; 
        10'b0000110111: data <= 16'h001b; 
        10'b0000111000: data <= 16'hffeb; 
        10'b0000111001: data <= 16'hffe6; 
        10'b0000111010: data <= 16'hffe0; 
        10'b0000111011: data <= 16'hfffd; 
        10'b0000111100: data <= 16'h0012; 
        10'b0000111101: data <= 16'h000b; 
        10'b0000111110: data <= 16'h0013; 
        10'b0000111111: data <= 16'h0034; 
        10'b0001000000: data <= 16'h0025; 
        10'b0001000001: data <= 16'h0050; 
        10'b0001000010: data <= 16'h0064; 
        10'b0001000011: data <= 16'h0071; 
        10'b0001000100: data <= 16'h0071; 
        10'b0001000101: data <= 16'h0077; 
        10'b0001000110: data <= 16'h003c; 
        10'b0001000111: data <= 16'h002b; 
        10'b0001001000: data <= 16'h0063; 
        10'b0001001001: data <= 16'h002c; 
        10'b0001001010: data <= 16'h002b; 
        10'b0001001011: data <= 16'h002f; 
        10'b0001001100: data <= 16'h002e; 
        10'b0001001101: data <= 16'h0017; 
        10'b0001001110: data <= 16'h001e; 
        10'b0001001111: data <= 16'h0006; 
        10'b0001010000: data <= 16'h0011; 
        10'b0001010001: data <= 16'hfff6; 
        10'b0001010010: data <= 16'hffde; 
        10'b0001010011: data <= 16'h000a; 
        10'b0001010100: data <= 16'hffe3; 
        10'b0001010101: data <= 16'h0003; 
        10'b0001010110: data <= 16'h001b; 
        10'b0001010111: data <= 16'h0010; 
        10'b0001011000: data <= 16'h0023; 
        10'b0001011001: data <= 16'hffe1; 
        10'b0001011010: data <= 16'h0026; 
        10'b0001011011: data <= 16'h002a; 
        10'b0001011100: data <= 16'h0032; 
        10'b0001011101: data <= 16'h0065; 
        10'b0001011110: data <= 16'h005a; 
        10'b0001011111: data <= 16'h0070; 
        10'b0001100000: data <= 16'h006e; 
        10'b0001100001: data <= 16'h006a; 
        10'b0001100010: data <= 16'h009b; 
        10'b0001100011: data <= 16'h0093; 
        10'b0001100100: data <= 16'h005b; 
        10'b0001100101: data <= 16'h0073; 
        10'b0001100110: data <= 16'h00b9; 
        10'b0001100111: data <= 16'h00b8; 
        10'b0001101000: data <= 16'h00c5; 
        10'b0001101001: data <= 16'h00ae; 
        10'b0001101010: data <= 16'h00b0; 
        10'b0001101011: data <= 16'h0066; 
        10'b0001101100: data <= 16'h005b; 
        10'b0001101101: data <= 16'h0016; 
        10'b0001101110: data <= 16'hfff0; 
        10'b0001101111: data <= 16'h0014; 
        10'b0001110000: data <= 16'h0005; 
        10'b0001110001: data <= 16'hfff9; 
        10'b0001110010: data <= 16'hfffe; 
        10'b0001110011: data <= 16'h001f; 
        10'b0001110100: data <= 16'h001b; 
        10'b0001110101: data <= 16'h000a; 
        10'b0001110110: data <= 16'h000a; 
        10'b0001110111: data <= 16'h003f; 
        10'b0001111000: data <= 16'hfff9; 
        10'b0001111001: data <= 16'hfff3; 
        10'b0001111010: data <= 16'h003d; 
        10'b0001111011: data <= 16'h0017; 
        10'b0001111100: data <= 16'h001c; 
        10'b0001111101: data <= 16'h000a; 
        10'b0001111110: data <= 16'h0018; 
        10'b0001111111: data <= 16'h0024; 
        10'b0010000000: data <= 16'h007b; 
        10'b0010000001: data <= 16'h007a; 
        10'b0010000010: data <= 16'h00bf; 
        10'b0010000011: data <= 16'h00c2; 
        10'b0010000100: data <= 16'h00f5; 
        10'b0010000101: data <= 16'h0110; 
        10'b0010000110: data <= 16'h00ea; 
        10'b0010000111: data <= 16'h009d; 
        10'b0010001000: data <= 16'h0016; 
        10'b0010001001: data <= 16'h002a; 
        10'b0010001010: data <= 16'h0006; 
        10'b0010001011: data <= 16'h0000; 
        10'b0010001100: data <= 16'h0006; 
        10'b0010001101: data <= 16'h0013; 
        10'b0010001110: data <= 16'h000b; 
        10'b0010001111: data <= 16'hfff2; 
        10'b0010010000: data <= 16'hffe6; 
        10'b0010010001: data <= 16'hfffd; 
        10'b0010010010: data <= 16'hffea; 
        10'b0010010011: data <= 16'hffd5; 
        10'b0010010100: data <= 16'h0020; 
        10'b0010010101: data <= 16'hffd6; 
        10'b0010010110: data <= 16'h000f; 
        10'b0010010111: data <= 16'hff71; 
        10'b0010011000: data <= 16'hffb4; 
        10'b0010011001: data <= 16'hffcc; 
        10'b0010011010: data <= 16'hffed; 
        10'b0010011011: data <= 16'hffbd; 
        10'b0010011100: data <= 16'hffbd; 
        10'b0010011101: data <= 16'h000d; 
        10'b0010011110: data <= 16'h005c; 
        10'b0010011111: data <= 16'h00ac; 
        10'b0010100000: data <= 16'h0095; 
        10'b0010100001: data <= 16'h0085; 
        10'b0010100010: data <= 16'h0069; 
        10'b0010100011: data <= 16'h0048; 
        10'b0010100100: data <= 16'hfff8; 
        10'b0010100101: data <= 16'h0004; 
        10'b0010100110: data <= 16'hffdc; 
        10'b0010100111: data <= 16'h0022; 
        10'b0010101000: data <= 16'hfffb; 
        10'b0010101001: data <= 16'h001f; 
        10'b0010101010: data <= 16'h001d; 
        10'b0010101011: data <= 16'hffdb; 
        10'b0010101100: data <= 16'h000d; 
        10'b0010101101: data <= 16'hfffa; 
        10'b0010101110: data <= 16'h000c; 
        10'b0010101111: data <= 16'h0001; 
        10'b0010110000: data <= 16'hffcb; 
        10'b0010110001: data <= 16'hffbf; 
        10'b0010110010: data <= 16'hff5c; 
        10'b0010110011: data <= 16'hff29; 
        10'b0010110100: data <= 16'hff83; 
        10'b0010110101: data <= 16'hff0b; 
        10'b0010110110: data <= 16'hff94; 
        10'b0010110111: data <= 16'hffb1; 
        10'b0010111000: data <= 16'hff8f; 
        10'b0010111001: data <= 16'hff9c; 
        10'b0010111010: data <= 16'hffe4; 
        10'b0010111011: data <= 16'hffbd; 
        10'b0010111100: data <= 16'hff93; 
        10'b0010111101: data <= 16'hff98; 
        10'b0010111110: data <= 16'hff5f; 
        10'b0010111111: data <= 16'hff97; 
        10'b0011000000: data <= 16'hffa9; 
        10'b0011000001: data <= 16'hffa4; 
        10'b0011000010: data <= 16'hfff2; 
        10'b0011000011: data <= 16'h001e; 
        10'b0011000100: data <= 16'h000c; 
        10'b0011000101: data <= 16'h0012; 
        10'b0011000110: data <= 16'h0001; 
        10'b0011000111: data <= 16'hfffa; 
        10'b0011001000: data <= 16'h0002; 
        10'b0011001001: data <= 16'hffe0; 
        10'b0011001010: data <= 16'hffbf; 
        10'b0011001011: data <= 16'hfff6; 
        10'b0011001100: data <= 16'hffa4; 
        10'b0011001101: data <= 16'hff8e; 
        10'b0011001110: data <= 16'hff5a; 
        10'b0011001111: data <= 16'hff7e; 
        10'b0011010000: data <= 16'hff16; 
        10'b0011010001: data <= 16'hfefa; 
        10'b0011010010: data <= 16'hff77; 
        10'b0011010011: data <= 16'hff7e; 
        10'b0011010100: data <= 16'hff34; 
        10'b0011010101: data <= 16'hff3f; 
        10'b0011010110: data <= 16'hff10; 
        10'b0011010111: data <= 16'hfebb; 
        10'b0011011000: data <= 16'hfeb4; 
        10'b0011011001: data <= 16'hfeea; 
        10'b0011011010: data <= 16'hfedd; 
        10'b0011011011: data <= 16'hff1a; 
        10'b0011011100: data <= 16'hffa8; 
        10'b0011011101: data <= 16'hffb1; 
        10'b0011011110: data <= 16'hffe1; 
        10'b0011011111: data <= 16'hffe8; 
        10'b0011100000: data <= 16'hfff4; 
        10'b0011100001: data <= 16'hfff6; 
        10'b0011100010: data <= 16'h0023; 
        10'b0011100011: data <= 16'hffd3; 
        10'b0011100100: data <= 16'hffdb; 
        10'b0011100101: data <= 16'hffce; 
        10'b0011100110: data <= 16'hff83; 
        10'b0011100111: data <= 16'hffe5; 
        10'b0011101000: data <= 16'hffd2; 
        10'b0011101001: data <= 16'hff7e; 
        10'b0011101010: data <= 16'hff68; 
        10'b0011101011: data <= 16'hff51; 
        10'b0011101100: data <= 16'hff2e; 
        10'b0011101101: data <= 16'hff0c; 
        10'b0011101110: data <= 16'hff12; 
        10'b0011101111: data <= 16'hff02; 
        10'b0011110000: data <= 16'hfed3; 
        10'b0011110001: data <= 16'hfea5; 
        10'b0011110010: data <= 16'hfe16; 
        10'b0011110011: data <= 16'hfe38; 
        10'b0011110100: data <= 16'hfe68; 
        10'b0011110101: data <= 16'hfe6c; 
        10'b0011110110: data <= 16'hfee6; 
        10'b0011110111: data <= 16'hff08; 
        10'b0011111000: data <= 16'hff65; 
        10'b0011111001: data <= 16'hff9e; 
        10'b0011111010: data <= 16'hffba; 
        10'b0011111011: data <= 16'h000a; 
        10'b0011111100: data <= 16'hfffb; 
        10'b0011111101: data <= 16'hffe5; 
        10'b0011111110: data <= 16'hfff0; 
        10'b0011111111: data <= 16'hffe1; 
        10'b0100000000: data <= 16'h0001; 
        10'b0100000001: data <= 16'hffe3; 
        10'b0100000010: data <= 16'hffd4; 
        10'b0100000011: data <= 16'hffe7; 
        10'b0100000100: data <= 16'h001e; 
        10'b0100000101: data <= 16'hffb1; 
        10'b0100000110: data <= 16'hff6b; 
        10'b0100000111: data <= 16'hff8e; 
        10'b0100001000: data <= 16'hffb6; 
        10'b0100001001: data <= 16'hff75; 
        10'b0100001010: data <= 16'hff81; 
        10'b0100001011: data <= 16'hfeea; 
        10'b0100001100: data <= 16'hfebc; 
        10'b0100001101: data <= 16'hfe2b; 
        10'b0100001110: data <= 16'hfe0b; 
        10'b0100001111: data <= 16'hfe67; 
        10'b0100010000: data <= 16'hfeb1; 
        10'b0100010001: data <= 16'hfef5; 
        10'b0100010010: data <= 16'hfecb; 
        10'b0100010011: data <= 16'hff39; 
        10'b0100010100: data <= 16'hff69; 
        10'b0100010101: data <= 16'hff90; 
        10'b0100010110: data <= 16'hffd2; 
        10'b0100010111: data <= 16'h0018; 
        10'b0100011000: data <= 16'hffe8; 
        10'b0100011001: data <= 16'h001f; 
        10'b0100011010: data <= 16'h0015; 
        10'b0100011011: data <= 16'hffdc; 
        10'b0100011100: data <= 16'hffcc; 
        10'b0100011101: data <= 16'h000d; 
        10'b0100011110: data <= 16'h002b; 
        10'b0100011111: data <= 16'h002a; 
        10'b0100100000: data <= 16'h0098; 
        10'b0100100001: data <= 16'hfffd; 
        10'b0100100010: data <= 16'h001e; 
        10'b0100100011: data <= 16'h000d; 
        10'b0100100100: data <= 16'hffa4; 
        10'b0100100101: data <= 16'hffc2; 
        10'b0100100110: data <= 16'hff77; 
        10'b0100100111: data <= 16'hfee0; 
        10'b0100101000: data <= 16'hfedb; 
        10'b0100101001: data <= 16'hfea9; 
        10'b0100101010: data <= 16'hfe9b; 
        10'b0100101011: data <= 16'hfee3; 
        10'b0100101100: data <= 16'hff3e; 
        10'b0100101101: data <= 16'hff75; 
        10'b0100101110: data <= 16'hff4a; 
        10'b0100101111: data <= 16'hffed; 
        10'b0100110000: data <= 16'hff89; 
        10'b0100110001: data <= 16'hffad; 
        10'b0100110010: data <= 16'hffe7; 
        10'b0100110011: data <= 16'hfff4; 
        10'b0100110100: data <= 16'hffed; 
        10'b0100110101: data <= 16'h000c; 
        10'b0100110110: data <= 16'hffeb; 
        10'b0100110111: data <= 16'hfffd; 
        10'b0100111000: data <= 16'hffeb; 
        10'b0100111001: data <= 16'h0005; 
        10'b0100111010: data <= 16'hfff5; 
        10'b0100111011: data <= 16'h007f; 
        10'b0100111100: data <= 16'h005b; 
        10'b0100111101: data <= 16'h002c; 
        10'b0100111110: data <= 16'h0037; 
        10'b0100111111: data <= 16'h0027; 
        10'b0101000000: data <= 16'h0027; 
        10'b0101000001: data <= 16'h0006; 
        10'b0101000010: data <= 16'hffbe; 
        10'b0101000011: data <= 16'hff1c; 
        10'b0101000100: data <= 16'hff2a; 
        10'b0101000101: data <= 16'hff4a; 
        10'b0101000110: data <= 16'hff49; 
        10'b0101000111: data <= 16'hff72; 
        10'b0101001000: data <= 16'hffbd; 
        10'b0101001001: data <= 16'h001a; 
        10'b0101001010: data <= 16'h0057; 
        10'b0101001011: data <= 16'h0088; 
        10'b0101001100: data <= 16'h0000; 
        10'b0101001101: data <= 16'hffb8; 
        10'b0101001110: data <= 16'hffe2; 
        10'b0101001111: data <= 16'hfff5; 
        10'b0101010000: data <= 16'hffed; 
        10'b0101010001: data <= 16'hfff6; 
        10'b0101010010: data <= 16'hffe1; 
        10'b0101010011: data <= 16'hfff1; 
        10'b0101010100: data <= 16'h0012; 
        10'b0101010101: data <= 16'h003c; 
        10'b0101010110: data <= 16'h005b; 
        10'b0101010111: data <= 16'h0077; 
        10'b0101011000: data <= 16'h0037; 
        10'b0101011001: data <= 16'h004d; 
        10'b0101011010: data <= 16'h0037; 
        10'b0101011011: data <= 16'h0090; 
        10'b0101011100: data <= 16'h008a; 
        10'b0101011101: data <= 16'h0063; 
        10'b0101011110: data <= 16'hffab; 
        10'b0101011111: data <= 16'hff67; 
        10'b0101100000: data <= 16'hfffa; 
        10'b0101100001: data <= 16'hfff2; 
        10'b0101100010: data <= 16'hff6a; 
        10'b0101100011: data <= 16'hff70; 
        10'b0101100100: data <= 16'hffee; 
        10'b0101100101: data <= 16'h0051; 
        10'b0101100110: data <= 16'h00c4; 
        10'b0101100111: data <= 16'h015c; 
        10'b0101101000: data <= 16'h00bb; 
        10'b0101101001: data <= 16'hffcb; 
        10'b0101101010: data <= 16'hffc3; 
        10'b0101101011: data <= 16'hffed; 
        10'b0101101100: data <= 16'hffee; 
        10'b0101101101: data <= 16'h0020; 
        10'b0101101110: data <= 16'h0019; 
        10'b0101101111: data <= 16'hffdd; 
        10'b0101110000: data <= 16'hffd0; 
        10'b0101110001: data <= 16'h0013; 
        10'b0101110010: data <= 16'h0097; 
        10'b0101110011: data <= 16'h0051; 
        10'b0101110100: data <= 16'h0046; 
        10'b0101110101: data <= 16'h0022; 
        10'b0101110110: data <= 16'h0092; 
        10'b0101110111: data <= 16'h007a; 
        10'b0101111000: data <= 16'h0070; 
        10'b0101111001: data <= 16'h0014; 
        10'b0101111010: data <= 16'hffeb; 
        10'b0101111011: data <= 16'hfffc; 
        10'b0101111100: data <= 16'h000b; 
        10'b0101111101: data <= 16'hffdf; 
        10'b0101111110: data <= 16'hff7e; 
        10'b0101111111: data <= 16'hffef; 
        10'b0110000000: data <= 16'hffc1; 
        10'b0110000001: data <= 16'h0068; 
        10'b0110000010: data <= 16'h010f; 
        10'b0110000011: data <= 16'h01ae; 
        10'b0110000100: data <= 16'h00e8; 
        10'b0110000101: data <= 16'hffed; 
        10'b0110000110: data <= 16'h0001; 
        10'b0110000111: data <= 16'h0015; 
        10'b0110001000: data <= 16'hfff1; 
        10'b0110001001: data <= 16'h0003; 
        10'b0110001010: data <= 16'h0018; 
        10'b0110001011: data <= 16'h0001; 
        10'b0110001100: data <= 16'hffcd; 
        10'b0110001101: data <= 16'h0036; 
        10'b0110001110: data <= 16'h008a; 
        10'b0110001111: data <= 16'h0077; 
        10'b0110010000: data <= 16'h00a4; 
        10'b0110010001: data <= 16'h009a; 
        10'b0110010010: data <= 16'h00a6; 
        10'b0110010011: data <= 16'h00b4; 
        10'b0110010100: data <= 16'h003d; 
        10'b0110010101: data <= 16'hffa8; 
        10'b0110010110: data <= 16'h0006; 
        10'b0110010111: data <= 16'h0049; 
        10'b0110011000: data <= 16'h0023; 
        10'b0110011001: data <= 16'hffc7; 
        10'b0110011010: data <= 16'hffc8; 
        10'b0110011011: data <= 16'hfff8; 
        10'b0110011100: data <= 16'h0076; 
        10'b0110011101: data <= 16'h0074; 
        10'b0110011110: data <= 16'h0133; 
        10'b0110011111: data <= 16'h0166; 
        10'b0110100000: data <= 16'h00ea; 
        10'b0110100001: data <= 16'hfffd; 
        10'b0110100010: data <= 16'hffbd; 
        10'b0110100011: data <= 16'hffdf; 
        10'b0110100100: data <= 16'h0019; 
        10'b0110100101: data <= 16'hfff3; 
        10'b0110100110: data <= 16'h0005; 
        10'b0110100111: data <= 16'hffe4; 
        10'b0110101000: data <= 16'hff9f; 
        10'b0110101001: data <= 16'hfff4; 
        10'b0110101010: data <= 16'h0090; 
        10'b0110101011: data <= 16'h00c0; 
        10'b0110101100: data <= 16'h007c; 
        10'b0110101101: data <= 16'h00c2; 
        10'b0110101110: data <= 16'h00f4; 
        10'b0110101111: data <= 16'h012a; 
        10'b0110110000: data <= 16'h004e; 
        10'b0110110001: data <= 16'hffea; 
        10'b0110110010: data <= 16'h0073; 
        10'b0110110011: data <= 16'h006a; 
        10'b0110110100: data <= 16'h0010; 
        10'b0110110101: data <= 16'hffca; 
        10'b0110110110: data <= 16'h000b; 
        10'b0110110111: data <= 16'h003b; 
        10'b0110111000: data <= 16'h008a; 
        10'b0110111001: data <= 16'h00bd; 
        10'b0110111010: data <= 16'h00ae; 
        10'b0110111011: data <= 16'h00d7; 
        10'b0110111100: data <= 16'h0073; 
        10'b0110111101: data <= 16'hffc5; 
        10'b0110111110: data <= 16'hffdb; 
        10'b0110111111: data <= 16'hffda; 
        10'b0111000000: data <= 16'h0007; 
        10'b0111000001: data <= 16'hffe5; 
        10'b0111000010: data <= 16'hffe4; 
        10'b0111000011: data <= 16'hffe1; 
        10'b0111000100: data <= 16'hff80; 
        10'b0111000101: data <= 16'hffba; 
        10'b0111000110: data <= 16'h00d6; 
        10'b0111000111: data <= 16'h00da; 
        10'b0111001000: data <= 16'h0091; 
        10'b0111001001: data <= 16'h00df; 
        10'b0111001010: data <= 16'h017a; 
        10'b0111001011: data <= 16'h0177; 
        10'b0111001100: data <= 16'h0072; 
        10'b0111001101: data <= 16'h0044; 
        10'b0111001110: data <= 16'h00a3; 
        10'b0111001111: data <= 16'h0056; 
        10'b0111010000: data <= 16'hffd3; 
        10'b0111010001: data <= 16'hffa7; 
        10'b0111010010: data <= 16'h001f; 
        10'b0111010011: data <= 16'h005f; 
        10'b0111010100: data <= 16'h002c; 
        10'b0111010101: data <= 16'h0001; 
        10'b0111010110: data <= 16'h0059; 
        10'b0111010111: data <= 16'h0035; 
        10'b0111011000: data <= 16'hffe6; 
        10'b0111011001: data <= 16'hffbb; 
        10'b0111011010: data <= 16'hffd5; 
        10'b0111011011: data <= 16'hfffa; 
        10'b0111011100: data <= 16'h0006; 
        10'b0111011101: data <= 16'h0015; 
        10'b0111011110: data <= 16'h001d; 
        10'b0111011111: data <= 16'hfffb; 
        10'b0111100000: data <= 16'hff49; 
        10'b0111100001: data <= 16'hffa0; 
        10'b0111100010: data <= 16'h0059; 
        10'b0111100011: data <= 16'h00aa; 
        10'b0111100100: data <= 16'h00c1; 
        10'b0111100101: data <= 16'h00f4; 
        10'b0111100110: data <= 16'h01a5; 
        10'b0111100111: data <= 16'h01ac; 
        10'b0111101000: data <= 16'h00dd; 
        10'b0111101001: data <= 16'h007c; 
        10'b0111101010: data <= 16'h007e; 
        10'b0111101011: data <= 16'h004f; 
        10'b0111101100: data <= 16'h0000; 
        10'b0111101101: data <= 16'h0017; 
        10'b0111101110: data <= 16'h00af; 
        10'b0111101111: data <= 16'h003c; 
        10'b0111110000: data <= 16'h0019; 
        10'b0111110001: data <= 16'hffd3; 
        10'b0111110010: data <= 16'h0028; 
        10'b0111110011: data <= 16'hfff7; 
        10'b0111110100: data <= 16'hffce; 
        10'b0111110101: data <= 16'hff9f; 
        10'b0111110110: data <= 16'hfff2; 
        10'b0111110111: data <= 16'h0010; 
        10'b0111111000: data <= 16'hfff2; 
        10'b0111111001: data <= 16'hffec; 
        10'b0111111010: data <= 16'hffff; 
        10'b0111111011: data <= 16'hffcb; 
        10'b0111111100: data <= 16'hff54; 
        10'b0111111101: data <= 16'hff59; 
        10'b0111111110: data <= 16'hffaf; 
        10'b0111111111: data <= 16'h0075; 
        10'b1000000000: data <= 16'h00bb; 
        10'b1000000001: data <= 16'h00aa; 
        10'b1000000010: data <= 16'h0127; 
        10'b1000000011: data <= 16'h016b; 
        10'b1000000100: data <= 16'h01ac; 
        10'b1000000101: data <= 16'h00c7; 
        10'b1000000110: data <= 16'h0036; 
        10'b1000000111: data <= 16'h006f; 
        10'b1000001000: data <= 16'h00bf; 
        10'b1000001001: data <= 16'h007c; 
        10'b1000001010: data <= 16'h009a; 
        10'b1000001011: data <= 16'h0051; 
        10'b1000001100: data <= 16'h000a; 
        10'b1000001101: data <= 16'h001b; 
        10'b1000001110: data <= 16'h001e; 
        10'b1000001111: data <= 16'hffef; 
        10'b1000010000: data <= 16'hffc3; 
        10'b1000010001: data <= 16'hffd3; 
        10'b1000010010: data <= 16'hffdd; 
        10'b1000010011: data <= 16'hffdb; 
        10'b1000010100: data <= 16'h0009; 
        10'b1000010101: data <= 16'hffe6; 
        10'b1000010110: data <= 16'h0010; 
        10'b1000010111: data <= 16'hffbc; 
        10'b1000011000: data <= 16'hff91; 
        10'b1000011001: data <= 16'hff4e; 
        10'b1000011010: data <= 16'hff76; 
        10'b1000011011: data <= 16'h000a; 
        10'b1000011100: data <= 16'h007a; 
        10'b1000011101: data <= 16'h00bf; 
        10'b1000011110: data <= 16'h00fe; 
        10'b1000011111: data <= 16'h0195; 
        10'b1000100000: data <= 16'h01c8; 
        10'b1000100001: data <= 16'h00eb; 
        10'b1000100010: data <= 16'h00d2; 
        10'b1000100011: data <= 16'h00db; 
        10'b1000100100: data <= 16'h009c; 
        10'b1000100101: data <= 16'h0080; 
        10'b1000100110: data <= 16'h00c8; 
        10'b1000100111: data <= 16'h0088; 
        10'b1000101000: data <= 16'h0058; 
        10'b1000101001: data <= 16'h0013; 
        10'b1000101010: data <= 16'hffe0; 
        10'b1000101011: data <= 16'hffd9; 
        10'b1000101100: data <= 16'hffd7; 
        10'b1000101101: data <= 16'hfff9; 
        10'b1000101110: data <= 16'hffec; 
        10'b1000101111: data <= 16'h001d; 
        10'b1000110000: data <= 16'hffee; 
        10'b1000110001: data <= 16'hffe6; 
        10'b1000110010: data <= 16'hfff7; 
        10'b1000110011: data <= 16'hffe1; 
        10'b1000110100: data <= 16'hff72; 
        10'b1000110101: data <= 16'hff56; 
        10'b1000110110: data <= 16'hff6d; 
        10'b1000110111: data <= 16'hffc4; 
        10'b1000111000: data <= 16'h0028; 
        10'b1000111001: data <= 16'h0080; 
        10'b1000111010: data <= 16'h00d2; 
        10'b1000111011: data <= 16'h008c; 
        10'b1000111100: data <= 16'h0114; 
        10'b1000111101: data <= 16'h014b; 
        10'b1000111110: data <= 16'h0189; 
        10'b1000111111: data <= 16'h014f; 
        10'b1001000000: data <= 16'h00b5; 
        10'b1001000001: data <= 16'h0074; 
        10'b1001000010: data <= 16'h00e1; 
        10'b1001000011: data <= 16'h009f; 
        10'b1001000100: data <= 16'h006c; 
        10'b1001000101: data <= 16'hffea; 
        10'b1001000110: data <= 16'hffad; 
        10'b1001000111: data <= 16'h0005; 
        10'b1001001000: data <= 16'hffec; 
        10'b1001001001: data <= 16'hfff6; 
        10'b1001001010: data <= 16'hffe7; 
        10'b1001001011: data <= 16'h0005; 
        10'b1001001100: data <= 16'hfffd; 
        10'b1001001101: data <= 16'h0003; 
        10'b1001001110: data <= 16'h000b; 
        10'b1001001111: data <= 16'hfff5; 
        10'b1001010000: data <= 16'hffca; 
        10'b1001010001: data <= 16'hff8b; 
        10'b1001010010: data <= 16'hff39; 
        10'b1001010011: data <= 16'hffa6; 
        10'b1001010100: data <= 16'hffca; 
        10'b1001010101: data <= 16'h0060; 
        10'b1001010110: data <= 16'h00af; 
        10'b1001010111: data <= 16'h00f8; 
        10'b1001011000: data <= 16'h013f; 
        10'b1001011001: data <= 16'h0144; 
        10'b1001011010: data <= 16'h0110; 
        10'b1001011011: data <= 16'h00eb; 
        10'b1001011100: data <= 16'h0093; 
        10'b1001011101: data <= 16'h00c8; 
        10'b1001011110: data <= 16'h00bb; 
        10'b1001011111: data <= 16'h0077; 
        10'b1001100000: data <= 16'h0010; 
        10'b1001100001: data <= 16'hffc1; 
        10'b1001100010: data <= 16'hffa7; 
        10'b1001100011: data <= 16'hffcc; 
        10'b1001100100: data <= 16'h0003; 
        10'b1001100101: data <= 16'hffdf; 
        10'b1001100110: data <= 16'hfff9; 
        10'b1001100111: data <= 16'hffed; 
        10'b1001101000: data <= 16'hffed; 
        10'b1001101001: data <= 16'hfffd; 
        10'b1001101010: data <= 16'h0020; 
        10'b1001101011: data <= 16'h0009; 
        10'b1001101100: data <= 16'hffed; 
        10'b1001101101: data <= 16'hff9a; 
        10'b1001101110: data <= 16'hff87; 
        10'b1001101111: data <= 16'hff5e; 
        10'b1001110000: data <= 16'hff94; 
        10'b1001110001: data <= 16'hffcf; 
        10'b1001110010: data <= 16'hffd8; 
        10'b1001110011: data <= 16'h0014; 
        10'b1001110100: data <= 16'h005d; 
        10'b1001110101: data <= 16'h0028; 
        10'b1001110110: data <= 16'h0022; 
        10'b1001110111: data <= 16'h0065; 
        10'b1001111000: data <= 16'h004b; 
        10'b1001111001: data <= 16'h0001; 
        10'b1001111010: data <= 16'hffe7; 
        10'b1001111011: data <= 16'hff8f; 
        10'b1001111100: data <= 16'hff94; 
        10'b1001111101: data <= 16'hffa6; 
        10'b1001111110: data <= 16'hffac; 
        10'b1001111111: data <= 16'hfff8; 
        10'b1010000000: data <= 16'hfff1; 
        10'b1010000001: data <= 16'hffe1; 
        10'b1010000010: data <= 16'h0022; 
        10'b1010000011: data <= 16'h000d; 
        10'b1010000100: data <= 16'h001c; 
        10'b1010000101: data <= 16'hfff5; 
        10'b1010000110: data <= 16'hfff1; 
        10'b1010000111: data <= 16'h0003; 
        10'b1010001000: data <= 16'h000a; 
        10'b1010001001: data <= 16'hffd6; 
        10'b1010001010: data <= 16'hffbe; 
        10'b1010001011: data <= 16'hff6f; 
        10'b1010001100: data <= 16'hff49; 
        10'b1010001101: data <= 16'hfef9; 
        10'b1010001110: data <= 16'hfefa; 
        10'b1010001111: data <= 16'hfecf; 
        10'b1010010000: data <= 16'hff44; 
        10'b1010010001: data <= 16'hff6c; 
        10'b1010010010: data <= 16'hff8c; 
        10'b1010010011: data <= 16'hff54; 
        10'b1010010100: data <= 16'hff1e; 
        10'b1010010101: data <= 16'hff00; 
        10'b1010010110: data <= 16'hff36; 
        10'b1010010111: data <= 16'hffa4; 
        10'b1010011000: data <= 16'hffa2; 
        10'b1010011001: data <= 16'hffae; 
        10'b1010011010: data <= 16'hffe3; 
        10'b1010011011: data <= 16'h0004; 
        10'b1010011100: data <= 16'hffde; 
        10'b1010011101: data <= 16'hffe4; 
        10'b1010011110: data <= 16'hfff4; 
        10'b1010011111: data <= 16'hfffd; 
        10'b1010100000: data <= 16'h0014; 
        10'b1010100001: data <= 16'h0010; 
        10'b1010100010: data <= 16'h000b; 
        10'b1010100011: data <= 16'hffe0; 
        10'b1010100100: data <= 16'hffe6; 
        10'b1010100101: data <= 16'hfff4; 
        10'b1010100110: data <= 16'hffe1; 
        10'b1010100111: data <= 16'hffce; 
        10'b1010101000: data <= 16'hffd8; 
        10'b1010101001: data <= 16'hffc0; 
        10'b1010101010: data <= 16'hffa0; 
        10'b1010101011: data <= 16'hff87; 
        10'b1010101100: data <= 16'hff73; 
        10'b1010101101: data <= 16'hff76; 
        10'b1010101110: data <= 16'hff5f; 
        10'b1010101111: data <= 16'hff60; 
        10'b1010110000: data <= 16'hff58; 
        10'b1010110001: data <= 16'hff80; 
        10'b1010110010: data <= 16'hffd4; 
        10'b1010110011: data <= 16'hffd7; 
        10'b1010110100: data <= 16'hfff2; 
        10'b1010110101: data <= 16'hffe9; 
        10'b1010110110: data <= 16'h0011; 
        10'b1010110111: data <= 16'hfff9; 
        10'b1010111000: data <= 16'hffdf; 
        10'b1010111001: data <= 16'hfff5; 
        10'b1010111010: data <= 16'hffe7; 
        10'b1010111011: data <= 16'hffe8; 
        10'b1010111100: data <= 16'h001f; 
        10'b1010111101: data <= 16'hffe3; 
        10'b1010111110: data <= 16'h0009; 
        10'b1010111111: data <= 16'hfff1; 
        10'b1011000000: data <= 16'hffe9; 
        10'b1011000001: data <= 16'hfffc; 
        10'b1011000010: data <= 16'h0015; 
        10'b1011000011: data <= 16'hfffe; 
        10'b1011000100: data <= 16'hffdd; 
        10'b1011000101: data <= 16'h000d; 
        10'b1011000110: data <= 16'hffdd; 
        10'b1011000111: data <= 16'hfffb; 
        10'b1011001000: data <= 16'h0002; 
        10'b1011001001: data <= 16'hffdb; 
        10'b1011001010: data <= 16'hffec; 
        10'b1011001011: data <= 16'hfff4; 
        10'b1011001100: data <= 16'hfffd; 
        10'b1011001101: data <= 16'hffe0; 
        10'b1011001110: data <= 16'hffed; 
        10'b1011001111: data <= 16'hffdd; 
        10'b1011010000: data <= 16'hffe4; 
        10'b1011010001: data <= 16'h0004; 
        10'b1011010010: data <= 16'hfff3; 
        10'b1011010011: data <= 16'h0019; 
        10'b1011010100: data <= 16'h0024; 
        10'b1011010101: data <= 16'h0020; 
        10'b1011010110: data <= 16'h0001; 
        10'b1011010111: data <= 16'h0018; 
        10'b1011011000: data <= 16'h0022; 
        10'b1011011001: data <= 16'hfffe; 
        10'b1011011010: data <= 16'h0006; 
        10'b1011011011: data <= 16'hfffa; 
        10'b1011011100: data <= 16'hffed; 
        10'b1011011101: data <= 16'h001c; 
        10'b1011011110: data <= 16'h0015; 
        10'b1011011111: data <= 16'hffee; 
        10'b1011100000: data <= 16'hfff5; 
        10'b1011100001: data <= 16'h0010; 
        10'b1011100010: data <= 16'hfff3; 
        10'b1011100011: data <= 16'h0007; 
        10'b1011100100: data <= 16'hfff2; 
        10'b1011100101: data <= 16'h0015; 
        10'b1011100110: data <= 16'h0016; 
        10'b1011100111: data <= 16'hffe4; 
        10'b1011101000: data <= 16'hffea; 
        10'b1011101001: data <= 16'h001d; 
        10'b1011101010: data <= 16'h0017; 
        10'b1011101011: data <= 16'hfff5; 
        10'b1011101100: data <= 16'h0014; 
        10'b1011101101: data <= 16'hfff8; 
        10'b1011101110: data <= 16'hfff8; 
        10'b1011101111: data <= 16'h000d; 
        10'b1011110000: data <= 16'h000e; 
        10'b1011110001: data <= 16'hfff9; 
        10'b1011110010: data <= 16'hffef; 
        10'b1011110011: data <= 16'hfff6; 
        10'b1011110100: data <= 16'h0021; 
        10'b1011110101: data <= 16'hfffe; 
        10'b1011110110: data <= 16'h0012; 
        10'b1011110111: data <= 16'hffed; 
        10'b1011111000: data <= 16'h000b; 
        10'b1011111001: data <= 16'hffff; 
        10'b1011111010: data <= 16'h001f; 
        10'b1011111011: data <= 16'h0004; 
        10'b1011111100: data <= 16'hfffc; 
        10'b1011111101: data <= 16'hffdc; 
        10'b1011111110: data <= 16'hffe8; 
        10'b1011111111: data <= 16'h000b; 
        10'b1100000000: data <= 16'hffdf; 
        10'b1100000001: data <= 16'hffe5; 
        10'b1100000010: data <= 16'hffeb; 
        10'b1100000011: data <= 16'hffdf; 
        10'b1100000100: data <= 16'hffe9; 
        10'b1100000101: data <= 16'hfff5; 
        10'b1100000110: data <= 16'hffe2; 
        10'b1100000111: data <= 16'hffe9; 
        10'b1100001000: data <= 16'hffed; 
        10'b1100001001: data <= 16'hfff0; 
        10'b1100001010: data <= 16'h001e; 
        10'b1100001011: data <= 16'hffe3; 
        10'b1100001100: data <= 16'hffed; 
        10'b1100001101: data <= 16'hffe4; 
        10'b1100001110: data <= 16'hffec; 
        10'b1100001111: data <= 16'h0006; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 11) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 17'h1ffe9; 
        10'b0000000001: data <= 17'h0002e; 
        10'b0000000010: data <= 17'h1ffcc; 
        10'b0000000011: data <= 17'h1fffc; 
        10'b0000000100: data <= 17'h1fffe; 
        10'b0000000101: data <= 17'h1fff9; 
        10'b0000000110: data <= 17'h00018; 
        10'b0000000111: data <= 17'h0004a; 
        10'b0000001000: data <= 17'h1ffd0; 
        10'b0000001001: data <= 17'h1ffe0; 
        10'b0000001010: data <= 17'h1ffe2; 
        10'b0000001011: data <= 17'h1ffd2; 
        10'b0000001100: data <= 17'h00018; 
        10'b0000001101: data <= 17'h00043; 
        10'b0000001110: data <= 17'h00026; 
        10'b0000001111: data <= 17'h1ffc2; 
        10'b0000010000: data <= 17'h1fff8; 
        10'b0000010001: data <= 17'h0004a; 
        10'b0000010010: data <= 17'h0000c; 
        10'b0000010011: data <= 17'h1fff9; 
        10'b0000010100: data <= 17'h1ffc7; 
        10'b0000010101: data <= 17'h1ffda; 
        10'b0000010110: data <= 17'h00011; 
        10'b0000010111: data <= 17'h00041; 
        10'b0000011000: data <= 17'h00023; 
        10'b0000011001: data <= 17'h0002a; 
        10'b0000011010: data <= 17'h1ffc6; 
        10'b0000011011: data <= 17'h1ffc9; 
        10'b0000011100: data <= 17'h0002f; 
        10'b0000011101: data <= 17'h00026; 
        10'b0000011110: data <= 17'h00030; 
        10'b0000011111: data <= 17'h1fff4; 
        10'b0000100000: data <= 17'h1ffbf; 
        10'b0000100001: data <= 17'h1ffd9; 
        10'b0000100010: data <= 17'h00021; 
        10'b0000100011: data <= 17'h0006b; 
        10'b0000100100: data <= 17'h00049; 
        10'b0000100101: data <= 17'h00016; 
        10'b0000100110: data <= 17'h00058; 
        10'b0000100111: data <= 17'h0005e; 
        10'b0000101000: data <= 17'h00064; 
        10'b0000101001: data <= 17'h0005e; 
        10'b0000101010: data <= 17'h0003b; 
        10'b0000101011: data <= 17'h00040; 
        10'b0000101100: data <= 17'h1ffbc; 
        10'b0000101101: data <= 17'h0003d; 
        10'b0000101110: data <= 17'h00052; 
        10'b0000101111: data <= 17'h0002f; 
        10'b0000110000: data <= 17'h1fff3; 
        10'b0000110001: data <= 17'h1ffd6; 
        10'b0000110010: data <= 17'h00057; 
        10'b0000110011: data <= 17'h00042; 
        10'b0000110100: data <= 17'h1ffe5; 
        10'b0000110101: data <= 17'h00049; 
        10'b0000110110: data <= 17'h1fff3; 
        10'b0000110111: data <= 17'h00036; 
        10'b0000111000: data <= 17'h1ffd5; 
        10'b0000111001: data <= 17'h1ffcd; 
        10'b0000111010: data <= 17'h1ffbf; 
        10'b0000111011: data <= 17'h1fffa; 
        10'b0000111100: data <= 17'h00024; 
        10'b0000111101: data <= 17'h00016; 
        10'b0000111110: data <= 17'h00025; 
        10'b0000111111: data <= 17'h00069; 
        10'b0001000000: data <= 17'h0004b; 
        10'b0001000001: data <= 17'h0009f; 
        10'b0001000010: data <= 17'h000c8; 
        10'b0001000011: data <= 17'h000e2; 
        10'b0001000100: data <= 17'h000e3; 
        10'b0001000101: data <= 17'h000ee; 
        10'b0001000110: data <= 17'h00079; 
        10'b0001000111: data <= 17'h00056; 
        10'b0001001000: data <= 17'h000c7; 
        10'b0001001001: data <= 17'h00058; 
        10'b0001001010: data <= 17'h00055; 
        10'b0001001011: data <= 17'h0005d; 
        10'b0001001100: data <= 17'h0005b; 
        10'b0001001101: data <= 17'h0002e; 
        10'b0001001110: data <= 17'h0003d; 
        10'b0001001111: data <= 17'h0000b; 
        10'b0001010000: data <= 17'h00021; 
        10'b0001010001: data <= 17'h1ffed; 
        10'b0001010010: data <= 17'h1ffbd; 
        10'b0001010011: data <= 17'h00015; 
        10'b0001010100: data <= 17'h1ffc7; 
        10'b0001010101: data <= 17'h00007; 
        10'b0001010110: data <= 17'h00036; 
        10'b0001010111: data <= 17'h0001f; 
        10'b0001011000: data <= 17'h00047; 
        10'b0001011001: data <= 17'h1ffc2; 
        10'b0001011010: data <= 17'h0004d; 
        10'b0001011011: data <= 17'h00054; 
        10'b0001011100: data <= 17'h00064; 
        10'b0001011101: data <= 17'h000cb; 
        10'b0001011110: data <= 17'h000b4; 
        10'b0001011111: data <= 17'h000e1; 
        10'b0001100000: data <= 17'h000dc; 
        10'b0001100001: data <= 17'h000d3; 
        10'b0001100010: data <= 17'h00137; 
        10'b0001100011: data <= 17'h00125; 
        10'b0001100100: data <= 17'h000b6; 
        10'b0001100101: data <= 17'h000e6; 
        10'b0001100110: data <= 17'h00172; 
        10'b0001100111: data <= 17'h00171; 
        10'b0001101000: data <= 17'h00189; 
        10'b0001101001: data <= 17'h0015c; 
        10'b0001101010: data <= 17'h00161; 
        10'b0001101011: data <= 17'h000cd; 
        10'b0001101100: data <= 17'h000b6; 
        10'b0001101101: data <= 17'h0002c; 
        10'b0001101110: data <= 17'h1ffe1; 
        10'b0001101111: data <= 17'h00028; 
        10'b0001110000: data <= 17'h0000b; 
        10'b0001110001: data <= 17'h1fff3; 
        10'b0001110010: data <= 17'h1fffb; 
        10'b0001110011: data <= 17'h0003e; 
        10'b0001110100: data <= 17'h00036; 
        10'b0001110101: data <= 17'h00014; 
        10'b0001110110: data <= 17'h00014; 
        10'b0001110111: data <= 17'h0007e; 
        10'b0001111000: data <= 17'h1fff2; 
        10'b0001111001: data <= 17'h1ffe6; 
        10'b0001111010: data <= 17'h0007a; 
        10'b0001111011: data <= 17'h0002e; 
        10'b0001111100: data <= 17'h00038; 
        10'b0001111101: data <= 17'h00014; 
        10'b0001111110: data <= 17'h00030; 
        10'b0001111111: data <= 17'h00048; 
        10'b0010000000: data <= 17'h000f6; 
        10'b0010000001: data <= 17'h000f4; 
        10'b0010000010: data <= 17'h0017e; 
        10'b0010000011: data <= 17'h00185; 
        10'b0010000100: data <= 17'h001ea; 
        10'b0010000101: data <= 17'h00220; 
        10'b0010000110: data <= 17'h001d4; 
        10'b0010000111: data <= 17'h0013a; 
        10'b0010001000: data <= 17'h0002d; 
        10'b0010001001: data <= 17'h00053; 
        10'b0010001010: data <= 17'h0000c; 
        10'b0010001011: data <= 17'h00000; 
        10'b0010001100: data <= 17'h0000d; 
        10'b0010001101: data <= 17'h00026; 
        10'b0010001110: data <= 17'h00016; 
        10'b0010001111: data <= 17'h1ffe3; 
        10'b0010010000: data <= 17'h1ffcc; 
        10'b0010010001: data <= 17'h1fffa; 
        10'b0010010010: data <= 17'h1ffd5; 
        10'b0010010011: data <= 17'h1ffaa; 
        10'b0010010100: data <= 17'h00041; 
        10'b0010010101: data <= 17'h1ffad; 
        10'b0010010110: data <= 17'h0001e; 
        10'b0010010111: data <= 17'h1fee3; 
        10'b0010011000: data <= 17'h1ff69; 
        10'b0010011001: data <= 17'h1ff98; 
        10'b0010011010: data <= 17'h1ffda; 
        10'b0010011011: data <= 17'h1ff79; 
        10'b0010011100: data <= 17'h1ff79; 
        10'b0010011101: data <= 17'h0001a; 
        10'b0010011110: data <= 17'h000b7; 
        10'b0010011111: data <= 17'h00158; 
        10'b0010100000: data <= 17'h0012a; 
        10'b0010100001: data <= 17'h0010b; 
        10'b0010100010: data <= 17'h000d2; 
        10'b0010100011: data <= 17'h00090; 
        10'b0010100100: data <= 17'h1ffef; 
        10'b0010100101: data <= 17'h00007; 
        10'b0010100110: data <= 17'h1ffb7; 
        10'b0010100111: data <= 17'h00044; 
        10'b0010101000: data <= 17'h1fff7; 
        10'b0010101001: data <= 17'h0003e; 
        10'b0010101010: data <= 17'h00039; 
        10'b0010101011: data <= 17'h1ffb6; 
        10'b0010101100: data <= 17'h0001a; 
        10'b0010101101: data <= 17'h1fff4; 
        10'b0010101110: data <= 17'h00018; 
        10'b0010101111: data <= 17'h00002; 
        10'b0010110000: data <= 17'h1ff96; 
        10'b0010110001: data <= 17'h1ff7f; 
        10'b0010110010: data <= 17'h1feb7; 
        10'b0010110011: data <= 17'h1fe52; 
        10'b0010110100: data <= 17'h1ff06; 
        10'b0010110101: data <= 17'h1fe16; 
        10'b0010110110: data <= 17'h1ff28; 
        10'b0010110111: data <= 17'h1ff61; 
        10'b0010111000: data <= 17'h1ff1e; 
        10'b0010111001: data <= 17'h1ff38; 
        10'b0010111010: data <= 17'h1ffc9; 
        10'b0010111011: data <= 17'h1ff7a; 
        10'b0010111100: data <= 17'h1ff27; 
        10'b0010111101: data <= 17'h1ff31; 
        10'b0010111110: data <= 17'h1febe; 
        10'b0010111111: data <= 17'h1ff2e; 
        10'b0011000000: data <= 17'h1ff52; 
        10'b0011000001: data <= 17'h1ff48; 
        10'b0011000010: data <= 17'h1ffe5; 
        10'b0011000011: data <= 17'h0003c; 
        10'b0011000100: data <= 17'h00018; 
        10'b0011000101: data <= 17'h00024; 
        10'b0011000110: data <= 17'h00002; 
        10'b0011000111: data <= 17'h1fff4; 
        10'b0011001000: data <= 17'h00004; 
        10'b0011001001: data <= 17'h1ffc0; 
        10'b0011001010: data <= 17'h1ff7f; 
        10'b0011001011: data <= 17'h1ffeb; 
        10'b0011001100: data <= 17'h1ff49; 
        10'b0011001101: data <= 17'h1ff1c; 
        10'b0011001110: data <= 17'h1feb5; 
        10'b0011001111: data <= 17'h1fefc; 
        10'b0011010000: data <= 17'h1fe2c; 
        10'b0011010001: data <= 17'h1fdf4; 
        10'b0011010010: data <= 17'h1feed; 
        10'b0011010011: data <= 17'h1fefb; 
        10'b0011010100: data <= 17'h1fe67; 
        10'b0011010101: data <= 17'h1fe7d; 
        10'b0011010110: data <= 17'h1fe20; 
        10'b0011010111: data <= 17'h1fd75; 
        10'b0011011000: data <= 17'h1fd68; 
        10'b0011011001: data <= 17'h1fdd4; 
        10'b0011011010: data <= 17'h1fdbb; 
        10'b0011011011: data <= 17'h1fe35; 
        10'b0011011100: data <= 17'h1ff51; 
        10'b0011011101: data <= 17'h1ff61; 
        10'b0011011110: data <= 17'h1ffc1; 
        10'b0011011111: data <= 17'h1ffd0; 
        10'b0011100000: data <= 17'h1ffe9; 
        10'b0011100001: data <= 17'h1ffec; 
        10'b0011100010: data <= 17'h00046; 
        10'b0011100011: data <= 17'h1ffa6; 
        10'b0011100100: data <= 17'h1ffb5; 
        10'b0011100101: data <= 17'h1ff9d; 
        10'b0011100110: data <= 17'h1ff07; 
        10'b0011100111: data <= 17'h1ffc9; 
        10'b0011101000: data <= 17'h1ffa4; 
        10'b0011101001: data <= 17'h1fefb; 
        10'b0011101010: data <= 17'h1fecf; 
        10'b0011101011: data <= 17'h1fea3; 
        10'b0011101100: data <= 17'h1fe5c; 
        10'b0011101101: data <= 17'h1fe18; 
        10'b0011101110: data <= 17'h1fe25; 
        10'b0011101111: data <= 17'h1fe04; 
        10'b0011110000: data <= 17'h1fda6; 
        10'b0011110001: data <= 17'h1fd4b; 
        10'b0011110010: data <= 17'h1fc2c; 
        10'b0011110011: data <= 17'h1fc70; 
        10'b0011110100: data <= 17'h1fcd1; 
        10'b0011110101: data <= 17'h1fcd9; 
        10'b0011110110: data <= 17'h1fdcc; 
        10'b0011110111: data <= 17'h1fe0f; 
        10'b0011111000: data <= 17'h1feca; 
        10'b0011111001: data <= 17'h1ff3d; 
        10'b0011111010: data <= 17'h1ff74; 
        10'b0011111011: data <= 17'h00015; 
        10'b0011111100: data <= 17'h1fff6; 
        10'b0011111101: data <= 17'h1ffc9; 
        10'b0011111110: data <= 17'h1ffe1; 
        10'b0011111111: data <= 17'h1ffc2; 
        10'b0100000000: data <= 17'h00002; 
        10'b0100000001: data <= 17'h1ffc7; 
        10'b0100000010: data <= 17'h1ffa9; 
        10'b0100000011: data <= 17'h1ffce; 
        10'b0100000100: data <= 17'h0003c; 
        10'b0100000101: data <= 17'h1ff63; 
        10'b0100000110: data <= 17'h1fed6; 
        10'b0100000111: data <= 17'h1ff1c; 
        10'b0100001000: data <= 17'h1ff6d; 
        10'b0100001001: data <= 17'h1feeb; 
        10'b0100001010: data <= 17'h1ff02; 
        10'b0100001011: data <= 17'h1fdd4; 
        10'b0100001100: data <= 17'h1fd78; 
        10'b0100001101: data <= 17'h1fc56; 
        10'b0100001110: data <= 17'h1fc17; 
        10'b0100001111: data <= 17'h1fccf; 
        10'b0100010000: data <= 17'h1fd61; 
        10'b0100010001: data <= 17'h1fdeb; 
        10'b0100010010: data <= 17'h1fd96; 
        10'b0100010011: data <= 17'h1fe73; 
        10'b0100010100: data <= 17'h1fed1; 
        10'b0100010101: data <= 17'h1ff1f; 
        10'b0100010110: data <= 17'h1ffa4; 
        10'b0100010111: data <= 17'h00031; 
        10'b0100011000: data <= 17'h1ffd1; 
        10'b0100011001: data <= 17'h0003d; 
        10'b0100011010: data <= 17'h0002a; 
        10'b0100011011: data <= 17'h1ffb8; 
        10'b0100011100: data <= 17'h1ff97; 
        10'b0100011101: data <= 17'h0001b; 
        10'b0100011110: data <= 17'h00056; 
        10'b0100011111: data <= 17'h00053; 
        10'b0100100000: data <= 17'h00130; 
        10'b0100100001: data <= 17'h1fffa; 
        10'b0100100010: data <= 17'h0003c; 
        10'b0100100011: data <= 17'h00019; 
        10'b0100100100: data <= 17'h1ff48; 
        10'b0100100101: data <= 17'h1ff83; 
        10'b0100100110: data <= 17'h1feee; 
        10'b0100100111: data <= 17'h1fdc1; 
        10'b0100101000: data <= 17'h1fdb7; 
        10'b0100101001: data <= 17'h1fd52; 
        10'b0100101010: data <= 17'h1fd36; 
        10'b0100101011: data <= 17'h1fdc6; 
        10'b0100101100: data <= 17'h1fe7d; 
        10'b0100101101: data <= 17'h1feeb; 
        10'b0100101110: data <= 17'h1fe93; 
        10'b0100101111: data <= 17'h1ffda; 
        10'b0100110000: data <= 17'h1ff13; 
        10'b0100110001: data <= 17'h1ff5b; 
        10'b0100110010: data <= 17'h1ffcf; 
        10'b0100110011: data <= 17'h1ffe8; 
        10'b0100110100: data <= 17'h1ffda; 
        10'b0100110101: data <= 17'h00019; 
        10'b0100110110: data <= 17'h1ffd6; 
        10'b0100110111: data <= 17'h1fffa; 
        10'b0100111000: data <= 17'h1ffd6; 
        10'b0100111001: data <= 17'h0000b; 
        10'b0100111010: data <= 17'h1ffe9; 
        10'b0100111011: data <= 17'h000fe; 
        10'b0100111100: data <= 17'h000b6; 
        10'b0100111101: data <= 17'h00058; 
        10'b0100111110: data <= 17'h0006e; 
        10'b0100111111: data <= 17'h0004e; 
        10'b0101000000: data <= 17'h0004e; 
        10'b0101000001: data <= 17'h0000c; 
        10'b0101000010: data <= 17'h1ff7b; 
        10'b0101000011: data <= 17'h1fe38; 
        10'b0101000100: data <= 17'h1fe54; 
        10'b0101000101: data <= 17'h1fe94; 
        10'b0101000110: data <= 17'h1fe92; 
        10'b0101000111: data <= 17'h1fee3; 
        10'b0101001000: data <= 17'h1ff7b; 
        10'b0101001001: data <= 17'h00033; 
        10'b0101001010: data <= 17'h000af; 
        10'b0101001011: data <= 17'h00110; 
        10'b0101001100: data <= 17'h1ffff; 
        10'b0101001101: data <= 17'h1ff70; 
        10'b0101001110: data <= 17'h1ffc4; 
        10'b0101001111: data <= 17'h1ffea; 
        10'b0101010000: data <= 17'h1ffda; 
        10'b0101010001: data <= 17'h1ffeb; 
        10'b0101010010: data <= 17'h1ffc2; 
        10'b0101010011: data <= 17'h1ffe2; 
        10'b0101010100: data <= 17'h00024; 
        10'b0101010101: data <= 17'h00077; 
        10'b0101010110: data <= 17'h000b6; 
        10'b0101010111: data <= 17'h000ef; 
        10'b0101011000: data <= 17'h0006f; 
        10'b0101011001: data <= 17'h0009b; 
        10'b0101011010: data <= 17'h0006d; 
        10'b0101011011: data <= 17'h0011f; 
        10'b0101011100: data <= 17'h00115; 
        10'b0101011101: data <= 17'h000c6; 
        10'b0101011110: data <= 17'h1ff56; 
        10'b0101011111: data <= 17'h1fece; 
        10'b0101100000: data <= 17'h1fff3; 
        10'b0101100001: data <= 17'h1ffe4; 
        10'b0101100010: data <= 17'h1fed4; 
        10'b0101100011: data <= 17'h1fee1; 
        10'b0101100100: data <= 17'h1ffdc; 
        10'b0101100101: data <= 17'h000a2; 
        10'b0101100110: data <= 17'h00188; 
        10'b0101100111: data <= 17'h002b8; 
        10'b0101101000: data <= 17'h00176; 
        10'b0101101001: data <= 17'h1ff95; 
        10'b0101101010: data <= 17'h1ff85; 
        10'b0101101011: data <= 17'h1ffdb; 
        10'b0101101100: data <= 17'h1ffdc; 
        10'b0101101101: data <= 17'h00041; 
        10'b0101101110: data <= 17'h00031; 
        10'b0101101111: data <= 17'h1ffba; 
        10'b0101110000: data <= 17'h1ffa0; 
        10'b0101110001: data <= 17'h00027; 
        10'b0101110010: data <= 17'h0012e; 
        10'b0101110011: data <= 17'h000a2; 
        10'b0101110100: data <= 17'h0008c; 
        10'b0101110101: data <= 17'h00045; 
        10'b0101110110: data <= 17'h00125; 
        10'b0101110111: data <= 17'h000f5; 
        10'b0101111000: data <= 17'h000e0; 
        10'b0101111001: data <= 17'h00028; 
        10'b0101111010: data <= 17'h1ffd7; 
        10'b0101111011: data <= 17'h1fff9; 
        10'b0101111100: data <= 17'h00017; 
        10'b0101111101: data <= 17'h1ffbe; 
        10'b0101111110: data <= 17'h1fefb; 
        10'b0101111111: data <= 17'h1ffde; 
        10'b0110000000: data <= 17'h1ff82; 
        10'b0110000001: data <= 17'h000d1; 
        10'b0110000010: data <= 17'h0021f; 
        10'b0110000011: data <= 17'h0035c; 
        10'b0110000100: data <= 17'h001d1; 
        10'b0110000101: data <= 17'h1ffdb; 
        10'b0110000110: data <= 17'h00001; 
        10'b0110000111: data <= 17'h0002a; 
        10'b0110001000: data <= 17'h1ffe1; 
        10'b0110001001: data <= 17'h00007; 
        10'b0110001010: data <= 17'h00031; 
        10'b0110001011: data <= 17'h00003; 
        10'b0110001100: data <= 17'h1ff9a; 
        10'b0110001101: data <= 17'h0006c; 
        10'b0110001110: data <= 17'h00115; 
        10'b0110001111: data <= 17'h000ef; 
        10'b0110010000: data <= 17'h00148; 
        10'b0110010001: data <= 17'h00134; 
        10'b0110010010: data <= 17'h0014d; 
        10'b0110010011: data <= 17'h00168; 
        10'b0110010100: data <= 17'h00079; 
        10'b0110010101: data <= 17'h1ff50; 
        10'b0110010110: data <= 17'h0000c; 
        10'b0110010111: data <= 17'h00093; 
        10'b0110011000: data <= 17'h00046; 
        10'b0110011001: data <= 17'h1ff8e; 
        10'b0110011010: data <= 17'h1ff91; 
        10'b0110011011: data <= 17'h1fff0; 
        10'b0110011100: data <= 17'h000eb; 
        10'b0110011101: data <= 17'h000e9; 
        10'b0110011110: data <= 17'h00267; 
        10'b0110011111: data <= 17'h002cb; 
        10'b0110100000: data <= 17'h001d5; 
        10'b0110100001: data <= 17'h1fff9; 
        10'b0110100010: data <= 17'h1ff7a; 
        10'b0110100011: data <= 17'h1ffbe; 
        10'b0110100100: data <= 17'h00032; 
        10'b0110100101: data <= 17'h1ffe7; 
        10'b0110100110: data <= 17'h0000a; 
        10'b0110100111: data <= 17'h1ffc9; 
        10'b0110101000: data <= 17'h1ff3e; 
        10'b0110101001: data <= 17'h1ffe8; 
        10'b0110101010: data <= 17'h00121; 
        10'b0110101011: data <= 17'h00180; 
        10'b0110101100: data <= 17'h000f7; 
        10'b0110101101: data <= 17'h00184; 
        10'b0110101110: data <= 17'h001e9; 
        10'b0110101111: data <= 17'h00254; 
        10'b0110110000: data <= 17'h0009c; 
        10'b0110110001: data <= 17'h1ffd5; 
        10'b0110110010: data <= 17'h000e6; 
        10'b0110110011: data <= 17'h000d4; 
        10'b0110110100: data <= 17'h00021; 
        10'b0110110101: data <= 17'h1ff94; 
        10'b0110110110: data <= 17'h00016; 
        10'b0110110111: data <= 17'h00077; 
        10'b0110111000: data <= 17'h00113; 
        10'b0110111001: data <= 17'h0017a; 
        10'b0110111010: data <= 17'h0015b; 
        10'b0110111011: data <= 17'h001af; 
        10'b0110111100: data <= 17'h000e6; 
        10'b0110111101: data <= 17'h1ff8a; 
        10'b0110111110: data <= 17'h1ffb7; 
        10'b0110111111: data <= 17'h1ffb5; 
        10'b0111000000: data <= 17'h0000d; 
        10'b0111000001: data <= 17'h1ffc9; 
        10'b0111000010: data <= 17'h1ffc7; 
        10'b0111000011: data <= 17'h1ffc1; 
        10'b0111000100: data <= 17'h1ff00; 
        10'b0111000101: data <= 17'h1ff75; 
        10'b0111000110: data <= 17'h001ac; 
        10'b0111000111: data <= 17'h001b5; 
        10'b0111001000: data <= 17'h00121; 
        10'b0111001001: data <= 17'h001be; 
        10'b0111001010: data <= 17'h002f4; 
        10'b0111001011: data <= 17'h002ee; 
        10'b0111001100: data <= 17'h000e5; 
        10'b0111001101: data <= 17'h00088; 
        10'b0111001110: data <= 17'h00146; 
        10'b0111001111: data <= 17'h000ac; 
        10'b0111010000: data <= 17'h1ffa6; 
        10'b0111010001: data <= 17'h1ff4e; 
        10'b0111010010: data <= 17'h0003e; 
        10'b0111010011: data <= 17'h000bf; 
        10'b0111010100: data <= 17'h00059; 
        10'b0111010101: data <= 17'h00003; 
        10'b0111010110: data <= 17'h000b2; 
        10'b0111010111: data <= 17'h0006b; 
        10'b0111011000: data <= 17'h1ffcc; 
        10'b0111011001: data <= 17'h1ff75; 
        10'b0111011010: data <= 17'h1ffab; 
        10'b0111011011: data <= 17'h1fff4; 
        10'b0111011100: data <= 17'h0000d; 
        10'b0111011101: data <= 17'h0002a; 
        10'b0111011110: data <= 17'h0003a; 
        10'b0111011111: data <= 17'h1fff6; 
        10'b0111100000: data <= 17'h1fe92; 
        10'b0111100001: data <= 17'h1ff41; 
        10'b0111100010: data <= 17'h000b3; 
        10'b0111100011: data <= 17'h00154; 
        10'b0111100100: data <= 17'h00183; 
        10'b0111100101: data <= 17'h001e8; 
        10'b0111100110: data <= 17'h00349; 
        10'b0111100111: data <= 17'h00357; 
        10'b0111101000: data <= 17'h001ba; 
        10'b0111101001: data <= 17'h000f9; 
        10'b0111101010: data <= 17'h000fc; 
        10'b0111101011: data <= 17'h0009f; 
        10'b0111101100: data <= 17'h00000; 
        10'b0111101101: data <= 17'h0002e; 
        10'b0111101110: data <= 17'h0015e; 
        10'b0111101111: data <= 17'h00079; 
        10'b0111110000: data <= 17'h00032; 
        10'b0111110001: data <= 17'h1ffa7; 
        10'b0111110010: data <= 17'h00050; 
        10'b0111110011: data <= 17'h1ffef; 
        10'b0111110100: data <= 17'h1ff9c; 
        10'b0111110101: data <= 17'h1ff3e; 
        10'b0111110110: data <= 17'h1ffe4; 
        10'b0111110111: data <= 17'h00020; 
        10'b0111111000: data <= 17'h1ffe3; 
        10'b0111111001: data <= 17'h1ffd8; 
        10'b0111111010: data <= 17'h1ffff; 
        10'b0111111011: data <= 17'h1ff95; 
        10'b0111111100: data <= 17'h1fea9; 
        10'b0111111101: data <= 17'h1feb1; 
        10'b0111111110: data <= 17'h1ff5e; 
        10'b0111111111: data <= 17'h000ea; 
        10'b1000000000: data <= 17'h00176; 
        10'b1000000001: data <= 17'h00154; 
        10'b1000000010: data <= 17'h0024d; 
        10'b1000000011: data <= 17'h002d7; 
        10'b1000000100: data <= 17'h00358; 
        10'b1000000101: data <= 17'h0018e; 
        10'b1000000110: data <= 17'h0006c; 
        10'b1000000111: data <= 17'h000dd; 
        10'b1000001000: data <= 17'h0017e; 
        10'b1000001001: data <= 17'h000f8; 
        10'b1000001010: data <= 17'h00135; 
        10'b1000001011: data <= 17'h000a2; 
        10'b1000001100: data <= 17'h00015; 
        10'b1000001101: data <= 17'h00036; 
        10'b1000001110: data <= 17'h0003c; 
        10'b1000001111: data <= 17'h1ffde; 
        10'b1000010000: data <= 17'h1ff86; 
        10'b1000010001: data <= 17'h1ffa6; 
        10'b1000010010: data <= 17'h1ffba; 
        10'b1000010011: data <= 17'h1ffb6; 
        10'b1000010100: data <= 17'h00012; 
        10'b1000010101: data <= 17'h1ffcc; 
        10'b1000010110: data <= 17'h00021; 
        10'b1000010111: data <= 17'h1ff79; 
        10'b1000011000: data <= 17'h1ff22; 
        10'b1000011001: data <= 17'h1fe9b; 
        10'b1000011010: data <= 17'h1feeb; 
        10'b1000011011: data <= 17'h00014; 
        10'b1000011100: data <= 17'h000f3; 
        10'b1000011101: data <= 17'h0017e; 
        10'b1000011110: data <= 17'h001fc; 
        10'b1000011111: data <= 17'h0032a; 
        10'b1000100000: data <= 17'h00390; 
        10'b1000100001: data <= 17'h001d6; 
        10'b1000100010: data <= 17'h001a4; 
        10'b1000100011: data <= 17'h001b7; 
        10'b1000100100: data <= 17'h00138; 
        10'b1000100101: data <= 17'h00101; 
        10'b1000100110: data <= 17'h00191; 
        10'b1000100111: data <= 17'h00111; 
        10'b1000101000: data <= 17'h000b1; 
        10'b1000101001: data <= 17'h00026; 
        10'b1000101010: data <= 17'h1ffc0; 
        10'b1000101011: data <= 17'h1ffb1; 
        10'b1000101100: data <= 17'h1ffad; 
        10'b1000101101: data <= 17'h1fff3; 
        10'b1000101110: data <= 17'h1ffd8; 
        10'b1000101111: data <= 17'h0003a; 
        10'b1000110000: data <= 17'h1ffdc; 
        10'b1000110001: data <= 17'h1ffcc; 
        10'b1000110010: data <= 17'h1ffee; 
        10'b1000110011: data <= 17'h1ffc3; 
        10'b1000110100: data <= 17'h1fee4; 
        10'b1000110101: data <= 17'h1feac; 
        10'b1000110110: data <= 17'h1feda; 
        10'b1000110111: data <= 17'h1ff88; 
        10'b1000111000: data <= 17'h00050; 
        10'b1000111001: data <= 17'h00100; 
        10'b1000111010: data <= 17'h001a5; 
        10'b1000111011: data <= 17'h00119; 
        10'b1000111100: data <= 17'h00228; 
        10'b1000111101: data <= 17'h00296; 
        10'b1000111110: data <= 17'h00312; 
        10'b1000111111: data <= 17'h0029d; 
        10'b1001000000: data <= 17'h0016b; 
        10'b1001000001: data <= 17'h000e8; 
        10'b1001000010: data <= 17'h001c2; 
        10'b1001000011: data <= 17'h0013e; 
        10'b1001000100: data <= 17'h000d7; 
        10'b1001000101: data <= 17'h1ffd4; 
        10'b1001000110: data <= 17'h1ff59; 
        10'b1001000111: data <= 17'h0000b; 
        10'b1001001000: data <= 17'h1ffd8; 
        10'b1001001001: data <= 17'h1ffec; 
        10'b1001001010: data <= 17'h1ffcd; 
        10'b1001001011: data <= 17'h0000b; 
        10'b1001001100: data <= 17'h1fff9; 
        10'b1001001101: data <= 17'h00007; 
        10'b1001001110: data <= 17'h00015; 
        10'b1001001111: data <= 17'h1ffea; 
        10'b1001010000: data <= 17'h1ff94; 
        10'b1001010001: data <= 17'h1ff16; 
        10'b1001010010: data <= 17'h1fe72; 
        10'b1001010011: data <= 17'h1ff4c; 
        10'b1001010100: data <= 17'h1ff94; 
        10'b1001010101: data <= 17'h000c0; 
        10'b1001010110: data <= 17'h0015d; 
        10'b1001010111: data <= 17'h001f1; 
        10'b1001011000: data <= 17'h0027f; 
        10'b1001011001: data <= 17'h00289; 
        10'b1001011010: data <= 17'h00221; 
        10'b1001011011: data <= 17'h001d6; 
        10'b1001011100: data <= 17'h00125; 
        10'b1001011101: data <= 17'h00191; 
        10'b1001011110: data <= 17'h00176; 
        10'b1001011111: data <= 17'h000ef; 
        10'b1001100000: data <= 17'h00020; 
        10'b1001100001: data <= 17'h1ff81; 
        10'b1001100010: data <= 17'h1ff4f; 
        10'b1001100011: data <= 17'h1ff99; 
        10'b1001100100: data <= 17'h00006; 
        10'b1001100101: data <= 17'h1ffbd; 
        10'b1001100110: data <= 17'h1fff2; 
        10'b1001100111: data <= 17'h1ffdb; 
        10'b1001101000: data <= 17'h1ffdb; 
        10'b1001101001: data <= 17'h1fffa; 
        10'b1001101010: data <= 17'h00040; 
        10'b1001101011: data <= 17'h00011; 
        10'b1001101100: data <= 17'h1ffda; 
        10'b1001101101: data <= 17'h1ff34; 
        10'b1001101110: data <= 17'h1ff0e; 
        10'b1001101111: data <= 17'h1febb; 
        10'b1001110000: data <= 17'h1ff27; 
        10'b1001110001: data <= 17'h1ff9e; 
        10'b1001110010: data <= 17'h1ffaf; 
        10'b1001110011: data <= 17'h00027; 
        10'b1001110100: data <= 17'h000bb; 
        10'b1001110101: data <= 17'h00051; 
        10'b1001110110: data <= 17'h00044; 
        10'b1001110111: data <= 17'h000ca; 
        10'b1001111000: data <= 17'h00096; 
        10'b1001111001: data <= 17'h00001; 
        10'b1001111010: data <= 17'h1ffce; 
        10'b1001111011: data <= 17'h1ff1f; 
        10'b1001111100: data <= 17'h1ff27; 
        10'b1001111101: data <= 17'h1ff4c; 
        10'b1001111110: data <= 17'h1ff57; 
        10'b1001111111: data <= 17'h1fff0; 
        10'b1010000000: data <= 17'h1ffe2; 
        10'b1010000001: data <= 17'h1ffc1; 
        10'b1010000010: data <= 17'h00045; 
        10'b1010000011: data <= 17'h0001a; 
        10'b1010000100: data <= 17'h00037; 
        10'b1010000101: data <= 17'h1ffea; 
        10'b1010000110: data <= 17'h1ffe1; 
        10'b1010000111: data <= 17'h00006; 
        10'b1010001000: data <= 17'h00013; 
        10'b1010001001: data <= 17'h1ffac; 
        10'b1010001010: data <= 17'h1ff7c; 
        10'b1010001011: data <= 17'h1fedf; 
        10'b1010001100: data <= 17'h1fe92; 
        10'b1010001101: data <= 17'h1fdf2; 
        10'b1010001110: data <= 17'h1fdf4; 
        10'b1010001111: data <= 17'h1fd9e; 
        10'b1010010000: data <= 17'h1fe88; 
        10'b1010010001: data <= 17'h1fed8; 
        10'b1010010010: data <= 17'h1ff19; 
        10'b1010010011: data <= 17'h1fea8; 
        10'b1010010100: data <= 17'h1fe3c; 
        10'b1010010101: data <= 17'h1fe00; 
        10'b1010010110: data <= 17'h1fe6c; 
        10'b1010010111: data <= 17'h1ff48; 
        10'b1010011000: data <= 17'h1ff45; 
        10'b1010011001: data <= 17'h1ff5c; 
        10'b1010011010: data <= 17'h1ffc6; 
        10'b1010011011: data <= 17'h00008; 
        10'b1010011100: data <= 17'h1ffbc; 
        10'b1010011101: data <= 17'h1ffc8; 
        10'b1010011110: data <= 17'h1ffe8; 
        10'b1010011111: data <= 17'h1fff9; 
        10'b1010100000: data <= 17'h00028; 
        10'b1010100001: data <= 17'h00020; 
        10'b1010100010: data <= 17'h00016; 
        10'b1010100011: data <= 17'h1ffbf; 
        10'b1010100100: data <= 17'h1ffcc; 
        10'b1010100101: data <= 17'h1ffe8; 
        10'b1010100110: data <= 17'h1ffc2; 
        10'b1010100111: data <= 17'h1ff9b; 
        10'b1010101000: data <= 17'h1ffb0; 
        10'b1010101001: data <= 17'h1ff80; 
        10'b1010101010: data <= 17'h1ff41; 
        10'b1010101011: data <= 17'h1ff0e; 
        10'b1010101100: data <= 17'h1fee7; 
        10'b1010101101: data <= 17'h1feed; 
        10'b1010101110: data <= 17'h1febf; 
        10'b1010101111: data <= 17'h1febf; 
        10'b1010110000: data <= 17'h1feb0; 
        10'b1010110001: data <= 17'h1ff00; 
        10'b1010110010: data <= 17'h1ffa7; 
        10'b1010110011: data <= 17'h1ffad; 
        10'b1010110100: data <= 17'h1ffe3; 
        10'b1010110101: data <= 17'h1ffd2; 
        10'b1010110110: data <= 17'h00022; 
        10'b1010110111: data <= 17'h1fff1; 
        10'b1010111000: data <= 17'h1ffbd; 
        10'b1010111001: data <= 17'h1ffeb; 
        10'b1010111010: data <= 17'h1ffce; 
        10'b1010111011: data <= 17'h1ffcf; 
        10'b1010111100: data <= 17'h0003f; 
        10'b1010111101: data <= 17'h1ffc6; 
        10'b1010111110: data <= 17'h00011; 
        10'b1010111111: data <= 17'h1ffe2; 
        10'b1011000000: data <= 17'h1ffd2; 
        10'b1011000001: data <= 17'h1fff7; 
        10'b1011000010: data <= 17'h0002a; 
        10'b1011000011: data <= 17'h1fffd; 
        10'b1011000100: data <= 17'h1ffb9; 
        10'b1011000101: data <= 17'h0001a; 
        10'b1011000110: data <= 17'h1ffbb; 
        10'b1011000111: data <= 17'h1fff5; 
        10'b1011001000: data <= 17'h00003; 
        10'b1011001001: data <= 17'h1ffb7; 
        10'b1011001010: data <= 17'h1ffd8; 
        10'b1011001011: data <= 17'h1ffe7; 
        10'b1011001100: data <= 17'h1fff9; 
        10'b1011001101: data <= 17'h1ffc0; 
        10'b1011001110: data <= 17'h1ffdb; 
        10'b1011001111: data <= 17'h1ffb9; 
        10'b1011010000: data <= 17'h1ffc8; 
        10'b1011010001: data <= 17'h00009; 
        10'b1011010010: data <= 17'h1ffe5; 
        10'b1011010011: data <= 17'h00033; 
        10'b1011010100: data <= 17'h00048; 
        10'b1011010101: data <= 17'h0003f; 
        10'b1011010110: data <= 17'h00003; 
        10'b1011010111: data <= 17'h00030; 
        10'b1011011000: data <= 17'h00043; 
        10'b1011011001: data <= 17'h1fffd; 
        10'b1011011010: data <= 17'h0000c; 
        10'b1011011011: data <= 17'h1fff3; 
        10'b1011011100: data <= 17'h1ffda; 
        10'b1011011101: data <= 17'h00039; 
        10'b1011011110: data <= 17'h0002b; 
        10'b1011011111: data <= 17'h1ffdb; 
        10'b1011100000: data <= 17'h1ffea; 
        10'b1011100001: data <= 17'h00020; 
        10'b1011100010: data <= 17'h1ffe5; 
        10'b1011100011: data <= 17'h0000e; 
        10'b1011100100: data <= 17'h1ffe4; 
        10'b1011100101: data <= 17'h0002a; 
        10'b1011100110: data <= 17'h0002c; 
        10'b1011100111: data <= 17'h1ffc7; 
        10'b1011101000: data <= 17'h1ffd5; 
        10'b1011101001: data <= 17'h0003a; 
        10'b1011101010: data <= 17'h0002d; 
        10'b1011101011: data <= 17'h1ffea; 
        10'b1011101100: data <= 17'h00029; 
        10'b1011101101: data <= 17'h1fff1; 
        10'b1011101110: data <= 17'h1fff0; 
        10'b1011101111: data <= 17'h00019; 
        10'b1011110000: data <= 17'h0001d; 
        10'b1011110001: data <= 17'h1fff2; 
        10'b1011110010: data <= 17'h1ffde; 
        10'b1011110011: data <= 17'h1ffed; 
        10'b1011110100: data <= 17'h00041; 
        10'b1011110101: data <= 17'h1fffd; 
        10'b1011110110: data <= 17'h00025; 
        10'b1011110111: data <= 17'h1ffdb; 
        10'b1011111000: data <= 17'h00017; 
        10'b1011111001: data <= 17'h1fffe; 
        10'b1011111010: data <= 17'h0003d; 
        10'b1011111011: data <= 17'h00009; 
        10'b1011111100: data <= 17'h1fff8; 
        10'b1011111101: data <= 17'h1ffb8; 
        10'b1011111110: data <= 17'h1ffcf; 
        10'b1011111111: data <= 17'h00016; 
        10'b1100000000: data <= 17'h1ffbf; 
        10'b1100000001: data <= 17'h1ffca; 
        10'b1100000010: data <= 17'h1ffd7; 
        10'b1100000011: data <= 17'h1ffbe; 
        10'b1100000100: data <= 17'h1ffd3; 
        10'b1100000101: data <= 17'h1ffea; 
        10'b1100000110: data <= 17'h1ffc4; 
        10'b1100000111: data <= 17'h1ffd3; 
        10'b1100001000: data <= 17'h1ffd9; 
        10'b1100001001: data <= 17'h1ffe0; 
        10'b1100001010: data <= 17'h0003c; 
        10'b1100001011: data <= 17'h1ffc5; 
        10'b1100001100: data <= 17'h1ffda; 
        10'b1100001101: data <= 17'h1ffc7; 
        10'b1100001110: data <= 17'h1ffd8; 
        10'b1100001111: data <= 17'h0000b; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 12) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 18'h3ffd2; 
        10'b0000000001: data <= 18'h0005d; 
        10'b0000000010: data <= 18'h3ff97; 
        10'b0000000011: data <= 18'h3fff8; 
        10'b0000000100: data <= 18'h3fffd; 
        10'b0000000101: data <= 18'h3fff2; 
        10'b0000000110: data <= 18'h00031; 
        10'b0000000111: data <= 18'h00093; 
        10'b0000001000: data <= 18'h3ff9f; 
        10'b0000001001: data <= 18'h3ffc0; 
        10'b0000001010: data <= 18'h3ffc4; 
        10'b0000001011: data <= 18'h3ffa3; 
        10'b0000001100: data <= 18'h00030; 
        10'b0000001101: data <= 18'h00087; 
        10'b0000001110: data <= 18'h0004c; 
        10'b0000001111: data <= 18'h3ff85; 
        10'b0000010000: data <= 18'h3ffef; 
        10'b0000010001: data <= 18'h00093; 
        10'b0000010010: data <= 18'h00019; 
        10'b0000010011: data <= 18'h3fff3; 
        10'b0000010100: data <= 18'h3ff8f; 
        10'b0000010101: data <= 18'h3ffb4; 
        10'b0000010110: data <= 18'h00023; 
        10'b0000010111: data <= 18'h00081; 
        10'b0000011000: data <= 18'h00046; 
        10'b0000011001: data <= 18'h00055; 
        10'b0000011010: data <= 18'h3ff8d; 
        10'b0000011011: data <= 18'h3ff92; 
        10'b0000011100: data <= 18'h0005f; 
        10'b0000011101: data <= 18'h0004b; 
        10'b0000011110: data <= 18'h00060; 
        10'b0000011111: data <= 18'h3ffe8; 
        10'b0000100000: data <= 18'h3ff7f; 
        10'b0000100001: data <= 18'h3ffb3; 
        10'b0000100010: data <= 18'h00042; 
        10'b0000100011: data <= 18'h000d7; 
        10'b0000100100: data <= 18'h00092; 
        10'b0000100101: data <= 18'h0002c; 
        10'b0000100110: data <= 18'h000b0; 
        10'b0000100111: data <= 18'h000bc; 
        10'b0000101000: data <= 18'h000c8; 
        10'b0000101001: data <= 18'h000bd; 
        10'b0000101010: data <= 18'h00077; 
        10'b0000101011: data <= 18'h0007f; 
        10'b0000101100: data <= 18'h3ff78; 
        10'b0000101101: data <= 18'h00079; 
        10'b0000101110: data <= 18'h000a4; 
        10'b0000101111: data <= 18'h0005d; 
        10'b0000110000: data <= 18'h3ffe6; 
        10'b0000110001: data <= 18'h3ffad; 
        10'b0000110010: data <= 18'h000ae; 
        10'b0000110011: data <= 18'h00083; 
        10'b0000110100: data <= 18'h3ffca; 
        10'b0000110101: data <= 18'h00093; 
        10'b0000110110: data <= 18'h3ffe7; 
        10'b0000110111: data <= 18'h0006d; 
        10'b0000111000: data <= 18'h3ffaa; 
        10'b0000111001: data <= 18'h3ff99; 
        10'b0000111010: data <= 18'h3ff7f; 
        10'b0000111011: data <= 18'h3fff3; 
        10'b0000111100: data <= 18'h00049; 
        10'b0000111101: data <= 18'h0002d; 
        10'b0000111110: data <= 18'h0004b; 
        10'b0000111111: data <= 18'h000d2; 
        10'b0001000000: data <= 18'h00095; 
        10'b0001000001: data <= 18'h0013e; 
        10'b0001000010: data <= 18'h00190; 
        10'b0001000011: data <= 18'h001c4; 
        10'b0001000100: data <= 18'h001c5; 
        10'b0001000101: data <= 18'h001dc; 
        10'b0001000110: data <= 18'h000f1; 
        10'b0001000111: data <= 18'h000ab; 
        10'b0001001000: data <= 18'h0018d; 
        10'b0001001001: data <= 18'h000af; 
        10'b0001001010: data <= 18'h000ab; 
        10'b0001001011: data <= 18'h000bb; 
        10'b0001001100: data <= 18'h000b7; 
        10'b0001001101: data <= 18'h0005c; 
        10'b0001001110: data <= 18'h0007a; 
        10'b0001001111: data <= 18'h00017; 
        10'b0001010000: data <= 18'h00043; 
        10'b0001010001: data <= 18'h3ffda; 
        10'b0001010010: data <= 18'h3ff79; 
        10'b0001010011: data <= 18'h00029; 
        10'b0001010100: data <= 18'h3ff8e; 
        10'b0001010101: data <= 18'h0000d; 
        10'b0001010110: data <= 18'h0006c; 
        10'b0001010111: data <= 18'h0003e; 
        10'b0001011000: data <= 18'h0008d; 
        10'b0001011001: data <= 18'h3ff85; 
        10'b0001011010: data <= 18'h00099; 
        10'b0001011011: data <= 18'h000a8; 
        10'b0001011100: data <= 18'h000c8; 
        10'b0001011101: data <= 18'h00196; 
        10'b0001011110: data <= 18'h00167; 
        10'b0001011111: data <= 18'h001c2; 
        10'b0001100000: data <= 18'h001b7; 
        10'b0001100001: data <= 18'h001a7; 
        10'b0001100010: data <= 18'h0026e; 
        10'b0001100011: data <= 18'h0024a; 
        10'b0001100100: data <= 18'h0016d; 
        10'b0001100101: data <= 18'h001cc; 
        10'b0001100110: data <= 18'h002e4; 
        10'b0001100111: data <= 18'h002e1; 
        10'b0001101000: data <= 18'h00313; 
        10'b0001101001: data <= 18'h002b9; 
        10'b0001101010: data <= 18'h002c2; 
        10'b0001101011: data <= 18'h0019a; 
        10'b0001101100: data <= 18'h0016c; 
        10'b0001101101: data <= 18'h00059; 
        10'b0001101110: data <= 18'h3ffc2; 
        10'b0001101111: data <= 18'h00050; 
        10'b0001110000: data <= 18'h00015; 
        10'b0001110001: data <= 18'h3ffe5; 
        10'b0001110010: data <= 18'h3fff7; 
        10'b0001110011: data <= 18'h0007d; 
        10'b0001110100: data <= 18'h0006c; 
        10'b0001110101: data <= 18'h00027; 
        10'b0001110110: data <= 18'h00028; 
        10'b0001110111: data <= 18'h000fb; 
        10'b0001111000: data <= 18'h3ffe4; 
        10'b0001111001: data <= 18'h3ffcc; 
        10'b0001111010: data <= 18'h000f3; 
        10'b0001111011: data <= 18'h0005b; 
        10'b0001111100: data <= 18'h00071; 
        10'b0001111101: data <= 18'h00029; 
        10'b0001111110: data <= 18'h00060; 
        10'b0001111111: data <= 18'h00090; 
        10'b0010000000: data <= 18'h001ed; 
        10'b0010000001: data <= 18'h001e8; 
        10'b0010000010: data <= 18'h002fc; 
        10'b0010000011: data <= 18'h00309; 
        10'b0010000100: data <= 18'h003d5; 
        10'b0010000101: data <= 18'h00440; 
        10'b0010000110: data <= 18'h003a8; 
        10'b0010000111: data <= 18'h00275; 
        10'b0010001000: data <= 18'h00059; 
        10'b0010001001: data <= 18'h000a7; 
        10'b0010001010: data <= 18'h00017; 
        10'b0010001011: data <= 18'h00000; 
        10'b0010001100: data <= 18'h00019; 
        10'b0010001101: data <= 18'h0004c; 
        10'b0010001110: data <= 18'h0002b; 
        10'b0010001111: data <= 18'h3ffc6; 
        10'b0010010000: data <= 18'h3ff98; 
        10'b0010010001: data <= 18'h3fff5; 
        10'b0010010010: data <= 18'h3ffa9; 
        10'b0010010011: data <= 18'h3ff54; 
        10'b0010010100: data <= 18'h00081; 
        10'b0010010101: data <= 18'h3ff5a; 
        10'b0010010110: data <= 18'h0003c; 
        10'b0010010111: data <= 18'h3fdc5; 
        10'b0010011000: data <= 18'h3fed2; 
        10'b0010011001: data <= 18'h3ff2f; 
        10'b0010011010: data <= 18'h3ffb3; 
        10'b0010011011: data <= 18'h3fef2; 
        10'b0010011100: data <= 18'h3fef2; 
        10'b0010011101: data <= 18'h00034; 
        10'b0010011110: data <= 18'h0016f; 
        10'b0010011111: data <= 18'h002af; 
        10'b0010100000: data <= 18'h00255; 
        10'b0010100001: data <= 18'h00215; 
        10'b0010100010: data <= 18'h001a5; 
        10'b0010100011: data <= 18'h00121; 
        10'b0010100100: data <= 18'h3ffdf; 
        10'b0010100101: data <= 18'h0000e; 
        10'b0010100110: data <= 18'h3ff6f; 
        10'b0010100111: data <= 18'h00089; 
        10'b0010101000: data <= 18'h3ffed; 
        10'b0010101001: data <= 18'h0007b; 
        10'b0010101010: data <= 18'h00073; 
        10'b0010101011: data <= 18'h3ff6c; 
        10'b0010101100: data <= 18'h00035; 
        10'b0010101101: data <= 18'h3ffe9; 
        10'b0010101110: data <= 18'h00030; 
        10'b0010101111: data <= 18'h00004; 
        10'b0010110000: data <= 18'h3ff2c; 
        10'b0010110001: data <= 18'h3fefe; 
        10'b0010110010: data <= 18'h3fd6f; 
        10'b0010110011: data <= 18'h3fca4; 
        10'b0010110100: data <= 18'h3fe0d; 
        10'b0010110101: data <= 18'h3fc2c; 
        10'b0010110110: data <= 18'h3fe50; 
        10'b0010110111: data <= 18'h3fec3; 
        10'b0010111000: data <= 18'h3fe3c; 
        10'b0010111001: data <= 18'h3fe70; 
        10'b0010111010: data <= 18'h3ff91; 
        10'b0010111011: data <= 18'h3fef4; 
        10'b0010111100: data <= 18'h3fe4e; 
        10'b0010111101: data <= 18'h3fe62; 
        10'b0010111110: data <= 18'h3fd7c; 
        10'b0010111111: data <= 18'h3fe5c; 
        10'b0011000000: data <= 18'h3fea4; 
        10'b0011000001: data <= 18'h3fe91; 
        10'b0011000010: data <= 18'h3ffc9; 
        10'b0011000011: data <= 18'h00078; 
        10'b0011000100: data <= 18'h00030; 
        10'b0011000101: data <= 18'h00047; 
        10'b0011000110: data <= 18'h00004; 
        10'b0011000111: data <= 18'h3ffe8; 
        10'b0011001000: data <= 18'h00008; 
        10'b0011001001: data <= 18'h3ff81; 
        10'b0011001010: data <= 18'h3fefe; 
        10'b0011001011: data <= 18'h3ffd6; 
        10'b0011001100: data <= 18'h3fe92; 
        10'b0011001101: data <= 18'h3fe39; 
        10'b0011001110: data <= 18'h3fd6a; 
        10'b0011001111: data <= 18'h3fdf7; 
        10'b0011010000: data <= 18'h3fc58; 
        10'b0011010001: data <= 18'h3fbe7; 
        10'b0011010010: data <= 18'h3fdda; 
        10'b0011010011: data <= 18'h3fdf6; 
        10'b0011010100: data <= 18'h3fccf; 
        10'b0011010101: data <= 18'h3fcfa; 
        10'b0011010110: data <= 18'h3fc40; 
        10'b0011010111: data <= 18'h3faea; 
        10'b0011011000: data <= 18'h3facf; 
        10'b0011011001: data <= 18'h3fba9; 
        10'b0011011010: data <= 18'h3fb76; 
        10'b0011011011: data <= 18'h3fc6a; 
        10'b0011011100: data <= 18'h3fea1; 
        10'b0011011101: data <= 18'h3fec3; 
        10'b0011011110: data <= 18'h3ff83; 
        10'b0011011111: data <= 18'h3ffa0; 
        10'b0011100000: data <= 18'h3ffd2; 
        10'b0011100001: data <= 18'h3ffd9; 
        10'b0011100010: data <= 18'h0008c; 
        10'b0011100011: data <= 18'h3ff4c; 
        10'b0011100100: data <= 18'h3ff6b; 
        10'b0011100101: data <= 18'h3ff39; 
        10'b0011100110: data <= 18'h3fe0d; 
        10'b0011100111: data <= 18'h3ff92; 
        10'b0011101000: data <= 18'h3ff48; 
        10'b0011101001: data <= 18'h3fdf6; 
        10'b0011101010: data <= 18'h3fd9f; 
        10'b0011101011: data <= 18'h3fd45; 
        10'b0011101100: data <= 18'h3fcb7; 
        10'b0011101101: data <= 18'h3fc31; 
        10'b0011101110: data <= 18'h3fc4a; 
        10'b0011101111: data <= 18'h3fc09; 
        10'b0011110000: data <= 18'h3fb4d; 
        10'b0011110001: data <= 18'h3fa96; 
        10'b0011110010: data <= 18'h3f859; 
        10'b0011110011: data <= 18'h3f8e0; 
        10'b0011110100: data <= 18'h3f9a1; 
        10'b0011110101: data <= 18'h3f9b1; 
        10'b0011110110: data <= 18'h3fb98; 
        10'b0011110111: data <= 18'h3fc1e; 
        10'b0011111000: data <= 18'h3fd94; 
        10'b0011111001: data <= 18'h3fe79; 
        10'b0011111010: data <= 18'h3fee7; 
        10'b0011111011: data <= 18'h0002a; 
        10'b0011111100: data <= 18'h3ffec; 
        10'b0011111101: data <= 18'h3ff93; 
        10'b0011111110: data <= 18'h3ffc1; 
        10'b0011111111: data <= 18'h3ff84; 
        10'b0100000000: data <= 18'h00004; 
        10'b0100000001: data <= 18'h3ff8e; 
        10'b0100000010: data <= 18'h3ff52; 
        10'b0100000011: data <= 18'h3ff9b; 
        10'b0100000100: data <= 18'h00077; 
        10'b0100000101: data <= 18'h3fec5; 
        10'b0100000110: data <= 18'h3fdac; 
        10'b0100000111: data <= 18'h3fe37; 
        10'b0100001000: data <= 18'h3feda; 
        10'b0100001001: data <= 18'h3fdd5; 
        10'b0100001010: data <= 18'h3fe04; 
        10'b0100001011: data <= 18'h3fba8; 
        10'b0100001100: data <= 18'h3faf0; 
        10'b0100001101: data <= 18'h3f8ab; 
        10'b0100001110: data <= 18'h3f82e; 
        10'b0100001111: data <= 18'h3f99d; 
        10'b0100010000: data <= 18'h3fac3; 
        10'b0100010001: data <= 18'h3fbd5; 
        10'b0100010010: data <= 18'h3fb2c; 
        10'b0100010011: data <= 18'h3fce6; 
        10'b0100010100: data <= 18'h3fda2; 
        10'b0100010101: data <= 18'h3fe3e; 
        10'b0100010110: data <= 18'h3ff47; 
        10'b0100010111: data <= 18'h00061; 
        10'b0100011000: data <= 18'h3ffa2; 
        10'b0100011001: data <= 18'h0007b; 
        10'b0100011010: data <= 18'h00053; 
        10'b0100011011: data <= 18'h3ff70; 
        10'b0100011100: data <= 18'h3ff2e; 
        10'b0100011101: data <= 18'h00035; 
        10'b0100011110: data <= 18'h000ad; 
        10'b0100011111: data <= 18'h000a6; 
        10'b0100100000: data <= 18'h00260; 
        10'b0100100001: data <= 18'h3fff3; 
        10'b0100100010: data <= 18'h00079; 
        10'b0100100011: data <= 18'h00032; 
        10'b0100100100: data <= 18'h3fe90; 
        10'b0100100101: data <= 18'h3ff06; 
        10'b0100100110: data <= 18'h3fddb; 
        10'b0100100111: data <= 18'h3fb81; 
        10'b0100101000: data <= 18'h3fb6e; 
        10'b0100101001: data <= 18'h3faa4; 
        10'b0100101010: data <= 18'h3fa6b; 
        10'b0100101011: data <= 18'h3fb8b; 
        10'b0100101100: data <= 18'h3fcf9; 
        10'b0100101101: data <= 18'h3fdd5; 
        10'b0100101110: data <= 18'h3fd26; 
        10'b0100101111: data <= 18'h3ffb4; 
        10'b0100110000: data <= 18'h3fe25; 
        10'b0100110001: data <= 18'h3feb6; 
        10'b0100110010: data <= 18'h3ff9e; 
        10'b0100110011: data <= 18'h3ffd1; 
        10'b0100110100: data <= 18'h3ffb4; 
        10'b0100110101: data <= 18'h00032; 
        10'b0100110110: data <= 18'h3ffac; 
        10'b0100110111: data <= 18'h3fff4; 
        10'b0100111000: data <= 18'h3ffad; 
        10'b0100111001: data <= 18'h00016; 
        10'b0100111010: data <= 18'h3ffd3; 
        10'b0100111011: data <= 18'h001fd; 
        10'b0100111100: data <= 18'h0016c; 
        10'b0100111101: data <= 18'h000af; 
        10'b0100111110: data <= 18'h000dc; 
        10'b0100111111: data <= 18'h0009c; 
        10'b0101000000: data <= 18'h0009c; 
        10'b0101000001: data <= 18'h00019; 
        10'b0101000010: data <= 18'h3fef7; 
        10'b0101000011: data <= 18'h3fc6f; 
        10'b0101000100: data <= 18'h3fca8; 
        10'b0101000101: data <= 18'h3fd27; 
        10'b0101000110: data <= 18'h3fd24; 
        10'b0101000111: data <= 18'h3fdc6; 
        10'b0101001000: data <= 18'h3fef6; 
        10'b0101001001: data <= 18'h00067; 
        10'b0101001010: data <= 18'h0015d; 
        10'b0101001011: data <= 18'h0021f; 
        10'b0101001100: data <= 18'h3ffff; 
        10'b0101001101: data <= 18'h3fedf; 
        10'b0101001110: data <= 18'h3ff87; 
        10'b0101001111: data <= 18'h3ffd4; 
        10'b0101010000: data <= 18'h3ffb3; 
        10'b0101010001: data <= 18'h3ffd7; 
        10'b0101010010: data <= 18'h3ff83; 
        10'b0101010011: data <= 18'h3ffc4; 
        10'b0101010100: data <= 18'h00049; 
        10'b0101010101: data <= 18'h000ee; 
        10'b0101010110: data <= 18'h0016c; 
        10'b0101010111: data <= 18'h001dd; 
        10'b0101011000: data <= 18'h000dd; 
        10'b0101011001: data <= 18'h00136; 
        10'b0101011010: data <= 18'h000db; 
        10'b0101011011: data <= 18'h0023f; 
        10'b0101011100: data <= 18'h00229; 
        10'b0101011101: data <= 18'h0018c; 
        10'b0101011110: data <= 18'h3fead; 
        10'b0101011111: data <= 18'h3fd9c; 
        10'b0101100000: data <= 18'h3ffe6; 
        10'b0101100001: data <= 18'h3ffc7; 
        10'b0101100010: data <= 18'h3fda8; 
        10'b0101100011: data <= 18'h3fdc1; 
        10'b0101100100: data <= 18'h3ffb9; 
        10'b0101100101: data <= 18'h00144; 
        10'b0101100110: data <= 18'h00310; 
        10'b0101100111: data <= 18'h0056f; 
        10'b0101101000: data <= 18'h002ec; 
        10'b0101101001: data <= 18'h3ff2b; 
        10'b0101101010: data <= 18'h3ff0b; 
        10'b0101101011: data <= 18'h3ffb6; 
        10'b0101101100: data <= 18'h3ffb7; 
        10'b0101101101: data <= 18'h00081; 
        10'b0101101110: data <= 18'h00063; 
        10'b0101101111: data <= 18'h3ff73; 
        10'b0101110000: data <= 18'h3ff40; 
        10'b0101110001: data <= 18'h0004d; 
        10'b0101110010: data <= 18'h0025c; 
        10'b0101110011: data <= 18'h00145; 
        10'b0101110100: data <= 18'h00117; 
        10'b0101110101: data <= 18'h0008a; 
        10'b0101110110: data <= 18'h0024a; 
        10'b0101110111: data <= 18'h001e9; 
        10'b0101111000: data <= 18'h001c1; 
        10'b0101111001: data <= 18'h0004f; 
        10'b0101111010: data <= 18'h3ffad; 
        10'b0101111011: data <= 18'h3fff2; 
        10'b0101111100: data <= 18'h0002d; 
        10'b0101111101: data <= 18'h3ff7c; 
        10'b0101111110: data <= 18'h3fdf6; 
        10'b0101111111: data <= 18'h3ffbb; 
        10'b0110000000: data <= 18'h3ff05; 
        10'b0110000001: data <= 18'h001a1; 
        10'b0110000010: data <= 18'h0043d; 
        10'b0110000011: data <= 18'h006b8; 
        10'b0110000100: data <= 18'h003a1; 
        10'b0110000101: data <= 18'h3ffb6; 
        10'b0110000110: data <= 18'h00003; 
        10'b0110000111: data <= 18'h00054; 
        10'b0110001000: data <= 18'h3ffc2; 
        10'b0110001001: data <= 18'h0000e; 
        10'b0110001010: data <= 18'h00061; 
        10'b0110001011: data <= 18'h00005; 
        10'b0110001100: data <= 18'h3ff35; 
        10'b0110001101: data <= 18'h000d8; 
        10'b0110001110: data <= 18'h0022a; 
        10'b0110001111: data <= 18'h001dd; 
        10'b0110010000: data <= 18'h00291; 
        10'b0110010001: data <= 18'h00267; 
        10'b0110010010: data <= 18'h0029a; 
        10'b0110010011: data <= 18'h002d1; 
        10'b0110010100: data <= 18'h000f3; 
        10'b0110010101: data <= 18'h3fea0; 
        10'b0110010110: data <= 18'h00017; 
        10'b0110010111: data <= 18'h00126; 
        10'b0110011000: data <= 18'h0008b; 
        10'b0110011001: data <= 18'h3ff1b; 
        10'b0110011010: data <= 18'h3ff22; 
        10'b0110011011: data <= 18'h3ffe0; 
        10'b0110011100: data <= 18'h001d7; 
        10'b0110011101: data <= 18'h001d2; 
        10'b0110011110: data <= 18'h004cd; 
        10'b0110011111: data <= 18'h00596; 
        10'b0110100000: data <= 18'h003aa; 
        10'b0110100001: data <= 18'h3fff3; 
        10'b0110100010: data <= 18'h3fef4; 
        10'b0110100011: data <= 18'h3ff7c; 
        10'b0110100100: data <= 18'h00064; 
        10'b0110100101: data <= 18'h3ffcd; 
        10'b0110100110: data <= 18'h00014; 
        10'b0110100111: data <= 18'h3ff91; 
        10'b0110101000: data <= 18'h3fe7c; 
        10'b0110101001: data <= 18'h3ffcf; 
        10'b0110101010: data <= 18'h00241; 
        10'b0110101011: data <= 18'h002ff; 
        10'b0110101100: data <= 18'h001ee; 
        10'b0110101101: data <= 18'h00307; 
        10'b0110101110: data <= 18'h003d1; 
        10'b0110101111: data <= 18'h004a9; 
        10'b0110110000: data <= 18'h00138; 
        10'b0110110001: data <= 18'h3ffaa; 
        10'b0110110010: data <= 18'h001cc; 
        10'b0110110011: data <= 18'h001a7; 
        10'b0110110100: data <= 18'h00042; 
        10'b0110110101: data <= 18'h3ff27; 
        10'b0110110110: data <= 18'h0002c; 
        10'b0110110111: data <= 18'h000ed; 
        10'b0110111000: data <= 18'h00227; 
        10'b0110111001: data <= 18'h002f4; 
        10'b0110111010: data <= 18'h002b7; 
        10'b0110111011: data <= 18'h0035d; 
        10'b0110111100: data <= 18'h001cb; 
        10'b0110111101: data <= 18'h3ff14; 
        10'b0110111110: data <= 18'h3ff6d; 
        10'b0110111111: data <= 18'h3ff6a; 
        10'b0111000000: data <= 18'h0001b; 
        10'b0111000001: data <= 18'h3ff92; 
        10'b0111000010: data <= 18'h3ff8e; 
        10'b0111000011: data <= 18'h3ff82; 
        10'b0111000100: data <= 18'h3fdff; 
        10'b0111000101: data <= 18'h3feea; 
        10'b0111000110: data <= 18'h00357; 
        10'b0111000111: data <= 18'h0036a; 
        10'b0111001000: data <= 18'h00242; 
        10'b0111001001: data <= 18'h0037c; 
        10'b0111001010: data <= 18'h005e9; 
        10'b0111001011: data <= 18'h005dc; 
        10'b0111001100: data <= 18'h001ca; 
        10'b0111001101: data <= 18'h00110; 
        10'b0111001110: data <= 18'h0028c; 
        10'b0111001111: data <= 18'h00158; 
        10'b0111010000: data <= 18'h3ff4c; 
        10'b0111010001: data <= 18'h3fe9b; 
        10'b0111010010: data <= 18'h0007b; 
        10'b0111010011: data <= 18'h0017d; 
        10'b0111010100: data <= 18'h000b1; 
        10'b0111010101: data <= 18'h00005; 
        10'b0111010110: data <= 18'h00164; 
        10'b0111010111: data <= 18'h000d5; 
        10'b0111011000: data <= 18'h3ff98; 
        10'b0111011001: data <= 18'h3feeb; 
        10'b0111011010: data <= 18'h3ff56; 
        10'b0111011011: data <= 18'h3ffe9; 
        10'b0111011100: data <= 18'h00019; 
        10'b0111011101: data <= 18'h00054; 
        10'b0111011110: data <= 18'h00074; 
        10'b0111011111: data <= 18'h3ffec; 
        10'b0111100000: data <= 18'h3fd24; 
        10'b0111100001: data <= 18'h3fe81; 
        10'b0111100010: data <= 18'h00166; 
        10'b0111100011: data <= 18'h002a7; 
        10'b0111100100: data <= 18'h00305; 
        10'b0111100101: data <= 18'h003cf; 
        10'b0111100110: data <= 18'h00693; 
        10'b0111100111: data <= 18'h006ae; 
        10'b0111101000: data <= 18'h00374; 
        10'b0111101001: data <= 18'h001f2; 
        10'b0111101010: data <= 18'h001f8; 
        10'b0111101011: data <= 18'h0013e; 
        10'b0111101100: data <= 18'h00000; 
        10'b0111101101: data <= 18'h0005c; 
        10'b0111101110: data <= 18'h002bd; 
        10'b0111101111: data <= 18'h000f2; 
        10'b0111110000: data <= 18'h00064; 
        10'b0111110001: data <= 18'h3ff4d; 
        10'b0111110010: data <= 18'h000a0; 
        10'b0111110011: data <= 18'h3ffde; 
        10'b0111110100: data <= 18'h3ff39; 
        10'b0111110101: data <= 18'h3fe7c; 
        10'b0111110110: data <= 18'h3ffc8; 
        10'b0111110111: data <= 18'h0003f; 
        10'b0111111000: data <= 18'h3ffc7; 
        10'b0111111001: data <= 18'h3ffb1; 
        10'b0111111010: data <= 18'h3fffe; 
        10'b0111111011: data <= 18'h3ff2b; 
        10'b0111111100: data <= 18'h3fd52; 
        10'b0111111101: data <= 18'h3fd62; 
        10'b0111111110: data <= 18'h3febc; 
        10'b0111111111: data <= 18'h001d3; 
        10'b1000000000: data <= 18'h002ed; 
        10'b1000000001: data <= 18'h002a9; 
        10'b1000000010: data <= 18'h0049a; 
        10'b1000000011: data <= 18'h005ae; 
        10'b1000000100: data <= 18'h006b1; 
        10'b1000000101: data <= 18'h0031c; 
        10'b1000000110: data <= 18'h000d7; 
        10'b1000000111: data <= 18'h001bb; 
        10'b1000001000: data <= 18'h002fc; 
        10'b1000001001: data <= 18'h001f0; 
        10'b1000001010: data <= 18'h00269; 
        10'b1000001011: data <= 18'h00145; 
        10'b1000001100: data <= 18'h0002a; 
        10'b1000001101: data <= 18'h0006c; 
        10'b1000001110: data <= 18'h00078; 
        10'b1000001111: data <= 18'h3ffbc; 
        10'b1000010000: data <= 18'h3ff0c; 
        10'b1000010001: data <= 18'h3ff4c; 
        10'b1000010010: data <= 18'h3ff74; 
        10'b1000010011: data <= 18'h3ff6b; 
        10'b1000010100: data <= 18'h00025; 
        10'b1000010101: data <= 18'h3ff98; 
        10'b1000010110: data <= 18'h00041; 
        10'b1000010111: data <= 18'h3fef1; 
        10'b1000011000: data <= 18'h3fe44; 
        10'b1000011001: data <= 18'h3fd37; 
        10'b1000011010: data <= 18'h3fdd6; 
        10'b1000011011: data <= 18'h00027; 
        10'b1000011100: data <= 18'h001e6; 
        10'b1000011101: data <= 18'h002fb; 
        10'b1000011110: data <= 18'h003f9; 
        10'b1000011111: data <= 18'h00654; 
        10'b1000100000: data <= 18'h0071f; 
        10'b1000100001: data <= 18'h003ac; 
        10'b1000100010: data <= 18'h00348; 
        10'b1000100011: data <= 18'h0036e; 
        10'b1000100100: data <= 18'h00271; 
        10'b1000100101: data <= 18'h00202; 
        10'b1000100110: data <= 18'h00321; 
        10'b1000100111: data <= 18'h00222; 
        10'b1000101000: data <= 18'h00161; 
        10'b1000101001: data <= 18'h0004c; 
        10'b1000101010: data <= 18'h3ff80; 
        10'b1000101011: data <= 18'h3ff62; 
        10'b1000101100: data <= 18'h3ff5b; 
        10'b1000101101: data <= 18'h3ffe5; 
        10'b1000101110: data <= 18'h3ffb1; 
        10'b1000101111: data <= 18'h00075; 
        10'b1000110000: data <= 18'h3ffb8; 
        10'b1000110001: data <= 18'h3ff98; 
        10'b1000110010: data <= 18'h3ffdb; 
        10'b1000110011: data <= 18'h3ff85; 
        10'b1000110100: data <= 18'h3fdc7; 
        10'b1000110101: data <= 18'h3fd58; 
        10'b1000110110: data <= 18'h3fdb3; 
        10'b1000110111: data <= 18'h3ff0f; 
        10'b1000111000: data <= 18'h000a1; 
        10'b1000111001: data <= 18'h001ff; 
        10'b1000111010: data <= 18'h0034a; 
        10'b1000111011: data <= 18'h00231; 
        10'b1000111100: data <= 18'h00451; 
        10'b1000111101: data <= 18'h0052c; 
        10'b1000111110: data <= 18'h00624; 
        10'b1000111111: data <= 18'h0053a; 
        10'b1001000000: data <= 18'h002d5; 
        10'b1001000001: data <= 18'h001d0; 
        10'b1001000010: data <= 18'h00385; 
        10'b1001000011: data <= 18'h0027b; 
        10'b1001000100: data <= 18'h001af; 
        10'b1001000101: data <= 18'h3ffa8; 
        10'b1001000110: data <= 18'h3feb2; 
        10'b1001000111: data <= 18'h00016; 
        10'b1001001000: data <= 18'h3ffaf; 
        10'b1001001001: data <= 18'h3ffd8; 
        10'b1001001010: data <= 18'h3ff9b; 
        10'b1001001011: data <= 18'h00015; 
        10'b1001001100: data <= 18'h3fff3; 
        10'b1001001101: data <= 18'h0000d; 
        10'b1001001110: data <= 18'h0002b; 
        10'b1001001111: data <= 18'h3ffd5; 
        10'b1001010000: data <= 18'h3ff28; 
        10'b1001010001: data <= 18'h3fe2c; 
        10'b1001010010: data <= 18'h3fce5; 
        10'b1001010011: data <= 18'h3fe98; 
        10'b1001010100: data <= 18'h3ff28; 
        10'b1001010101: data <= 18'h00181; 
        10'b1001010110: data <= 18'h002bb; 
        10'b1001010111: data <= 18'h003e2; 
        10'b1001011000: data <= 18'h004fe; 
        10'b1001011001: data <= 18'h00512; 
        10'b1001011010: data <= 18'h00441; 
        10'b1001011011: data <= 18'h003ab; 
        10'b1001011100: data <= 18'h0024a; 
        10'b1001011101: data <= 18'h00321; 
        10'b1001011110: data <= 18'h002eb; 
        10'b1001011111: data <= 18'h001de; 
        10'b1001100000: data <= 18'h00040; 
        10'b1001100001: data <= 18'h3ff03; 
        10'b1001100010: data <= 18'h3fe9e; 
        10'b1001100011: data <= 18'h3ff32; 
        10'b1001100100: data <= 18'h0000c; 
        10'b1001100101: data <= 18'h3ff7b; 
        10'b1001100110: data <= 18'h3ffe3; 
        10'b1001100111: data <= 18'h3ffb6; 
        10'b1001101000: data <= 18'h3ffb5; 
        10'b1001101001: data <= 18'h3fff3; 
        10'b1001101010: data <= 18'h0007f; 
        10'b1001101011: data <= 18'h00023; 
        10'b1001101100: data <= 18'h3ffb5; 
        10'b1001101101: data <= 18'h3fe68; 
        10'b1001101110: data <= 18'h3fe1c; 
        10'b1001101111: data <= 18'h3fd76; 
        10'b1001110000: data <= 18'h3fe4f; 
        10'b1001110001: data <= 18'h3ff3b; 
        10'b1001110010: data <= 18'h3ff5e; 
        10'b1001110011: data <= 18'h0004e; 
        10'b1001110100: data <= 18'h00176; 
        10'b1001110101: data <= 18'h000a2; 
        10'b1001110110: data <= 18'h00088; 
        10'b1001110111: data <= 18'h00193; 
        10'b1001111000: data <= 18'h0012c; 
        10'b1001111001: data <= 18'h00003; 
        10'b1001111010: data <= 18'h3ff9c; 
        10'b1001111011: data <= 18'h3fe3d; 
        10'b1001111100: data <= 18'h3fe4e; 
        10'b1001111101: data <= 18'h3fe97; 
        10'b1001111110: data <= 18'h3feaf; 
        10'b1001111111: data <= 18'h3ffdf; 
        10'b1010000000: data <= 18'h3ffc5; 
        10'b1010000001: data <= 18'h3ff82; 
        10'b1010000010: data <= 18'h0008a; 
        10'b1010000011: data <= 18'h00035; 
        10'b1010000100: data <= 18'h0006e; 
        10'b1010000101: data <= 18'h3ffd4; 
        10'b1010000110: data <= 18'h3ffc2; 
        10'b1010000111: data <= 18'h0000d; 
        10'b1010001000: data <= 18'h00027; 
        10'b1010001001: data <= 18'h3ff57; 
        10'b1010001010: data <= 18'h3fef8; 
        10'b1010001011: data <= 18'h3fdbd; 
        10'b1010001100: data <= 18'h3fd24; 
        10'b1010001101: data <= 18'h3fbe3; 
        10'b1010001110: data <= 18'h3fbe8; 
        10'b1010001111: data <= 18'h3fb3b; 
        10'b1010010000: data <= 18'h3fd10; 
        10'b1010010001: data <= 18'h3fdaf; 
        10'b1010010010: data <= 18'h3fe32; 
        10'b1010010011: data <= 18'h3fd51; 
        10'b1010010100: data <= 18'h3fc79; 
        10'b1010010101: data <= 18'h3fc00; 
        10'b1010010110: data <= 18'h3fcd9; 
        10'b1010010111: data <= 18'h3fe90; 
        10'b1010011000: data <= 18'h3fe89; 
        10'b1010011001: data <= 18'h3feb8; 
        10'b1010011010: data <= 18'h3ff8b; 
        10'b1010011011: data <= 18'h00010; 
        10'b1010011100: data <= 18'h3ff77; 
        10'b1010011101: data <= 18'h3ff8f; 
        10'b1010011110: data <= 18'h3ffd0; 
        10'b1010011111: data <= 18'h3fff2; 
        10'b1010100000: data <= 18'h0004f; 
        10'b1010100001: data <= 18'h00040; 
        10'b1010100010: data <= 18'h0002b; 
        10'b1010100011: data <= 18'h3ff7e; 
        10'b1010100100: data <= 18'h3ff99; 
        10'b1010100101: data <= 18'h3ffcf; 
        10'b1010100110: data <= 18'h3ff83; 
        10'b1010100111: data <= 18'h3ff36; 
        10'b1010101000: data <= 18'h3ff60; 
        10'b1010101001: data <= 18'h3ff01; 
        10'b1010101010: data <= 18'h3fe82; 
        10'b1010101011: data <= 18'h3fe1c; 
        10'b1010101100: data <= 18'h3fdce; 
        10'b1010101101: data <= 18'h3fdda; 
        10'b1010101110: data <= 18'h3fd7d; 
        10'b1010101111: data <= 18'h3fd7e; 
        10'b1010110000: data <= 18'h3fd61; 
        10'b1010110001: data <= 18'h3fe00; 
        10'b1010110010: data <= 18'h3ff4e; 
        10'b1010110011: data <= 18'h3ff5b; 
        10'b1010110100: data <= 18'h3ffc6; 
        10'b1010110101: data <= 18'h3ffa5; 
        10'b1010110110: data <= 18'h00044; 
        10'b1010110111: data <= 18'h3ffe2; 
        10'b1010111000: data <= 18'h3ff7a; 
        10'b1010111001: data <= 18'h3ffd6; 
        10'b1010111010: data <= 18'h3ff9c; 
        10'b1010111011: data <= 18'h3ff9f; 
        10'b1010111100: data <= 18'h0007d; 
        10'b1010111101: data <= 18'h3ff8c; 
        10'b1010111110: data <= 18'h00022; 
        10'b1010111111: data <= 18'h3ffc5; 
        10'b1011000000: data <= 18'h3ffa5; 
        10'b1011000001: data <= 18'h3ffef; 
        10'b1011000010: data <= 18'h00053; 
        10'b1011000011: data <= 18'h3fff9; 
        10'b1011000100: data <= 18'h3ff72; 
        10'b1011000101: data <= 18'h00033; 
        10'b1011000110: data <= 18'h3ff75; 
        10'b1011000111: data <= 18'h3ffeb; 
        10'b1011001000: data <= 18'h00007; 
        10'b1011001001: data <= 18'h3ff6d; 
        10'b1011001010: data <= 18'h3ffaf; 
        10'b1011001011: data <= 18'h3ffcf; 
        10'b1011001100: data <= 18'h3fff3; 
        10'b1011001101: data <= 18'h3ff80; 
        10'b1011001110: data <= 18'h3ffb5; 
        10'b1011001111: data <= 18'h3ff73; 
        10'b1011010000: data <= 18'h3ff91; 
        10'b1011010001: data <= 18'h00012; 
        10'b1011010010: data <= 18'h3ffcb; 
        10'b1011010011: data <= 18'h00066; 
        10'b1011010100: data <= 18'h00090; 
        10'b1011010101: data <= 18'h0007f; 
        10'b1011010110: data <= 18'h00006; 
        10'b1011010111: data <= 18'h0005f; 
        10'b1011011000: data <= 18'h00087; 
        10'b1011011001: data <= 18'h3fffa; 
        10'b1011011010: data <= 18'h00019; 
        10'b1011011011: data <= 18'h3ffe6; 
        10'b1011011100: data <= 18'h3ffb4; 
        10'b1011011101: data <= 18'h00072; 
        10'b1011011110: data <= 18'h00056; 
        10'b1011011111: data <= 18'h3ffb6; 
        10'b1011100000: data <= 18'h3ffd4; 
        10'b1011100001: data <= 18'h00040; 
        10'b1011100010: data <= 18'h3ffcb; 
        10'b1011100011: data <= 18'h0001c; 
        10'b1011100100: data <= 18'h3ffc8; 
        10'b1011100101: data <= 18'h00054; 
        10'b1011100110: data <= 18'h00058; 
        10'b1011100111: data <= 18'h3ff8e; 
        10'b1011101000: data <= 18'h3ffa9; 
        10'b1011101001: data <= 18'h00073; 
        10'b1011101010: data <= 18'h0005a; 
        10'b1011101011: data <= 18'h3ffd4; 
        10'b1011101100: data <= 18'h00051; 
        10'b1011101101: data <= 18'h3ffe1; 
        10'b1011101110: data <= 18'h3ffe0; 
        10'b1011101111: data <= 18'h00032; 
        10'b1011110000: data <= 18'h0003a; 
        10'b1011110001: data <= 18'h3ffe4; 
        10'b1011110010: data <= 18'h3ffbc; 
        10'b1011110011: data <= 18'h3ffd9; 
        10'b1011110100: data <= 18'h00082; 
        10'b1011110101: data <= 18'h3fffa; 
        10'b1011110110: data <= 18'h0004a; 
        10'b1011110111: data <= 18'h3ffb5; 
        10'b1011111000: data <= 18'h0002e; 
        10'b1011111001: data <= 18'h3fffc; 
        10'b1011111010: data <= 18'h0007a; 
        10'b1011111011: data <= 18'h00011; 
        10'b1011111100: data <= 18'h3fff0; 
        10'b1011111101: data <= 18'h3ff70; 
        10'b1011111110: data <= 18'h3ff9e; 
        10'b1011111111: data <= 18'h0002c; 
        10'b1100000000: data <= 18'h3ff7e; 
        10'b1100000001: data <= 18'h3ff93; 
        10'b1100000010: data <= 18'h3ffad; 
        10'b1100000011: data <= 18'h3ff7b; 
        10'b1100000100: data <= 18'h3ffa6; 
        10'b1100000101: data <= 18'h3ffd3; 
        10'b1100000110: data <= 18'h3ff89; 
        10'b1100000111: data <= 18'h3ffa6; 
        10'b1100001000: data <= 18'h3ffb2; 
        10'b1100001001: data <= 18'h3ffc0; 
        10'b1100001010: data <= 18'h00079; 
        10'b1100001011: data <= 18'h3ff8a; 
        10'b1100001100: data <= 18'h3ffb3; 
        10'b1100001101: data <= 18'h3ff8e; 
        10'b1100001110: data <= 18'h3ffb0; 
        10'b1100001111: data <= 18'h00016; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 13) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 19'h7ffa5; 
        10'b0000000001: data <= 19'h000ba; 
        10'b0000000010: data <= 19'h7ff2e; 
        10'b0000000011: data <= 19'h7fff0; 
        10'b0000000100: data <= 19'h7fff9; 
        10'b0000000101: data <= 19'h7ffe4; 
        10'b0000000110: data <= 19'h00062; 
        10'b0000000111: data <= 19'h00127; 
        10'b0000001000: data <= 19'h7ff3e; 
        10'b0000001001: data <= 19'h7ff7f; 
        10'b0000001010: data <= 19'h7ff88; 
        10'b0000001011: data <= 19'h7ff47; 
        10'b0000001100: data <= 19'h00060; 
        10'b0000001101: data <= 19'h0010d; 
        10'b0000001110: data <= 19'h00097; 
        10'b0000001111: data <= 19'h7ff0a; 
        10'b0000010000: data <= 19'h7ffde; 
        10'b0000010001: data <= 19'h00127; 
        10'b0000010010: data <= 19'h00032; 
        10'b0000010011: data <= 19'h7ffe6; 
        10'b0000010100: data <= 19'h7ff1d; 
        10'b0000010101: data <= 19'h7ff68; 
        10'b0000010110: data <= 19'h00046; 
        10'b0000010111: data <= 19'h00103; 
        10'b0000011000: data <= 19'h0008b; 
        10'b0000011001: data <= 19'h000aa; 
        10'b0000011010: data <= 19'h7ff1a; 
        10'b0000011011: data <= 19'h7ff23; 
        10'b0000011100: data <= 19'h000be; 
        10'b0000011101: data <= 19'h00096; 
        10'b0000011110: data <= 19'h000bf; 
        10'b0000011111: data <= 19'h7ffcf; 
        10'b0000100000: data <= 19'h7fefe; 
        10'b0000100001: data <= 19'h7ff66; 
        10'b0000100010: data <= 19'h00084; 
        10'b0000100011: data <= 19'h001ad; 
        10'b0000100100: data <= 19'h00123; 
        10'b0000100101: data <= 19'h00057; 
        10'b0000100110: data <= 19'h00160; 
        10'b0000100111: data <= 19'h00178; 
        10'b0000101000: data <= 19'h00191; 
        10'b0000101001: data <= 19'h00179; 
        10'b0000101010: data <= 19'h000ee; 
        10'b0000101011: data <= 19'h000fe; 
        10'b0000101100: data <= 19'h7fef1; 
        10'b0000101101: data <= 19'h000f2; 
        10'b0000101110: data <= 19'h00148; 
        10'b0000101111: data <= 19'h000bb; 
        10'b0000110000: data <= 19'h7ffcb; 
        10'b0000110001: data <= 19'h7ff59; 
        10'b0000110010: data <= 19'h0015c; 
        10'b0000110011: data <= 19'h00107; 
        10'b0000110100: data <= 19'h7ff94; 
        10'b0000110101: data <= 19'h00125; 
        10'b0000110110: data <= 19'h7ffcd; 
        10'b0000110111: data <= 19'h000d9; 
        10'b0000111000: data <= 19'h7ff55; 
        10'b0000111001: data <= 19'h7ff32; 
        10'b0000111010: data <= 19'h7fefd; 
        10'b0000111011: data <= 19'h7ffe7; 
        10'b0000111100: data <= 19'h00092; 
        10'b0000111101: data <= 19'h0005a; 
        10'b0000111110: data <= 19'h00095; 
        10'b0000111111: data <= 19'h001a4; 
        10'b0001000000: data <= 19'h0012b; 
        10'b0001000001: data <= 19'h0027c; 
        10'b0001000010: data <= 19'h00321; 
        10'b0001000011: data <= 19'h00389; 
        10'b0001000100: data <= 19'h0038b; 
        10'b0001000101: data <= 19'h003b8; 
        10'b0001000110: data <= 19'h001e3; 
        10'b0001000111: data <= 19'h00156; 
        10'b0001001000: data <= 19'h0031b; 
        10'b0001001001: data <= 19'h0015f; 
        10'b0001001010: data <= 19'h00155; 
        10'b0001001011: data <= 19'h00176; 
        10'b0001001100: data <= 19'h0016d; 
        10'b0001001101: data <= 19'h000b9; 
        10'b0001001110: data <= 19'h000f4; 
        10'b0001001111: data <= 19'h0002e; 
        10'b0001010000: data <= 19'h00086; 
        10'b0001010001: data <= 19'h7ffb4; 
        10'b0001010010: data <= 19'h7fef2; 
        10'b0001010011: data <= 19'h00053; 
        10'b0001010100: data <= 19'h7ff1b; 
        10'b0001010101: data <= 19'h0001b; 
        10'b0001010110: data <= 19'h000d8; 
        10'b0001010111: data <= 19'h0007d; 
        10'b0001011000: data <= 19'h0011b; 
        10'b0001011001: data <= 19'h7ff0a; 
        10'b0001011010: data <= 19'h00133; 
        10'b0001011011: data <= 19'h00150; 
        10'b0001011100: data <= 19'h00190; 
        10'b0001011101: data <= 19'h0032b; 
        10'b0001011110: data <= 19'h002cf; 
        10'b0001011111: data <= 19'h00384; 
        10'b0001100000: data <= 19'h0036e; 
        10'b0001100001: data <= 19'h0034d; 
        10'b0001100010: data <= 19'h004dc; 
        10'b0001100011: data <= 19'h00495; 
        10'b0001100100: data <= 19'h002d9; 
        10'b0001100101: data <= 19'h00399; 
        10'b0001100110: data <= 19'h005c7; 
        10'b0001100111: data <= 19'h005c3; 
        10'b0001101000: data <= 19'h00625; 
        10'b0001101001: data <= 19'h00572; 
        10'b0001101010: data <= 19'h00583; 
        10'b0001101011: data <= 19'h00334; 
        10'b0001101100: data <= 19'h002d7; 
        10'b0001101101: data <= 19'h000b2; 
        10'b0001101110: data <= 19'h7ff83; 
        10'b0001101111: data <= 19'h000a1; 
        10'b0001110000: data <= 19'h0002a; 
        10'b0001110001: data <= 19'h7ffca; 
        10'b0001110010: data <= 19'h7ffed; 
        10'b0001110011: data <= 19'h000fa; 
        10'b0001110100: data <= 19'h000d7; 
        10'b0001110101: data <= 19'h0004f; 
        10'b0001110110: data <= 19'h00050; 
        10'b0001110111: data <= 19'h001f7; 
        10'b0001111000: data <= 19'h7ffc8; 
        10'b0001111001: data <= 19'h7ff97; 
        10'b0001111010: data <= 19'h001e6; 
        10'b0001111011: data <= 19'h000b7; 
        10'b0001111100: data <= 19'h000e1; 
        10'b0001111101: data <= 19'h00051; 
        10'b0001111110: data <= 19'h000bf; 
        10'b0001111111: data <= 19'h00120; 
        10'b0010000000: data <= 19'h003da; 
        10'b0010000001: data <= 19'h003d0; 
        10'b0010000010: data <= 19'h005f9; 
        10'b0010000011: data <= 19'h00612; 
        10'b0010000100: data <= 19'h007a9; 
        10'b0010000101: data <= 19'h00880; 
        10'b0010000110: data <= 19'h00750; 
        10'b0010000111: data <= 19'h004e9; 
        10'b0010001000: data <= 19'h000b2; 
        10'b0010001001: data <= 19'h0014e; 
        10'b0010001010: data <= 19'h0002e; 
        10'b0010001011: data <= 19'h00000; 
        10'b0010001100: data <= 19'h00032; 
        10'b0010001101: data <= 19'h00098; 
        10'b0010001110: data <= 19'h00057; 
        10'b0010001111: data <= 19'h7ff8c; 
        10'b0010010000: data <= 19'h7ff30; 
        10'b0010010001: data <= 19'h7ffe9; 
        10'b0010010010: data <= 19'h7ff52; 
        10'b0010010011: data <= 19'h7fea8; 
        10'b0010010100: data <= 19'h00102; 
        10'b0010010101: data <= 19'h7feb3; 
        10'b0010010110: data <= 19'h00078; 
        10'b0010010111: data <= 19'h7fb8a; 
        10'b0010011000: data <= 19'h7fda4; 
        10'b0010011001: data <= 19'h7fe5e; 
        10'b0010011010: data <= 19'h7ff67; 
        10'b0010011011: data <= 19'h7fde5; 
        10'b0010011100: data <= 19'h7fde5; 
        10'b0010011101: data <= 19'h00068; 
        10'b0010011110: data <= 19'h002dd; 
        10'b0010011111: data <= 19'h0055f; 
        10'b0010100000: data <= 19'h004a9; 
        10'b0010100001: data <= 19'h0042a; 
        10'b0010100010: data <= 19'h00349; 
        10'b0010100011: data <= 19'h00241; 
        10'b0010100100: data <= 19'h7ffbd; 
        10'b0010100101: data <= 19'h0001d; 
        10'b0010100110: data <= 19'h7fede; 
        10'b0010100111: data <= 19'h00112; 
        10'b0010101000: data <= 19'h7ffda; 
        10'b0010101001: data <= 19'h000f7; 
        10'b0010101010: data <= 19'h000e6; 
        10'b0010101011: data <= 19'h7fed7; 
        10'b0010101100: data <= 19'h00069; 
        10'b0010101101: data <= 19'h7ffd1; 
        10'b0010101110: data <= 19'h0005f; 
        10'b0010101111: data <= 19'h00007; 
        10'b0010110000: data <= 19'h7fe58; 
        10'b0010110001: data <= 19'h7fdfb; 
        10'b0010110010: data <= 19'h7fadd; 
        10'b0010110011: data <= 19'h7f949; 
        10'b0010110100: data <= 19'h7fc19; 
        10'b0010110101: data <= 19'h7f858; 
        10'b0010110110: data <= 19'h7fc9f; 
        10'b0010110111: data <= 19'h7fd85; 
        10'b0010111000: data <= 19'h7fc78; 
        10'b0010111001: data <= 19'h7fce1; 
        10'b0010111010: data <= 19'h7ff22; 
        10'b0010111011: data <= 19'h7fde8; 
        10'b0010111100: data <= 19'h7fc9b; 
        10'b0010111101: data <= 19'h7fcc4; 
        10'b0010111110: data <= 19'h7faf8; 
        10'b0010111111: data <= 19'h7fcb8; 
        10'b0011000000: data <= 19'h7fd47; 
        10'b0011000001: data <= 19'h7fd22; 
        10'b0011000010: data <= 19'h7ff92; 
        10'b0011000011: data <= 19'h000ef; 
        10'b0011000100: data <= 19'h0005f; 
        10'b0011000101: data <= 19'h0008e; 
        10'b0011000110: data <= 19'h00009; 
        10'b0011000111: data <= 19'h7ffd1; 
        10'b0011001000: data <= 19'h00010; 
        10'b0011001001: data <= 19'h7ff01; 
        10'b0011001010: data <= 19'h7fdfc; 
        10'b0011001011: data <= 19'h7ffad; 
        10'b0011001100: data <= 19'h7fd23; 
        10'b0011001101: data <= 19'h7fc72; 
        10'b0011001110: data <= 19'h7fad3; 
        10'b0011001111: data <= 19'h7fbef; 
        10'b0011010000: data <= 19'h7f8b1; 
        10'b0011010001: data <= 19'h7f7cf; 
        10'b0011010010: data <= 19'h7fbb4; 
        10'b0011010011: data <= 19'h7fbed; 
        10'b0011010100: data <= 19'h7f99d; 
        10'b0011010101: data <= 19'h7f9f4; 
        10'b0011010110: data <= 19'h7f881; 
        10'b0011010111: data <= 19'h7f5d4; 
        10'b0011011000: data <= 19'h7f59f; 
        10'b0011011001: data <= 19'h7f752; 
        10'b0011011010: data <= 19'h7f6eb; 
        10'b0011011011: data <= 19'h7f8d4; 
        10'b0011011100: data <= 19'h7fd42; 
        10'b0011011101: data <= 19'h7fd85; 
        10'b0011011110: data <= 19'h7ff05; 
        10'b0011011111: data <= 19'h7ff41; 
        10'b0011100000: data <= 19'h7ffa4; 
        10'b0011100001: data <= 19'h7ffb2; 
        10'b0011100010: data <= 19'h00119; 
        10'b0011100011: data <= 19'h7fe99; 
        10'b0011100100: data <= 19'h7fed5; 
        10'b0011100101: data <= 19'h7fe72; 
        10'b0011100110: data <= 19'h7fc1a; 
        10'b0011100111: data <= 19'h7ff25; 
        10'b0011101000: data <= 19'h7fe90; 
        10'b0011101001: data <= 19'h7fbec; 
        10'b0011101010: data <= 19'h7fb3d; 
        10'b0011101011: data <= 19'h7fa8b; 
        10'b0011101100: data <= 19'h7f96e; 
        10'b0011101101: data <= 19'h7f862; 
        10'b0011101110: data <= 19'h7f894; 
        10'b0011101111: data <= 19'h7f812; 
        10'b0011110000: data <= 19'h7f699; 
        10'b0011110001: data <= 19'h7f52b; 
        10'b0011110010: data <= 19'h7f0b2; 
        10'b0011110011: data <= 19'h7f1c1; 
        10'b0011110100: data <= 19'h7f343; 
        10'b0011110101: data <= 19'h7f363; 
        10'b0011110110: data <= 19'h7f72f; 
        10'b0011110111: data <= 19'h7f83c; 
        10'b0011111000: data <= 19'h7fb27; 
        10'b0011111001: data <= 19'h7fcf2; 
        10'b0011111010: data <= 19'h7fdcf; 
        10'b0011111011: data <= 19'h00053; 
        10'b0011111100: data <= 19'h7ffd7; 
        10'b0011111101: data <= 19'h7ff26; 
        10'b0011111110: data <= 19'h7ff83; 
        10'b0011111111: data <= 19'h7ff07; 
        10'b0100000000: data <= 19'h00007; 
        10'b0100000001: data <= 19'h7ff1b; 
        10'b0100000010: data <= 19'h7fea4; 
        10'b0100000011: data <= 19'h7ff36; 
        10'b0100000100: data <= 19'h000ee; 
        10'b0100000101: data <= 19'h7fd8a; 
        10'b0100000110: data <= 19'h7fb59; 
        10'b0100000111: data <= 19'h7fc6e; 
        10'b0100001000: data <= 19'h7fdb4; 
        10'b0100001001: data <= 19'h7fbaa; 
        10'b0100001010: data <= 19'h7fc07; 
        10'b0100001011: data <= 19'h7f750; 
        10'b0100001100: data <= 19'h7f5e1; 
        10'b0100001101: data <= 19'h7f156; 
        10'b0100001110: data <= 19'h7f05c; 
        10'b0100001111: data <= 19'h7f33a; 
        10'b0100010000: data <= 19'h7f586; 
        10'b0100010001: data <= 19'h7f7aa; 
        10'b0100010010: data <= 19'h7f659; 
        10'b0100010011: data <= 19'h7f9cc; 
        10'b0100010100: data <= 19'h7fb44; 
        10'b0100010101: data <= 19'h7fc7d; 
        10'b0100010110: data <= 19'h7fe8e; 
        10'b0100010111: data <= 19'h000c2; 
        10'b0100011000: data <= 19'h7ff44; 
        10'b0100011001: data <= 19'h000f6; 
        10'b0100011010: data <= 19'h000a6; 
        10'b0100011011: data <= 19'h7fee0; 
        10'b0100011100: data <= 19'h7fe5d; 
        10'b0100011101: data <= 19'h0006a; 
        10'b0100011110: data <= 19'h0015a; 
        10'b0100011111: data <= 19'h0014c; 
        10'b0100100000: data <= 19'h004c0; 
        10'b0100100001: data <= 19'h7ffe7; 
        10'b0100100010: data <= 19'h000f2; 
        10'b0100100011: data <= 19'h00065; 
        10'b0100100100: data <= 19'h7fd20; 
        10'b0100100101: data <= 19'h7fe0c; 
        10'b0100100110: data <= 19'h7fbb7; 
        10'b0100100111: data <= 19'h7f702; 
        10'b0100101000: data <= 19'h7f6db; 
        10'b0100101001: data <= 19'h7f547; 
        10'b0100101010: data <= 19'h7f4d6; 
        10'b0100101011: data <= 19'h7f716; 
        10'b0100101100: data <= 19'h7f9f3; 
        10'b0100101101: data <= 19'h7fbab; 
        10'b0100101110: data <= 19'h7fa4c; 
        10'b0100101111: data <= 19'h7ff67; 
        10'b0100110000: data <= 19'h7fc4a; 
        10'b0100110001: data <= 19'h7fd6c; 
        10'b0100110010: data <= 19'h7ff3c; 
        10'b0100110011: data <= 19'h7ffa1; 
        10'b0100110100: data <= 19'h7ff67; 
        10'b0100110101: data <= 19'h00064; 
        10'b0100110110: data <= 19'h7ff58; 
        10'b0100110111: data <= 19'h7ffe8; 
        10'b0100111000: data <= 19'h7ff5a; 
        10'b0100111001: data <= 19'h0002b; 
        10'b0100111010: data <= 19'h7ffa6; 
        10'b0100111011: data <= 19'h003f9; 
        10'b0100111100: data <= 19'h002d8; 
        10'b0100111101: data <= 19'h0015e; 
        10'b0100111110: data <= 19'h001b8; 
        10'b0100111111: data <= 19'h00137; 
        10'b0101000000: data <= 19'h00138; 
        10'b0101000001: data <= 19'h00032; 
        10'b0101000010: data <= 19'h7fdee; 
        10'b0101000011: data <= 19'h7f8de; 
        10'b0101000100: data <= 19'h7f950; 
        10'b0101000101: data <= 19'h7fa4f; 
        10'b0101000110: data <= 19'h7fa48; 
        10'b0101000111: data <= 19'h7fb8d; 
        10'b0101001000: data <= 19'h7fdec; 
        10'b0101001001: data <= 19'h000cd; 
        10'b0101001010: data <= 19'h002ba; 
        10'b0101001011: data <= 19'h0043e; 
        10'b0101001100: data <= 19'h7fffd; 
        10'b0101001101: data <= 19'h7fdbe; 
        10'b0101001110: data <= 19'h7ff0f; 
        10'b0101001111: data <= 19'h7ffa8; 
        10'b0101010000: data <= 19'h7ff67; 
        10'b0101010001: data <= 19'h7ffae; 
        10'b0101010010: data <= 19'h7ff07; 
        10'b0101010011: data <= 19'h7ff89; 
        10'b0101010100: data <= 19'h00091; 
        10'b0101010101: data <= 19'h001dc; 
        10'b0101010110: data <= 19'h002d7; 
        10'b0101010111: data <= 19'h003ba; 
        10'b0101011000: data <= 19'h001ba; 
        10'b0101011001: data <= 19'h0026c; 
        10'b0101011010: data <= 19'h001b5; 
        10'b0101011011: data <= 19'h0047e; 
        10'b0101011100: data <= 19'h00452; 
        10'b0101011101: data <= 19'h00318; 
        10'b0101011110: data <= 19'h7fd5a; 
        10'b0101011111: data <= 19'h7fb37; 
        10'b0101100000: data <= 19'h7ffcd; 
        10'b0101100001: data <= 19'h7ff8f; 
        10'b0101100010: data <= 19'h7fb51; 
        10'b0101100011: data <= 19'h7fb83; 
        10'b0101100100: data <= 19'h7ff71; 
        10'b0101100101: data <= 19'h00289; 
        10'b0101100110: data <= 19'h00620; 
        10'b0101100111: data <= 19'h00ade; 
        10'b0101101000: data <= 19'h005d8; 
        10'b0101101001: data <= 19'h7fe55; 
        10'b0101101010: data <= 19'h7fe16; 
        10'b0101101011: data <= 19'h7ff6c; 
        10'b0101101100: data <= 19'h7ff6e; 
        10'b0101101101: data <= 19'h00102; 
        10'b0101101110: data <= 19'h000c5; 
        10'b0101101111: data <= 19'h7fee7; 
        10'b0101110000: data <= 19'h7fe80; 
        10'b0101110001: data <= 19'h0009b; 
        10'b0101110010: data <= 19'h004b7; 
        10'b0101110011: data <= 19'h0028a; 
        10'b0101110100: data <= 19'h0022e; 
        10'b0101110101: data <= 19'h00114; 
        10'b0101110110: data <= 19'h00494; 
        10'b0101110111: data <= 19'h003d2; 
        10'b0101111000: data <= 19'h00381; 
        10'b0101111001: data <= 19'h0009e; 
        10'b0101111010: data <= 19'h7ff5a; 
        10'b0101111011: data <= 19'h7ffe3; 
        10'b0101111100: data <= 19'h0005b; 
        10'b0101111101: data <= 19'h7fef8; 
        10'b0101111110: data <= 19'h7fbec; 
        10'b0101111111: data <= 19'h7ff77; 
        10'b0110000000: data <= 19'h7fe0a; 
        10'b0110000001: data <= 19'h00343; 
        10'b0110000010: data <= 19'h0087b; 
        10'b0110000011: data <= 19'h00d70; 
        10'b0110000100: data <= 19'h00742; 
        10'b0110000101: data <= 19'h7ff6c; 
        10'b0110000110: data <= 19'h00006; 
        10'b0110000111: data <= 19'h000a9; 
        10'b0110001000: data <= 19'h7ff85; 
        10'b0110001001: data <= 19'h0001b; 
        10'b0110001010: data <= 19'h000c3; 
        10'b0110001011: data <= 19'h0000a; 
        10'b0110001100: data <= 19'h7fe6a; 
        10'b0110001101: data <= 19'h001b1; 
        10'b0110001110: data <= 19'h00453; 
        10'b0110001111: data <= 19'h003ba; 
        10'b0110010000: data <= 19'h00521; 
        10'b0110010001: data <= 19'h004ce; 
        10'b0110010010: data <= 19'h00533; 
        10'b0110010011: data <= 19'h005a2; 
        10'b0110010100: data <= 19'h001e5; 
        10'b0110010101: data <= 19'h7fd41; 
        10'b0110010110: data <= 19'h0002f; 
        10'b0110010111: data <= 19'h0024b; 
        10'b0110011000: data <= 19'h00116; 
        10'b0110011001: data <= 19'h7fe37; 
        10'b0110011010: data <= 19'h7fe44; 
        10'b0110011011: data <= 19'h7ffc0; 
        10'b0110011100: data <= 19'h003ae; 
        10'b0110011101: data <= 19'h003a3; 
        10'b0110011110: data <= 19'h0099a; 
        10'b0110011111: data <= 19'h00b2c; 
        10'b0110100000: data <= 19'h00753; 
        10'b0110100001: data <= 19'h7ffe6; 
        10'b0110100010: data <= 19'h7fde7; 
        10'b0110100011: data <= 19'h7fef8; 
        10'b0110100100: data <= 19'h000c9; 
        10'b0110100101: data <= 19'h7ff9a; 
        10'b0110100110: data <= 19'h00027; 
        10'b0110100111: data <= 19'h7ff22; 
        10'b0110101000: data <= 19'h7fcf8; 
        10'b0110101001: data <= 19'h7ff9e; 
        10'b0110101010: data <= 19'h00482; 
        10'b0110101011: data <= 19'h005fe; 
        10'b0110101100: data <= 19'h003dc; 
        10'b0110101101: data <= 19'h0060f; 
        10'b0110101110: data <= 19'h007a3; 
        10'b0110101111: data <= 19'h00951; 
        10'b0110110000: data <= 19'h0026f; 
        10'b0110110001: data <= 19'h7ff53; 
        10'b0110110010: data <= 19'h00398; 
        10'b0110110011: data <= 19'h0034e; 
        10'b0110110100: data <= 19'h00083; 
        10'b0110110101: data <= 19'h7fe4e; 
        10'b0110110110: data <= 19'h00057; 
        10'b0110110111: data <= 19'h001db; 
        10'b0110111000: data <= 19'h0044e; 
        10'b0110111001: data <= 19'h005e9; 
        10'b0110111010: data <= 19'h0056e; 
        10'b0110111011: data <= 19'h006ba; 
        10'b0110111100: data <= 19'h00397; 
        10'b0110111101: data <= 19'h7fe29; 
        10'b0110111110: data <= 19'h7fedb; 
        10'b0110111111: data <= 19'h7fed4; 
        10'b0111000000: data <= 19'h00035; 
        10'b0111000001: data <= 19'h7ff25; 
        10'b0111000010: data <= 19'h7ff1d; 
        10'b0111000011: data <= 19'h7ff05; 
        10'b0111000100: data <= 19'h7fbfe; 
        10'b0111000101: data <= 19'h7fdd4; 
        10'b0111000110: data <= 19'h006ae; 
        10'b0111000111: data <= 19'h006d3; 
        10'b0111001000: data <= 19'h00484; 
        10'b0111001001: data <= 19'h006f8; 
        10'b0111001010: data <= 19'h00bd1; 
        10'b0111001011: data <= 19'h00bb9; 
        10'b0111001100: data <= 19'h00393; 
        10'b0111001101: data <= 19'h00220; 
        10'b0111001110: data <= 19'h00518; 
        10'b0111001111: data <= 19'h002b0; 
        10'b0111010000: data <= 19'h7fe98; 
        10'b0111010001: data <= 19'h7fd37; 
        10'b0111010010: data <= 19'h000f7; 
        10'b0111010011: data <= 19'h002fa; 
        10'b0111010100: data <= 19'h00163; 
        10'b0111010101: data <= 19'h0000a; 
        10'b0111010110: data <= 19'h002c8; 
        10'b0111010111: data <= 19'h001ab; 
        10'b0111011000: data <= 19'h7ff31; 
        10'b0111011001: data <= 19'h7fdd6; 
        10'b0111011010: data <= 19'h7feac; 
        10'b0111011011: data <= 19'h7ffd2; 
        10'b0111011100: data <= 19'h00032; 
        10'b0111011101: data <= 19'h000a8; 
        10'b0111011110: data <= 19'h000e8; 
        10'b0111011111: data <= 19'h7ffd7; 
        10'b0111100000: data <= 19'h7fa49; 
        10'b0111100001: data <= 19'h7fd03; 
        10'b0111100010: data <= 19'h002cb; 
        10'b0111100011: data <= 19'h0054f; 
        10'b0111100100: data <= 19'h0060a; 
        10'b0111100101: data <= 19'h0079e; 
        10'b0111100110: data <= 19'h00d26; 
        10'b0111100111: data <= 19'h00d5c; 
        10'b0111101000: data <= 19'h006e7; 
        10'b0111101001: data <= 19'h003e3; 
        10'b0111101010: data <= 19'h003ef; 
        10'b0111101011: data <= 19'h0027c; 
        10'b0111101100: data <= 19'h00000; 
        10'b0111101101: data <= 19'h000b8; 
        10'b0111101110: data <= 19'h0057a; 
        10'b0111101111: data <= 19'h001e4; 
        10'b0111110000: data <= 19'h000c9; 
        10'b0111110001: data <= 19'h7fe9a; 
        10'b0111110010: data <= 19'h00141; 
        10'b0111110011: data <= 19'h7ffbc; 
        10'b0111110100: data <= 19'h7fe72; 
        10'b0111110101: data <= 19'h7fcf8; 
        10'b0111110110: data <= 19'h7ff91; 
        10'b0111110111: data <= 19'h0007f; 
        10'b0111111000: data <= 19'h7ff8e; 
        10'b0111111001: data <= 19'h7ff62; 
        10'b0111111010: data <= 19'h7fffc; 
        10'b0111111011: data <= 19'h7fe55; 
        10'b0111111100: data <= 19'h7faa3; 
        10'b0111111101: data <= 19'h7fac4; 
        10'b0111111110: data <= 19'h7fd77; 
        10'b0111111111: data <= 19'h003a7; 
        10'b1000000000: data <= 19'h005da; 
        10'b1000000001: data <= 19'h00551; 
        10'b1000000010: data <= 19'h00935; 
        10'b1000000011: data <= 19'h00b5b; 
        10'b1000000100: data <= 19'h00d62; 
        10'b1000000101: data <= 19'h00637; 
        10'b1000000110: data <= 19'h001ae; 
        10'b1000000111: data <= 19'h00375; 
        10'b1000001000: data <= 19'h005f8; 
        10'b1000001001: data <= 19'h003e0; 
        10'b1000001010: data <= 19'h004d3; 
        10'b1000001011: data <= 19'h0028a; 
        10'b1000001100: data <= 19'h00054; 
        10'b1000001101: data <= 19'h000d9; 
        10'b1000001110: data <= 19'h000f0; 
        10'b1000001111: data <= 19'h7ff78; 
        10'b1000010000: data <= 19'h7fe17; 
        10'b1000010001: data <= 19'h7fe97; 
        10'b1000010010: data <= 19'h7fee9; 
        10'b1000010011: data <= 19'h7fed7; 
        10'b1000010100: data <= 19'h00049; 
        10'b1000010101: data <= 19'h7ff31; 
        10'b1000010110: data <= 19'h00083; 
        10'b1000010111: data <= 19'h7fde2; 
        10'b1000011000: data <= 19'h7fc87; 
        10'b1000011001: data <= 19'h7fa6e; 
        10'b1000011010: data <= 19'h7fbac; 
        10'b1000011011: data <= 19'h0004e; 
        10'b1000011100: data <= 19'h003cc; 
        10'b1000011101: data <= 19'h005f7; 
        10'b1000011110: data <= 19'h007f1; 
        10'b1000011111: data <= 19'h00ca9; 
        10'b1000100000: data <= 19'h00e3f; 
        10'b1000100001: data <= 19'h00758; 
        10'b1000100010: data <= 19'h0068f; 
        10'b1000100011: data <= 19'h006dc; 
        10'b1000100100: data <= 19'h004e2; 
        10'b1000100101: data <= 19'h00403; 
        10'b1000100110: data <= 19'h00643; 
        10'b1000100111: data <= 19'h00444; 
        10'b1000101000: data <= 19'h002c3; 
        10'b1000101001: data <= 19'h00098; 
        10'b1000101010: data <= 19'h7ff00; 
        10'b1000101011: data <= 19'h7fec4; 
        10'b1000101100: data <= 19'h7feb5; 
        10'b1000101101: data <= 19'h7ffcb; 
        10'b1000101110: data <= 19'h7ff62; 
        10'b1000101111: data <= 19'h000e9; 
        10'b1000110000: data <= 19'h7ff71; 
        10'b1000110001: data <= 19'h7ff30; 
        10'b1000110010: data <= 19'h7ffb7; 
        10'b1000110011: data <= 19'h7ff0a; 
        10'b1000110100: data <= 19'h7fb8f; 
        10'b1000110101: data <= 19'h7fab0; 
        10'b1000110110: data <= 19'h7fb66; 
        10'b1000110111: data <= 19'h7fe1f; 
        10'b1000111000: data <= 19'h00142; 
        10'b1000111001: data <= 19'h003fe; 
        10'b1000111010: data <= 19'h00693; 
        10'b1000111011: data <= 19'h00462; 
        10'b1000111100: data <= 19'h008a1; 
        10'b1000111101: data <= 19'h00a59; 
        10'b1000111110: data <= 19'h00c48; 
        10'b1000111111: data <= 19'h00a75; 
        10'b1001000000: data <= 19'h005ab; 
        10'b1001000001: data <= 19'h003a0; 
        10'b1001000010: data <= 19'h0070a; 
        10'b1001000011: data <= 19'h004f7; 
        10'b1001000100: data <= 19'h0035e; 
        10'b1001000101: data <= 19'h7ff4f; 
        10'b1001000110: data <= 19'h7fd64; 
        10'b1001000111: data <= 19'h0002b; 
        10'b1001001000: data <= 19'h7ff5e; 
        10'b1001001001: data <= 19'h7ffaf; 
        10'b1001001010: data <= 19'h7ff36; 
        10'b1001001011: data <= 19'h0002b; 
        10'b1001001100: data <= 19'h7ffe6; 
        10'b1001001101: data <= 19'h0001a; 
        10'b1001001110: data <= 19'h00055; 
        10'b1001001111: data <= 19'h7ffa9; 
        10'b1001010000: data <= 19'h7fe51; 
        10'b1001010001: data <= 19'h7fc57; 
        10'b1001010010: data <= 19'h7f9ca; 
        10'b1001010011: data <= 19'h7fd30; 
        10'b1001010100: data <= 19'h7fe51; 
        10'b1001010101: data <= 19'h00301; 
        10'b1001010110: data <= 19'h00575; 
        10'b1001010111: data <= 19'h007c3; 
        10'b1001011000: data <= 19'h009fc; 
        10'b1001011001: data <= 19'h00a23; 
        10'b1001011010: data <= 19'h00883; 
        10'b1001011011: data <= 19'h00756; 
        10'b1001011100: data <= 19'h00494; 
        10'b1001011101: data <= 19'h00643; 
        10'b1001011110: data <= 19'h005d6; 
        10'b1001011111: data <= 19'h003bb; 
        10'b1001100000: data <= 19'h0007f; 
        10'b1001100001: data <= 19'h7fe06; 
        10'b1001100010: data <= 19'h7fd3b; 
        10'b1001100011: data <= 19'h7fe64; 
        10'b1001100100: data <= 19'h00018; 
        10'b1001100101: data <= 19'h7fef5; 
        10'b1001100110: data <= 19'h7ffc6; 
        10'b1001100111: data <= 19'h7ff6c; 
        10'b1001101000: data <= 19'h7ff6b; 
        10'b1001101001: data <= 19'h7ffe6; 
        10'b1001101010: data <= 19'h000ff; 
        10'b1001101011: data <= 19'h00045; 
        10'b1001101100: data <= 19'h7ff6a; 
        10'b1001101101: data <= 19'h7fcd0; 
        10'b1001101110: data <= 19'h7fc37; 
        10'b1001101111: data <= 19'h7faec; 
        10'b1001110000: data <= 19'h7fc9d; 
        10'b1001110001: data <= 19'h7fe76; 
        10'b1001110010: data <= 19'h7febd; 
        10'b1001110011: data <= 19'h0009d; 
        10'b1001110100: data <= 19'h002eb; 
        10'b1001110101: data <= 19'h00144; 
        10'b1001110110: data <= 19'h00110; 
        10'b1001110111: data <= 19'h00327; 
        10'b1001111000: data <= 19'h00258; 
        10'b1001111001: data <= 19'h00005; 
        10'b1001111010: data <= 19'h7ff37; 
        10'b1001111011: data <= 19'h7fc7b; 
        10'b1001111100: data <= 19'h7fc9d; 
        10'b1001111101: data <= 19'h7fd2e; 
        10'b1001111110: data <= 19'h7fd5e; 
        10'b1001111111: data <= 19'h7ffbf; 
        10'b1010000000: data <= 19'h7ff8a; 
        10'b1010000001: data <= 19'h7ff05; 
        10'b1010000010: data <= 19'h00113; 
        10'b1010000011: data <= 19'h0006a; 
        10'b1010000100: data <= 19'h000dd; 
        10'b1010000101: data <= 19'h7ffa9; 
        10'b1010000110: data <= 19'h7ff85; 
        10'b1010000111: data <= 19'h00019; 
        10'b1010001000: data <= 19'h0004e; 
        10'b1010001001: data <= 19'h7feaf; 
        10'b1010001010: data <= 19'h7fdf1; 
        10'b1010001011: data <= 19'h7fb7a; 
        10'b1010001100: data <= 19'h7fa48; 
        10'b1010001101: data <= 19'h7f7c6; 
        10'b1010001110: data <= 19'h7f7d1; 
        10'b1010001111: data <= 19'h7f676; 
        10'b1010010000: data <= 19'h7fa1f; 
        10'b1010010001: data <= 19'h7fb5e; 
        10'b1010010010: data <= 19'h7fc64; 
        10'b1010010011: data <= 19'h7faa2; 
        10'b1010010100: data <= 19'h7f8f2; 
        10'b1010010101: data <= 19'h7f800; 
        10'b1010010110: data <= 19'h7f9b1; 
        10'b1010010111: data <= 19'h7fd20; 
        10'b1010011000: data <= 19'h7fd13; 
        10'b1010011001: data <= 19'h7fd70; 
        10'b1010011010: data <= 19'h7ff16; 
        10'b1010011011: data <= 19'h00021; 
        10'b1010011100: data <= 19'h7feef; 
        10'b1010011101: data <= 19'h7ff1f; 
        10'b1010011110: data <= 19'h7ffa0; 
        10'b1010011111: data <= 19'h7ffe4; 
        10'b1010100000: data <= 19'h0009e; 
        10'b1010100001: data <= 19'h0007f; 
        10'b1010100010: data <= 19'h00057; 
        10'b1010100011: data <= 19'h7fefc; 
        10'b1010100100: data <= 19'h7ff32; 
        10'b1010100101: data <= 19'h7ff9f; 
        10'b1010100110: data <= 19'h7ff07; 
        10'b1010100111: data <= 19'h7fe6c; 
        10'b1010101000: data <= 19'h7fec1; 
        10'b1010101001: data <= 19'h7fe02; 
        10'b1010101010: data <= 19'h7fd04; 
        10'b1010101011: data <= 19'h7fc39; 
        10'b1010101100: data <= 19'h7fb9b; 
        10'b1010101101: data <= 19'h7fbb3; 
        10'b1010101110: data <= 19'h7fafb; 
        10'b1010101111: data <= 19'h7fafc; 
        10'b1010110000: data <= 19'h7fac2; 
        10'b1010110001: data <= 19'h7fbff; 
        10'b1010110010: data <= 19'h7fe9c; 
        10'b1010110011: data <= 19'h7feb5; 
        10'b1010110100: data <= 19'h7ff8c; 
        10'b1010110101: data <= 19'h7ff49; 
        10'b1010110110: data <= 19'h00088; 
        10'b1010110111: data <= 19'h7ffc5; 
        10'b1010111000: data <= 19'h7fef4; 
        10'b1010111001: data <= 19'h7ffac; 
        10'b1010111010: data <= 19'h7ff38; 
        10'b1010111011: data <= 19'h7ff3e; 
        10'b1010111100: data <= 19'h000fa; 
        10'b1010111101: data <= 19'h7ff17; 
        10'b1010111110: data <= 19'h00044; 
        10'b1010111111: data <= 19'h7ff89; 
        10'b1011000000: data <= 19'h7ff4a; 
        10'b1011000001: data <= 19'h7ffde; 
        10'b1011000010: data <= 19'h000a7; 
        10'b1011000011: data <= 19'h7fff3; 
        10'b1011000100: data <= 19'h7fee4; 
        10'b1011000101: data <= 19'h00067; 
        10'b1011000110: data <= 19'h7feeb; 
        10'b1011000111: data <= 19'h7ffd5; 
        10'b1011001000: data <= 19'h0000e; 
        10'b1011001001: data <= 19'h7fedb; 
        10'b1011001010: data <= 19'h7ff5e; 
        10'b1011001011: data <= 19'h7ff9d; 
        10'b1011001100: data <= 19'h7ffe5; 
        10'b1011001101: data <= 19'h7ff00; 
        10'b1011001110: data <= 19'h7ff6a; 
        10'b1011001111: data <= 19'h7fee6; 
        10'b1011010000: data <= 19'h7ff22; 
        10'b1011010001: data <= 19'h00023; 
        10'b1011010010: data <= 19'h7ff95; 
        10'b1011010011: data <= 19'h000cb; 
        10'b1011010100: data <= 19'h00120; 
        10'b1011010101: data <= 19'h000fe; 
        10'b1011010110: data <= 19'h0000c; 
        10'b1011010111: data <= 19'h000bf; 
        10'b1011011000: data <= 19'h0010e; 
        10'b1011011001: data <= 19'h7fff3; 
        10'b1011011010: data <= 19'h00031; 
        10'b1011011011: data <= 19'h7ffcd; 
        10'b1011011100: data <= 19'h7ff68; 
        10'b1011011101: data <= 19'h000e3; 
        10'b1011011110: data <= 19'h000ab; 
        10'b1011011111: data <= 19'h7ff6c; 
        10'b1011100000: data <= 19'h7ffa8; 
        10'b1011100001: data <= 19'h00080; 
        10'b1011100010: data <= 19'h7ff95; 
        10'b1011100011: data <= 19'h00038; 
        10'b1011100100: data <= 19'h7ff90; 
        10'b1011100101: data <= 19'h000a7; 
        10'b1011100110: data <= 19'h000b0; 
        10'b1011100111: data <= 19'h7ff1c; 
        10'b1011101000: data <= 19'h7ff52; 
        10'b1011101001: data <= 19'h000e6; 
        10'b1011101010: data <= 19'h000b5; 
        10'b1011101011: data <= 19'h7ffa7; 
        10'b1011101100: data <= 19'h000a2; 
        10'b1011101101: data <= 19'h7ffc3; 
        10'b1011101110: data <= 19'h7ffc0; 
        10'b1011101111: data <= 19'h00065; 
        10'b1011110000: data <= 19'h00073; 
        10'b1011110001: data <= 19'h7ffc8; 
        10'b1011110010: data <= 19'h7ff78; 
        10'b1011110011: data <= 19'h7ffb2; 
        10'b1011110100: data <= 19'h00105; 
        10'b1011110101: data <= 19'h7fff3; 
        10'b1011110110: data <= 19'h00093; 
        10'b1011110111: data <= 19'h7ff6b; 
        10'b1011111000: data <= 19'h0005b; 
        10'b1011111001: data <= 19'h7fff9; 
        10'b1011111010: data <= 19'h000f5; 
        10'b1011111011: data <= 19'h00023; 
        10'b1011111100: data <= 19'h7ffdf; 
        10'b1011111101: data <= 19'h7fee0; 
        10'b1011111110: data <= 19'h7ff3d; 
        10'b1011111111: data <= 19'h00059; 
        10'b1100000000: data <= 19'h7fefb; 
        10'b1100000001: data <= 19'h7ff26; 
        10'b1100000010: data <= 19'h7ff5b; 
        10'b1100000011: data <= 19'h7fef6; 
        10'b1100000100: data <= 19'h7ff4c; 
        10'b1100000101: data <= 19'h7ffa7; 
        10'b1100000110: data <= 19'h7ff12; 
        10'b1100000111: data <= 19'h7ff4c; 
        10'b1100001000: data <= 19'h7ff64; 
        10'b1100001001: data <= 19'h7ff81; 
        10'b1100001010: data <= 19'h000f1; 
        10'b1100001011: data <= 19'h7ff14; 
        10'b1100001100: data <= 19'h7ff66; 
        10'b1100001101: data <= 19'h7ff1c; 
        10'b1100001110: data <= 19'h7ff60; 
        10'b1100001111: data <= 19'h0002c; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 14) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 20'hfff4a; 
        10'b0000000001: data <= 20'h00174; 
        10'b0000000010: data <= 20'hffe5c; 
        10'b0000000011: data <= 20'hfffe0; 
        10'b0000000100: data <= 20'hffff2; 
        10'b0000000101: data <= 20'hfffc7; 
        10'b0000000110: data <= 20'h000c3; 
        10'b0000000111: data <= 20'h0024e; 
        10'b0000001000: data <= 20'hffe7d; 
        10'b0000001001: data <= 20'hffeff; 
        10'b0000001010: data <= 20'hfff0f; 
        10'b0000001011: data <= 20'hffe8e; 
        10'b0000001100: data <= 20'h000bf; 
        10'b0000001101: data <= 20'h0021b; 
        10'b0000001110: data <= 20'h0012f; 
        10'b0000001111: data <= 20'hffe13; 
        10'b0000010000: data <= 20'hfffbc; 
        10'b0000010001: data <= 20'h0024e; 
        10'b0000010010: data <= 20'h00064; 
        10'b0000010011: data <= 20'hfffcc; 
        10'b0000010100: data <= 20'hffe3a; 
        10'b0000010101: data <= 20'hffed1; 
        10'b0000010110: data <= 20'h0008b; 
        10'b0000010111: data <= 20'h00205; 
        10'b0000011000: data <= 20'h00117; 
        10'b0000011001: data <= 20'h00154; 
        10'b0000011010: data <= 20'hffe33; 
        10'b0000011011: data <= 20'hffe46; 
        10'b0000011100: data <= 20'h0017b; 
        10'b0000011101: data <= 20'h0012d; 
        10'b0000011110: data <= 20'h0017e; 
        10'b0000011111: data <= 20'hfff9f; 
        10'b0000100000: data <= 20'hffdfb; 
        10'b0000100001: data <= 20'hffecb; 
        10'b0000100010: data <= 20'h00108; 
        10'b0000100011: data <= 20'h0035b; 
        10'b0000100100: data <= 20'h00246; 
        10'b0000100101: data <= 20'h000af; 
        10'b0000100110: data <= 20'h002c0; 
        10'b0000100111: data <= 20'h002f0; 
        10'b0000101000: data <= 20'h00321; 
        10'b0000101001: data <= 20'h002f3; 
        10'b0000101010: data <= 20'h001db; 
        10'b0000101011: data <= 20'h001fc; 
        10'b0000101100: data <= 20'hffde1; 
        10'b0000101101: data <= 20'h001e4; 
        10'b0000101110: data <= 20'h00290; 
        10'b0000101111: data <= 20'h00176; 
        10'b0000110000: data <= 20'hfff96; 
        10'b0000110001: data <= 20'hffeb2; 
        10'b0000110010: data <= 20'h002b9; 
        10'b0000110011: data <= 20'h0020e; 
        10'b0000110100: data <= 20'hfff28; 
        10'b0000110101: data <= 20'h0024b; 
        10'b0000110110: data <= 20'hfff9b; 
        10'b0000110111: data <= 20'h001b2; 
        10'b0000111000: data <= 20'hffeaa; 
        10'b0000111001: data <= 20'hffe64; 
        10'b0000111010: data <= 20'hffdfa; 
        10'b0000111011: data <= 20'hfffcd; 
        10'b0000111100: data <= 20'h00124; 
        10'b0000111101: data <= 20'h000b4; 
        10'b0000111110: data <= 20'h0012a; 
        10'b0000111111: data <= 20'h00348; 
        10'b0001000000: data <= 20'h00255; 
        10'b0001000001: data <= 20'h004f9; 
        10'b0001000010: data <= 20'h00641; 
        10'b0001000011: data <= 20'h00711; 
        10'b0001000100: data <= 20'h00715; 
        10'b0001000101: data <= 20'h00771; 
        10'b0001000110: data <= 20'h003c6; 
        10'b0001000111: data <= 20'h002ad; 
        10'b0001001000: data <= 20'h00636; 
        10'b0001001001: data <= 20'h002be; 
        10'b0001001010: data <= 20'h002aa; 
        10'b0001001011: data <= 20'h002eb; 
        10'b0001001100: data <= 20'h002db; 
        10'b0001001101: data <= 20'h00172; 
        10'b0001001110: data <= 20'h001e7; 
        10'b0001001111: data <= 20'h0005b; 
        10'b0001010000: data <= 20'h0010c; 
        10'b0001010001: data <= 20'hfff67; 
        10'b0001010010: data <= 20'hffde5; 
        10'b0001010011: data <= 20'h000a5; 
        10'b0001010100: data <= 20'hffe37; 
        10'b0001010101: data <= 20'h00036; 
        10'b0001010110: data <= 20'h001af; 
        10'b0001010111: data <= 20'h000f9; 
        10'b0001011000: data <= 20'h00236; 
        10'b0001011001: data <= 20'hffe14; 
        10'b0001011010: data <= 20'h00266; 
        10'b0001011011: data <= 20'h002a1; 
        10'b0001011100: data <= 20'h00320; 
        10'b0001011101: data <= 20'h00656; 
        10'b0001011110: data <= 20'h0059d; 
        10'b0001011111: data <= 20'h00708; 
        10'b0001100000: data <= 20'h006dc; 
        10'b0001100001: data <= 20'h0069a; 
        10'b0001100010: data <= 20'h009b7; 
        10'b0001100011: data <= 20'h0092a; 
        10'b0001100100: data <= 20'h005b2; 
        10'b0001100101: data <= 20'h00731; 
        10'b0001100110: data <= 20'h00b8e; 
        10'b0001100111: data <= 20'h00b86; 
        10'b0001101000: data <= 20'h00c4b; 
        10'b0001101001: data <= 20'h00ae3; 
        10'b0001101010: data <= 20'h00b06; 
        10'b0001101011: data <= 20'h00667; 
        10'b0001101100: data <= 20'h005af; 
        10'b0001101101: data <= 20'h00164; 
        10'b0001101110: data <= 20'hfff06; 
        10'b0001101111: data <= 20'h00142; 
        10'b0001110000: data <= 20'h00055; 
        10'b0001110001: data <= 20'hfff95; 
        10'b0001110010: data <= 20'hfffda; 
        10'b0001110011: data <= 20'h001f4; 
        10'b0001110100: data <= 20'h001ae; 
        10'b0001110101: data <= 20'h0009d; 
        10'b0001110110: data <= 20'h0009f; 
        10'b0001110111: data <= 20'h003ed; 
        10'b0001111000: data <= 20'hfff90; 
        10'b0001111001: data <= 20'hfff2e; 
        10'b0001111010: data <= 20'h003cc; 
        10'b0001111011: data <= 20'h0016e; 
        10'b0001111100: data <= 20'h001c3; 
        10'b0001111101: data <= 20'h000a3; 
        10'b0001111110: data <= 20'h0017f; 
        10'b0001111111: data <= 20'h00240; 
        10'b0010000000: data <= 20'h007b4; 
        10'b0010000001: data <= 20'h007a0; 
        10'b0010000010: data <= 20'h00bf2; 
        10'b0010000011: data <= 20'h00c25; 
        10'b0010000100: data <= 20'h00f53; 
        10'b0010000101: data <= 20'h01100; 
        10'b0010000110: data <= 20'h00ea0; 
        10'b0010000111: data <= 20'h009d2; 
        10'b0010001000: data <= 20'h00164; 
        10'b0010001001: data <= 20'h0029b; 
        10'b0010001010: data <= 20'h0005d; 
        10'b0010001011: data <= 20'h00000; 
        10'b0010001100: data <= 20'h00065; 
        10'b0010001101: data <= 20'h00130; 
        10'b0010001110: data <= 20'h000ad; 
        10'b0010001111: data <= 20'hfff19; 
        10'b0010010000: data <= 20'hffe61; 
        10'b0010010001: data <= 20'hfffd2; 
        10'b0010010010: data <= 20'hffea4; 
        10'b0010010011: data <= 20'hffd4f; 
        10'b0010010100: data <= 20'h00204; 
        10'b0010010101: data <= 20'hffd67; 
        10'b0010010110: data <= 20'h000f0; 
        10'b0010010111: data <= 20'hff715; 
        10'b0010011000: data <= 20'hffb47; 
        10'b0010011001: data <= 20'hffcbd; 
        10'b0010011010: data <= 20'hffecd; 
        10'b0010011011: data <= 20'hffbca; 
        10'b0010011100: data <= 20'hffbca; 
        10'b0010011101: data <= 20'h000d0; 
        10'b0010011110: data <= 20'h005bb; 
        10'b0010011111: data <= 20'h00abe; 
        10'b0010100000: data <= 20'h00952; 
        10'b0010100001: data <= 20'h00855; 
        10'b0010100010: data <= 20'h00693; 
        10'b0010100011: data <= 20'h00482; 
        10'b0010100100: data <= 20'hfff7a; 
        10'b0010100101: data <= 20'h0003a; 
        10'b0010100110: data <= 20'hffdbc; 
        10'b0010100111: data <= 20'h00224; 
        10'b0010101000: data <= 20'hfffb5; 
        10'b0010101001: data <= 20'h001ed; 
        10'b0010101010: data <= 20'h001cc; 
        10'b0010101011: data <= 20'hffdae; 
        10'b0010101100: data <= 20'h000d2; 
        10'b0010101101: data <= 20'hfffa2; 
        10'b0010101110: data <= 20'h000be; 
        10'b0010101111: data <= 20'h0000e; 
        10'b0010110000: data <= 20'hffcb0; 
        10'b0010110001: data <= 20'hffbf6; 
        10'b0010110010: data <= 20'hff5ba; 
        10'b0010110011: data <= 20'hff292; 
        10'b0010110100: data <= 20'hff832; 
        10'b0010110101: data <= 20'hff0b0; 
        10'b0010110110: data <= 20'hff93f; 
        10'b0010110111: data <= 20'hffb0a; 
        10'b0010111000: data <= 20'hff8f0; 
        10'b0010111001: data <= 20'hff9c2; 
        10'b0010111010: data <= 20'hffe44; 
        10'b0010111011: data <= 20'hffbd0; 
        10'b0010111100: data <= 20'hff937; 
        10'b0010111101: data <= 20'hff988; 
        10'b0010111110: data <= 20'hff5f1; 
        10'b0010111111: data <= 20'hff970; 
        10'b0011000000: data <= 20'hffa8f; 
        10'b0011000001: data <= 20'hffa43; 
        10'b0011000010: data <= 20'hfff25; 
        10'b0011000011: data <= 20'h001df; 
        10'b0011000100: data <= 20'h000be; 
        10'b0011000101: data <= 20'h0011c; 
        10'b0011000110: data <= 20'h00011; 
        10'b0011000111: data <= 20'hfffa2; 
        10'b0011001000: data <= 20'h00020; 
        10'b0011001001: data <= 20'hffe02; 
        10'b0011001010: data <= 20'hffbf7; 
        10'b0011001011: data <= 20'hfff5a; 
        10'b0011001100: data <= 20'hffa46; 
        10'b0011001101: data <= 20'hff8e3; 
        10'b0011001110: data <= 20'hff5a6; 
        10'b0011001111: data <= 20'hff7dd; 
        10'b0011010000: data <= 20'hff161; 
        10'b0011010001: data <= 20'hfef9e; 
        10'b0011010010: data <= 20'hff769; 
        10'b0011010011: data <= 20'hff7da; 
        10'b0011010100: data <= 20'hff33a; 
        10'b0011010101: data <= 20'hff3e9; 
        10'b0011010110: data <= 20'hff102; 
        10'b0011010111: data <= 20'hfeba9; 
        10'b0011011000: data <= 20'hfeb3e; 
        10'b0011011001: data <= 20'hfeea3; 
        10'b0011011010: data <= 20'hfedd7; 
        10'b0011011011: data <= 20'hff1a8; 
        10'b0011011100: data <= 20'hffa84; 
        10'b0011011101: data <= 20'hffb0a; 
        10'b0011011110: data <= 20'hffe0b; 
        10'b0011011111: data <= 20'hffe81; 
        10'b0011100000: data <= 20'hfff47; 
        10'b0011100001: data <= 20'hfff63; 
        10'b0011100010: data <= 20'h00232; 
        10'b0011100011: data <= 20'hffd32; 
        10'b0011100100: data <= 20'hffdab; 
        10'b0011100101: data <= 20'hffce5; 
        10'b0011100110: data <= 20'hff834; 
        10'b0011100111: data <= 20'hffe4a; 
        10'b0011101000: data <= 20'hffd1f; 
        10'b0011101001: data <= 20'hff7d9; 
        10'b0011101010: data <= 20'hff67a; 
        10'b0011101011: data <= 20'hff516; 
        10'b0011101100: data <= 20'hff2dc; 
        10'b0011101101: data <= 20'hff0c3; 
        10'b0011101110: data <= 20'hff127; 
        10'b0011101111: data <= 20'hff024; 
        10'b0011110000: data <= 20'hfed32; 
        10'b0011110001: data <= 20'hfea57; 
        10'b0011110010: data <= 20'hfe164; 
        10'b0011110011: data <= 20'hfe382; 
        10'b0011110100: data <= 20'hfe686; 
        10'b0011110101: data <= 20'hfe6c5; 
        10'b0011110110: data <= 20'hfee5e; 
        10'b0011110111: data <= 20'hff079; 
        10'b0011111000: data <= 20'hff64f; 
        10'b0011111001: data <= 20'hff9e5; 
        10'b0011111010: data <= 20'hffb9e; 
        10'b0011111011: data <= 20'h000a6; 
        10'b0011111100: data <= 20'hfffaf; 
        10'b0011111101: data <= 20'hffe4b; 
        10'b0011111110: data <= 20'hfff05; 
        10'b0011111111: data <= 20'hffe0f; 
        10'b0100000000: data <= 20'h0000f; 
        10'b0100000001: data <= 20'hffe36; 
        10'b0100000010: data <= 20'hffd48; 
        10'b0100000011: data <= 20'hffe6d; 
        10'b0100000100: data <= 20'h001dd; 
        10'b0100000101: data <= 20'hffb14; 
        10'b0100000110: data <= 20'hff6b1; 
        10'b0100000111: data <= 20'hff8dd; 
        10'b0100001000: data <= 20'hffb67; 
        10'b0100001001: data <= 20'hff754; 
        10'b0100001010: data <= 20'hff80f; 
        10'b0100001011: data <= 20'hfeea0; 
        10'b0100001100: data <= 20'hfebc2; 
        10'b0100001101: data <= 20'hfe2ac; 
        10'b0100001110: data <= 20'hfe0b8; 
        10'b0100001111: data <= 20'hfe674; 
        10'b0100010000: data <= 20'hfeb0c; 
        10'b0100010001: data <= 20'hfef55; 
        10'b0100010010: data <= 20'hfecb2; 
        10'b0100010011: data <= 20'hff397; 
        10'b0100010100: data <= 20'hff689; 
        10'b0100010101: data <= 20'hff8fa; 
        10'b0100010110: data <= 20'hffd1c; 
        10'b0100010111: data <= 20'h00185; 
        10'b0100011000: data <= 20'hffe88; 
        10'b0100011001: data <= 20'h001eb; 
        10'b0100011010: data <= 20'h0014c; 
        10'b0100011011: data <= 20'hffdc0; 
        10'b0100011100: data <= 20'hffcba; 
        10'b0100011101: data <= 20'h000d5; 
        10'b0100011110: data <= 20'h002b3; 
        10'b0100011111: data <= 20'h00298; 
        10'b0100100000: data <= 20'h00980; 
        10'b0100100001: data <= 20'hfffce; 
        10'b0100100010: data <= 20'h001e4; 
        10'b0100100011: data <= 20'h000c9; 
        10'b0100100100: data <= 20'hffa41; 
        10'b0100100101: data <= 20'hffc18; 
        10'b0100100110: data <= 20'hff76d; 
        10'b0100100111: data <= 20'hfee04; 
        10'b0100101000: data <= 20'hfedb7; 
        10'b0100101001: data <= 20'hfea8f; 
        10'b0100101010: data <= 20'hfe9ad; 
        10'b0100101011: data <= 20'hfee2c; 
        10'b0100101100: data <= 20'hff3e6; 
        10'b0100101101: data <= 20'hff755; 
        10'b0100101110: data <= 20'hff498; 
        10'b0100101111: data <= 20'hffece; 
        10'b0100110000: data <= 20'hff895; 
        10'b0100110001: data <= 20'hffad8; 
        10'b0100110010: data <= 20'hffe78; 
        10'b0100110011: data <= 20'hfff42; 
        10'b0100110100: data <= 20'hffecf; 
        10'b0100110101: data <= 20'h000c7; 
        10'b0100110110: data <= 20'hffeb1; 
        10'b0100110111: data <= 20'hfffd0; 
        10'b0100111000: data <= 20'hffeb4; 
        10'b0100111001: data <= 20'h00057; 
        10'b0100111010: data <= 20'hfff4c; 
        10'b0100111011: data <= 20'h007f3; 
        10'b0100111100: data <= 20'h005b0; 
        10'b0100111101: data <= 20'h002bc; 
        10'b0100111110: data <= 20'h00370; 
        10'b0100111111: data <= 20'h0026f; 
        10'b0101000000: data <= 20'h00270; 
        10'b0101000001: data <= 20'h00064; 
        10'b0101000010: data <= 20'hffbdc; 
        10'b0101000011: data <= 20'hff1bd; 
        10'b0101000100: data <= 20'hff29f; 
        10'b0101000101: data <= 20'hff49d; 
        10'b0101000110: data <= 20'hff491; 
        10'b0101000111: data <= 20'hff719; 
        10'b0101001000: data <= 20'hffbd8; 
        10'b0101001001: data <= 20'h0019a; 
        10'b0101001010: data <= 20'h00575; 
        10'b0101001011: data <= 20'h0087d; 
        10'b0101001100: data <= 20'hffffb; 
        10'b0101001101: data <= 20'hffb7c; 
        10'b0101001110: data <= 20'hffe1d; 
        10'b0101001111: data <= 20'hfff4f; 
        10'b0101010000: data <= 20'hffecd; 
        10'b0101010001: data <= 20'hfff5c; 
        10'b0101010010: data <= 20'hffe0d; 
        10'b0101010011: data <= 20'hfff12; 
        10'b0101010100: data <= 20'h00122; 
        10'b0101010101: data <= 20'h003b8; 
        10'b0101010110: data <= 20'h005af; 
        10'b0101010111: data <= 20'h00774; 
        10'b0101011000: data <= 20'h00375; 
        10'b0101011001: data <= 20'h004d7; 
        10'b0101011010: data <= 20'h0036b; 
        10'b0101011011: data <= 20'h008fb; 
        10'b0101011100: data <= 20'h008a5; 
        10'b0101011101: data <= 20'h0062f; 
        10'b0101011110: data <= 20'hffab3; 
        10'b0101011111: data <= 20'hff66e; 
        10'b0101100000: data <= 20'hfff99; 
        10'b0101100001: data <= 20'hfff1e; 
        10'b0101100010: data <= 20'hff6a2; 
        10'b0101100011: data <= 20'hff706; 
        10'b0101100100: data <= 20'hffee3; 
        10'b0101100101: data <= 20'h00512; 
        10'b0101100110: data <= 20'h00c40; 
        10'b0101100111: data <= 20'h015bc; 
        10'b0101101000: data <= 20'h00bb1; 
        10'b0101101001: data <= 20'hffcaa; 
        10'b0101101010: data <= 20'hffc2c; 
        10'b0101101011: data <= 20'hffed8; 
        10'b0101101100: data <= 20'hffedd; 
        10'b0101101101: data <= 20'h00205; 
        10'b0101101110: data <= 20'h0018b; 
        10'b0101101111: data <= 20'hffdce; 
        10'b0101110000: data <= 20'hffd00; 
        10'b0101110001: data <= 20'h00136; 
        10'b0101110010: data <= 20'h0096f; 
        10'b0101110011: data <= 20'h00513; 
        10'b0101110100: data <= 20'h0045d; 
        10'b0101110101: data <= 20'h00228; 
        10'b0101110110: data <= 20'h00928; 
        10'b0101110111: data <= 20'h007a4; 
        10'b0101111000: data <= 20'h00702; 
        10'b0101111001: data <= 20'h0013d; 
        10'b0101111010: data <= 20'hffeb4; 
        10'b0101111011: data <= 20'hfffc7; 
        10'b0101111100: data <= 20'h000b6; 
        10'b0101111101: data <= 20'hffdf1; 
        10'b0101111110: data <= 20'hff7d8; 
        10'b0101111111: data <= 20'hffeed; 
        10'b0110000000: data <= 20'hffc14; 
        10'b0110000001: data <= 20'h00685; 
        10'b0110000010: data <= 20'h010f6; 
        10'b0110000011: data <= 20'h01adf; 
        10'b0110000100: data <= 20'h00e84; 
        10'b0110000101: data <= 20'hffed7; 
        10'b0110000110: data <= 20'h0000b; 
        10'b0110000111: data <= 20'h00151; 
        10'b0110001000: data <= 20'hfff09; 
        10'b0110001001: data <= 20'h00036; 
        10'b0110001010: data <= 20'h00186; 
        10'b0110001011: data <= 20'h00014; 
        10'b0110001100: data <= 20'hffcd3; 
        10'b0110001101: data <= 20'h00361; 
        10'b0110001110: data <= 20'h008a6; 
        10'b0110001111: data <= 20'h00774; 
        10'b0110010000: data <= 20'h00a43; 
        10'b0110010001: data <= 20'h0099c; 
        10'b0110010010: data <= 20'h00a67; 
        10'b0110010011: data <= 20'h00b43; 
        10'b0110010100: data <= 20'h003cb; 
        10'b0110010101: data <= 20'hffa82; 
        10'b0110010110: data <= 20'h0005d; 
        10'b0110010111: data <= 20'h00497; 
        10'b0110011000: data <= 20'h0022c; 
        10'b0110011001: data <= 20'hffc6e; 
        10'b0110011010: data <= 20'hffc88; 
        10'b0110011011: data <= 20'hfff80; 
        10'b0110011100: data <= 20'h0075c; 
        10'b0110011101: data <= 20'h00747; 
        10'b0110011110: data <= 20'h01334; 
        10'b0110011111: data <= 20'h01659; 
        10'b0110100000: data <= 20'h00ea7; 
        10'b0110100001: data <= 20'hfffcc; 
        10'b0110100010: data <= 20'hffbce; 
        10'b0110100011: data <= 20'hffdef; 
        10'b0110100100: data <= 20'h00192; 
        10'b0110100101: data <= 20'hfff34; 
        10'b0110100110: data <= 20'h0004e; 
        10'b0110100111: data <= 20'hffe45; 
        10'b0110101000: data <= 20'hff9f0; 
        10'b0110101001: data <= 20'hfff3c; 
        10'b0110101010: data <= 20'h00905; 
        10'b0110101011: data <= 20'h00bfd; 
        10'b0110101100: data <= 20'h007b8; 
        10'b0110101101: data <= 20'h00c1e; 
        10'b0110101110: data <= 20'h00f45; 
        10'b0110101111: data <= 20'h012a2; 
        10'b0110110000: data <= 20'h004de; 
        10'b0110110001: data <= 20'hffea6; 
        10'b0110110010: data <= 20'h00730; 
        10'b0110110011: data <= 20'h0069d; 
        10'b0110110100: data <= 20'h00106; 
        10'b0110110101: data <= 20'hffc9d; 
        10'b0110110110: data <= 20'h000af; 
        10'b0110110111: data <= 20'h003b6; 
        10'b0110111000: data <= 20'h0089c; 
        10'b0110111001: data <= 20'h00bd1; 
        10'b0110111010: data <= 20'h00adc; 
        10'b0110111011: data <= 20'h00d75; 
        10'b0110111100: data <= 20'h0072e; 
        10'b0110111101: data <= 20'hffc51; 
        10'b0110111110: data <= 20'hffdb6; 
        10'b0110111111: data <= 20'hffda8; 
        10'b0111000000: data <= 20'h0006b; 
        10'b0111000001: data <= 20'hffe4a; 
        10'b0111000010: data <= 20'hffe39; 
        10'b0111000011: data <= 20'hffe09; 
        10'b0111000100: data <= 20'hff7fd; 
        10'b0111000101: data <= 20'hffba7; 
        10'b0111000110: data <= 20'h00d5c; 
        10'b0111000111: data <= 20'h00da7; 
        10'b0111001000: data <= 20'h00908; 
        10'b0111001001: data <= 20'h00df0; 
        10'b0111001010: data <= 20'h017a3; 
        10'b0111001011: data <= 20'h01772; 
        10'b0111001100: data <= 20'h00726; 
        10'b0111001101: data <= 20'h00440; 
        10'b0111001110: data <= 20'h00a30; 
        10'b0111001111: data <= 20'h00560; 
        10'b0111010000: data <= 20'hffd30; 
        10'b0111010001: data <= 20'hffa6d; 
        10'b0111010010: data <= 20'h001ed; 
        10'b0111010011: data <= 20'h005f4; 
        10'b0111010100: data <= 20'h002c5; 
        10'b0111010101: data <= 20'h00015; 
        10'b0111010110: data <= 20'h00590; 
        10'b0111010111: data <= 20'h00355; 
        10'b0111011000: data <= 20'hffe62; 
        10'b0111011001: data <= 20'hffbab; 
        10'b0111011010: data <= 20'hffd58; 
        10'b0111011011: data <= 20'hfffa3; 
        10'b0111011100: data <= 20'h00065; 
        10'b0111011101: data <= 20'h00151; 
        10'b0111011110: data <= 20'h001d1; 
        10'b0111011111: data <= 20'hfffae; 
        10'b0111100000: data <= 20'hff492; 
        10'b0111100001: data <= 20'hffa06; 
        10'b0111100010: data <= 20'h00596; 
        10'b0111100011: data <= 20'h00a9e; 
        10'b0111100100: data <= 20'h00c14; 
        10'b0111100101: data <= 20'h00f3c; 
        10'b0111100110: data <= 20'h01a4b; 
        10'b0111100111: data <= 20'h01ab9; 
        10'b0111101000: data <= 20'h00dce; 
        10'b0111101001: data <= 20'h007c6; 
        10'b0111101010: data <= 20'h007df; 
        10'b0111101011: data <= 20'h004f8; 
        10'b0111101100: data <= 20'hfffff; 
        10'b0111101101: data <= 20'h00170; 
        10'b0111101110: data <= 20'h00af3; 
        10'b0111101111: data <= 20'h003c8; 
        10'b0111110000: data <= 20'h00191; 
        10'b0111110001: data <= 20'hffd35; 
        10'b0111110010: data <= 20'h00281; 
        10'b0111110011: data <= 20'hfff77; 
        10'b0111110100: data <= 20'hffce3; 
        10'b0111110101: data <= 20'hff9f1; 
        10'b0111110110: data <= 20'hfff22; 
        10'b0111110111: data <= 20'h000fd; 
        10'b0111111000: data <= 20'hfff1b; 
        10'b0111111001: data <= 20'hffec4; 
        10'b0111111010: data <= 20'hffff7; 
        10'b0111111011: data <= 20'hffcaa; 
        10'b0111111100: data <= 20'hff547; 
        10'b0111111101: data <= 20'hff588; 
        10'b0111111110: data <= 20'hffaee; 
        10'b0111111111: data <= 20'h0074d; 
        10'b1000000000: data <= 20'h00bb3; 
        10'b1000000001: data <= 20'h00aa2; 
        10'b1000000010: data <= 20'h0126a; 
        10'b1000000011: data <= 20'h016b6; 
        10'b1000000100: data <= 20'h01ac3; 
        10'b1000000101: data <= 20'h00c6e; 
        10'b1000000110: data <= 20'h0035d; 
        10'b1000000111: data <= 20'h006eb; 
        10'b1000001000: data <= 20'h00bf1; 
        10'b1000001001: data <= 20'h007bf; 
        10'b1000001010: data <= 20'h009a6; 
        10'b1000001011: data <= 20'h00514; 
        10'b1000001100: data <= 20'h000a7; 
        10'b1000001101: data <= 20'h001b2; 
        10'b1000001110: data <= 20'h001e0; 
        10'b1000001111: data <= 20'hffef1; 
        10'b1000010000: data <= 20'hffc2e; 
        10'b1000010001: data <= 20'hffd2f; 
        10'b1000010010: data <= 20'hffdd2; 
        10'b1000010011: data <= 20'hffdae; 
        10'b1000010100: data <= 20'h00093; 
        10'b1000010101: data <= 20'hffe61; 
        10'b1000010110: data <= 20'h00106; 
        10'b1000010111: data <= 20'hffbc4; 
        10'b1000011000: data <= 20'hff90e; 
        10'b1000011001: data <= 20'hff4dc; 
        10'b1000011010: data <= 20'hff759; 
        10'b1000011011: data <= 20'h0009d; 
        10'b1000011100: data <= 20'h00798; 
        10'b1000011101: data <= 20'h00bee; 
        10'b1000011110: data <= 20'h00fe3; 
        10'b1000011111: data <= 20'h01952; 
        10'b1000100000: data <= 20'h01c7d; 
        10'b1000100001: data <= 20'h00eb0; 
        10'b1000100010: data <= 20'h00d1f; 
        10'b1000100011: data <= 20'h00db7; 
        10'b1000100100: data <= 20'h009c4; 
        10'b1000100101: data <= 20'h00807; 
        10'b1000100110: data <= 20'h00c86; 
        10'b1000100111: data <= 20'h00887; 
        10'b1000101000: data <= 20'h00585; 
        10'b1000101001: data <= 20'h00130; 
        10'b1000101010: data <= 20'hffe01; 
        10'b1000101011: data <= 20'hffd89; 
        10'b1000101100: data <= 20'hffd6b; 
        10'b1000101101: data <= 20'hfff96; 
        10'b1000101110: data <= 20'hffec3; 
        10'b1000101111: data <= 20'h001d3; 
        10'b1000110000: data <= 20'hffee1; 
        10'b1000110001: data <= 20'hffe5f; 
        10'b1000110010: data <= 20'hfff6e; 
        10'b1000110011: data <= 20'hffe15; 
        10'b1000110100: data <= 20'hff71d; 
        10'b1000110101: data <= 20'hff560; 
        10'b1000110110: data <= 20'hff6cd; 
        10'b1000110111: data <= 20'hffc3e; 
        10'b1000111000: data <= 20'h00283; 
        10'b1000111001: data <= 20'h007fc; 
        10'b1000111010: data <= 20'h00d27; 
        10'b1000111011: data <= 20'h008c4; 
        10'b1000111100: data <= 20'h01142; 
        10'b1000111101: data <= 20'h014b1; 
        10'b1000111110: data <= 20'h01890; 
        10'b1000111111: data <= 20'h014e9; 
        10'b1001000000: data <= 20'h00b56; 
        10'b1001000001: data <= 20'h00740; 
        10'b1001000010: data <= 20'h00e14; 
        10'b1001000011: data <= 20'h009ed; 
        10'b1001000100: data <= 20'h006bc; 
        10'b1001000101: data <= 20'hffe9e; 
        10'b1001000110: data <= 20'hffac8; 
        10'b1001000111: data <= 20'h00057; 
        10'b1001001000: data <= 20'hffebd; 
        10'b1001001001: data <= 20'hfff5f; 
        10'b1001001010: data <= 20'hffe6b; 
        10'b1001001011: data <= 20'h00055; 
        10'b1001001100: data <= 20'hfffcc; 
        10'b1001001101: data <= 20'h00035; 
        10'b1001001110: data <= 20'h000aa; 
        10'b1001001111: data <= 20'hfff52; 
        10'b1001010000: data <= 20'hffca2; 
        10'b1001010001: data <= 20'hff8af; 
        10'b1001010010: data <= 20'hff393; 
        10'b1001010011: data <= 20'hffa60; 
        10'b1001010100: data <= 20'hffca1; 
        10'b1001010101: data <= 20'h00603; 
        10'b1001010110: data <= 20'h00aea; 
        10'b1001010111: data <= 20'h00f86; 
        10'b1001011000: data <= 20'h013f8; 
        10'b1001011001: data <= 20'h01447; 
        10'b1001011010: data <= 20'h01105; 
        10'b1001011011: data <= 20'h00eac; 
        10'b1001011100: data <= 20'h00928; 
        10'b1001011101: data <= 20'h00c86; 
        10'b1001011110: data <= 20'h00bac; 
        10'b1001011111: data <= 20'h00776; 
        10'b1001100000: data <= 20'h000fe; 
        10'b1001100001: data <= 20'hffc0c; 
        10'b1001100010: data <= 20'hffa76; 
        10'b1001100011: data <= 20'hffcc8; 
        10'b1001100100: data <= 20'h00030; 
        10'b1001100101: data <= 20'hffdea; 
        10'b1001100110: data <= 20'hfff8d; 
        10'b1001100111: data <= 20'hffed8; 
        10'b1001101000: data <= 20'hffed5; 
        10'b1001101001: data <= 20'hfffcd; 
        10'b1001101010: data <= 20'h001fe; 
        10'b1001101011: data <= 20'h0008a; 
        10'b1001101100: data <= 20'hffed3; 
        10'b1001101101: data <= 20'hff9a0; 
        10'b1001101110: data <= 20'hff86e; 
        10'b1001101111: data <= 20'hff5d8; 
        10'b1001110000: data <= 20'hff93a; 
        10'b1001110001: data <= 20'hffced; 
        10'b1001110010: data <= 20'hffd79; 
        10'b1001110011: data <= 20'h0013a; 
        10'b1001110100: data <= 20'h005d6; 
        10'b1001110101: data <= 20'h00287; 
        10'b1001110110: data <= 20'h00221; 
        10'b1001110111: data <= 20'h0064d; 
        10'b1001111000: data <= 20'h004b1; 
        10'b1001111001: data <= 20'h0000a; 
        10'b1001111010: data <= 20'hffe6e; 
        10'b1001111011: data <= 20'hff8f5; 
        10'b1001111100: data <= 20'hff939; 
        10'b1001111101: data <= 20'hffa5d; 
        10'b1001111110: data <= 20'hffabb; 
        10'b1001111111: data <= 20'hfff7e; 
        10'b1010000000: data <= 20'hfff14; 
        10'b1010000001: data <= 20'hffe09; 
        10'b1010000010: data <= 20'h00226; 
        10'b1010000011: data <= 20'h000d4; 
        10'b1010000100: data <= 20'h001ba; 
        10'b1010000101: data <= 20'hfff52; 
        10'b1010000110: data <= 20'hfff09; 
        10'b1010000111: data <= 20'h00033; 
        10'b1010001000: data <= 20'h0009b; 
        10'b1010001001: data <= 20'hffd5e; 
        10'b1010001010: data <= 20'hffbe1; 
        10'b1010001011: data <= 20'hff6f5; 
        10'b1010001100: data <= 20'hff491; 
        10'b1010001101: data <= 20'hfef8d; 
        10'b1010001110: data <= 20'hfefa2; 
        10'b1010001111: data <= 20'hfecec; 
        10'b1010010000: data <= 20'hff43e; 
        10'b1010010001: data <= 20'hff6bd; 
        10'b1010010010: data <= 20'hff8c7; 
        10'b1010010011: data <= 20'hff543; 
        10'b1010010100: data <= 20'hff1e3; 
        10'b1010010101: data <= 20'hfefff; 
        10'b1010010110: data <= 20'hff363; 
        10'b1010010111: data <= 20'hffa3f; 
        10'b1010011000: data <= 20'hffa25; 
        10'b1010011001: data <= 20'hffae0; 
        10'b1010011010: data <= 20'hffe2c; 
        10'b1010011011: data <= 20'h00041; 
        10'b1010011100: data <= 20'hffdde; 
        10'b1010011101: data <= 20'hffe3d; 
        10'b1010011110: data <= 20'hfff3f; 
        10'b1010011111: data <= 20'hfffc8; 
        10'b1010100000: data <= 20'h0013d; 
        10'b1010100001: data <= 20'h000ff; 
        10'b1010100010: data <= 20'h000ae; 
        10'b1010100011: data <= 20'hffdf9; 
        10'b1010100100: data <= 20'hffe63; 
        10'b1010100101: data <= 20'hfff3e; 
        10'b1010100110: data <= 20'hffe0e; 
        10'b1010100111: data <= 20'hffcd9; 
        10'b1010101000: data <= 20'hffd82; 
        10'b1010101001: data <= 20'hffc04; 
        10'b1010101010: data <= 20'hffa07; 
        10'b1010101011: data <= 20'hff871; 
        10'b1010101100: data <= 20'hff736; 
        10'b1010101101: data <= 20'hff766; 
        10'b1010101110: data <= 20'hff5f6; 
        10'b1010101111: data <= 20'hff5f8; 
        10'b1010110000: data <= 20'hff583; 
        10'b1010110001: data <= 20'hff7ff; 
        10'b1010110010: data <= 20'hffd39; 
        10'b1010110011: data <= 20'hffd6b; 
        10'b1010110100: data <= 20'hfff19; 
        10'b1010110101: data <= 20'hffe93; 
        10'b1010110110: data <= 20'h0010f; 
        10'b1010110111: data <= 20'hfff89; 
        10'b1010111000: data <= 20'hffde8; 
        10'b1010111001: data <= 20'hfff57; 
        10'b1010111010: data <= 20'hffe71; 
        10'b1010111011: data <= 20'hffe7b; 
        10'b1010111100: data <= 20'h001f4; 
        10'b1010111101: data <= 20'hffe2e; 
        10'b1010111110: data <= 20'h00089; 
        10'b1010111111: data <= 20'hfff12; 
        10'b1011000000: data <= 20'hffe93; 
        10'b1011000001: data <= 20'hfffbb; 
        10'b1011000010: data <= 20'h0014d; 
        10'b1011000011: data <= 20'hfffe6; 
        10'b1011000100: data <= 20'hffdc8; 
        10'b1011000101: data <= 20'h000ce; 
        10'b1011000110: data <= 20'hffdd6; 
        10'b1011000111: data <= 20'hfffab; 
        10'b1011001000: data <= 20'h0001c; 
        10'b1011001001: data <= 20'hffdb5; 
        10'b1011001010: data <= 20'hffebd; 
        10'b1011001011: data <= 20'hfff3a; 
        10'b1011001100: data <= 20'hfffcb; 
        10'b1011001101: data <= 20'hffe01; 
        10'b1011001110: data <= 20'hffed5; 
        10'b1011001111: data <= 20'hffdcb; 
        10'b1011010000: data <= 20'hffe43; 
        10'b1011010001: data <= 20'h00046; 
        10'b1011010010: data <= 20'hfff2a; 
        10'b1011010011: data <= 20'h00196; 
        10'b1011010100: data <= 20'h0023f; 
        10'b1011010101: data <= 20'h001fc; 
        10'b1011010110: data <= 20'h00017; 
        10'b1011010111: data <= 20'h0017d; 
        10'b1011011000: data <= 20'h0021b; 
        10'b1011011001: data <= 20'hfffe7; 
        10'b1011011010: data <= 20'h00063; 
        10'b1011011011: data <= 20'hfff99; 
        10'b1011011100: data <= 20'hffed0; 
        10'b1011011101: data <= 20'h001c7; 
        10'b1011011110: data <= 20'h00156; 
        10'b1011011111: data <= 20'hffed9; 
        10'b1011100000: data <= 20'hfff50; 
        10'b1011100001: data <= 20'h00101; 
        10'b1011100010: data <= 20'hfff2b; 
        10'b1011100011: data <= 20'h00071; 
        10'b1011100100: data <= 20'hfff20; 
        10'b1011100101: data <= 20'h0014f; 
        10'b1011100110: data <= 20'h00160; 
        10'b1011100111: data <= 20'hffe38; 
        10'b1011101000: data <= 20'hffea5; 
        10'b1011101001: data <= 20'h001cd; 
        10'b1011101010: data <= 20'h0016a; 
        10'b1011101011: data <= 20'hfff4f; 
        10'b1011101100: data <= 20'h00144; 
        10'b1011101101: data <= 20'hfff85; 
        10'b1011101110: data <= 20'hfff7f; 
        10'b1011101111: data <= 20'h000ca; 
        10'b1011110000: data <= 20'h000e7; 
        10'b1011110001: data <= 20'hfff8f; 
        10'b1011110010: data <= 20'hffef1; 
        10'b1011110011: data <= 20'hfff65; 
        10'b1011110100: data <= 20'h00209; 
        10'b1011110101: data <= 20'hfffe6; 
        10'b1011110110: data <= 20'h00126; 
        10'b1011110111: data <= 20'hffed5; 
        10'b1011111000: data <= 20'h000b6; 
        10'b1011111001: data <= 20'hffff1; 
        10'b1011111010: data <= 20'h001ea; 
        10'b1011111011: data <= 20'h00046; 
        10'b1011111100: data <= 20'hfffbf; 
        10'b1011111101: data <= 20'hffdbf; 
        10'b1011111110: data <= 20'hffe7a; 
        10'b1011111111: data <= 20'h000b2; 
        10'b1100000000: data <= 20'hffdf7; 
        10'b1100000001: data <= 20'hffe4c; 
        10'b1100000010: data <= 20'hffeb6; 
        10'b1100000011: data <= 20'hffdec; 
        10'b1100000100: data <= 20'hffe97; 
        10'b1100000101: data <= 20'hfff4e; 
        10'b1100000110: data <= 20'hffe23; 
        10'b1100000111: data <= 20'hffe98; 
        10'b1100001000: data <= 20'hffec9; 
        10'b1100001001: data <= 20'hfff02; 
        10'b1100001010: data <= 20'h001e2; 
        10'b1100001011: data <= 20'hffe29; 
        10'b1100001100: data <= 20'hffecd; 
        10'b1100001101: data <= 20'hffe38; 
        10'b1100001110: data <= 20'hffec0; 
        10'b1100001111: data <= 20'h00059; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 15) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 21'h1ffe94; 
        10'b0000000001: data <= 21'h0002e7; 
        10'b0000000010: data <= 21'h1ffcb8; 
        10'b0000000011: data <= 21'h1fffbf; 
        10'b0000000100: data <= 21'h1fffe4; 
        10'b0000000101: data <= 21'h1fff8e; 
        10'b0000000110: data <= 21'h000187; 
        10'b0000000111: data <= 21'h00049c; 
        10'b0000001000: data <= 21'h1ffcf9; 
        10'b0000001001: data <= 21'h1ffdfe; 
        10'b0000001010: data <= 21'h1ffe1f; 
        10'b0000001011: data <= 21'h1ffd1c; 
        10'b0000001100: data <= 21'h00017e; 
        10'b0000001101: data <= 21'h000436; 
        10'b0000001110: data <= 21'h00025e; 
        10'b0000001111: data <= 21'h1ffc26; 
        10'b0000010000: data <= 21'h1fff79; 
        10'b0000010001: data <= 21'h00049b; 
        10'b0000010010: data <= 21'h0000c8; 
        10'b0000010011: data <= 21'h1fff98; 
        10'b0000010100: data <= 21'h1ffc74; 
        10'b0000010101: data <= 21'h1ffda2; 
        10'b0000010110: data <= 21'h000116; 
        10'b0000010111: data <= 21'h00040a; 
        10'b0000011000: data <= 21'h00022e; 
        10'b0000011001: data <= 21'h0002a8; 
        10'b0000011010: data <= 21'h1ffc66; 
        10'b0000011011: data <= 21'h1ffc8c; 
        10'b0000011100: data <= 21'h0002f7; 
        10'b0000011101: data <= 21'h000259; 
        10'b0000011110: data <= 21'h0002fc; 
        10'b0000011111: data <= 21'h1fff3d; 
        10'b0000100000: data <= 21'h1ffbf6; 
        10'b0000100001: data <= 21'h1ffd97; 
        10'b0000100010: data <= 21'h000210; 
        10'b0000100011: data <= 21'h0006b5; 
        10'b0000100100: data <= 21'h00048c; 
        10'b0000100101: data <= 21'h00015e; 
        10'b0000100110: data <= 21'h000581; 
        10'b0000100111: data <= 21'h0005e0; 
        10'b0000101000: data <= 21'h000642; 
        10'b0000101001: data <= 21'h0005e6; 
        10'b0000101010: data <= 21'h0003b7; 
        10'b0000101011: data <= 21'h0003f9; 
        10'b0000101100: data <= 21'h1ffbc2; 
        10'b0000101101: data <= 21'h0003c8; 
        10'b0000101110: data <= 21'h000521; 
        10'b0000101111: data <= 21'h0002eb; 
        10'b0000110000: data <= 21'h1fff2d; 
        10'b0000110001: data <= 21'h1ffd65; 
        10'b0000110010: data <= 21'h000571; 
        10'b0000110011: data <= 21'h00041c; 
        10'b0000110100: data <= 21'h1ffe4f; 
        10'b0000110101: data <= 21'h000496; 
        10'b0000110110: data <= 21'h1fff36; 
        10'b0000110111: data <= 21'h000365; 
        10'b0000111000: data <= 21'h1ffd53; 
        10'b0000111001: data <= 21'h1ffcc8; 
        10'b0000111010: data <= 21'h1ffbf4; 
        10'b0000111011: data <= 21'h1fff9b; 
        10'b0000111100: data <= 21'h000248; 
        10'b0000111101: data <= 21'h000168; 
        10'b0000111110: data <= 21'h000255; 
        10'b0000111111: data <= 21'h000690; 
        10'b0001000000: data <= 21'h0004aa; 
        10'b0001000001: data <= 21'h0009f1; 
        10'b0001000010: data <= 21'h000c82; 
        10'b0001000011: data <= 21'h000e22; 
        10'b0001000100: data <= 21'h000e2a; 
        10'b0001000101: data <= 21'h000ee2; 
        10'b0001000110: data <= 21'h00078b; 
        10'b0001000111: data <= 21'h000559; 
        10'b0001001000: data <= 21'h000c6c; 
        10'b0001001001: data <= 21'h00057b; 
        10'b0001001010: data <= 21'h000555; 
        10'b0001001011: data <= 21'h0005d7; 
        10'b0001001100: data <= 21'h0005b6; 
        10'b0001001101: data <= 21'h0002e4; 
        10'b0001001110: data <= 21'h0003ce; 
        10'b0001001111: data <= 21'h0000b6; 
        10'b0001010000: data <= 21'h000218; 
        10'b0001010001: data <= 21'h1ffece; 
        10'b0001010010: data <= 21'h1ffbca; 
        10'b0001010011: data <= 21'h00014a; 
        10'b0001010100: data <= 21'h1ffc6d; 
        10'b0001010101: data <= 21'h00006c; 
        10'b0001010110: data <= 21'h00035e; 
        10'b0001010111: data <= 21'h0001f2; 
        10'b0001011000: data <= 21'h00046b; 
        10'b0001011001: data <= 21'h1ffc28; 
        10'b0001011010: data <= 21'h0004cb; 
        10'b0001011011: data <= 21'h000541; 
        10'b0001011100: data <= 21'h000641; 
        10'b0001011101: data <= 21'h000cad; 
        10'b0001011110: data <= 21'h000b3b; 
        10'b0001011111: data <= 21'h000e10; 
        10'b0001100000: data <= 21'h000db8; 
        10'b0001100001: data <= 21'h000d35; 
        10'b0001100010: data <= 21'h00136e; 
        10'b0001100011: data <= 21'h001254; 
        10'b0001100100: data <= 21'h000b65; 
        10'b0001100101: data <= 21'h000e62; 
        10'b0001100110: data <= 21'h00171c; 
        10'b0001100111: data <= 21'h00170c; 
        10'b0001101000: data <= 21'h001895; 
        10'b0001101001: data <= 21'h0015c7; 
        10'b0001101010: data <= 21'h00160d; 
        10'b0001101011: data <= 21'h000ccf; 
        10'b0001101100: data <= 21'h000b5e; 
        10'b0001101101: data <= 21'h0002c7; 
        10'b0001101110: data <= 21'h1ffe0c; 
        10'b0001101111: data <= 21'h000283; 
        10'b0001110000: data <= 21'h0000aa; 
        10'b0001110001: data <= 21'h1fff29; 
        10'b0001110010: data <= 21'h1fffb4; 
        10'b0001110011: data <= 21'h0003e8; 
        10'b0001110100: data <= 21'h00035d; 
        10'b0001110101: data <= 21'h00013a; 
        10'b0001110110: data <= 21'h00013f; 
        10'b0001110111: data <= 21'h0007da; 
        10'b0001111000: data <= 21'h1fff20; 
        10'b0001111001: data <= 21'h1ffe5c; 
        10'b0001111010: data <= 21'h000798; 
        10'b0001111011: data <= 21'h0002dc; 
        10'b0001111100: data <= 21'h000386; 
        10'b0001111101: data <= 21'h000146; 
        10'b0001111110: data <= 21'h0002fe; 
        10'b0001111111: data <= 21'h00047f; 
        10'b0010000000: data <= 21'h000f68; 
        10'b0010000001: data <= 21'h000f41; 
        10'b0010000010: data <= 21'h0017e3; 
        10'b0010000011: data <= 21'h001849; 
        10'b0010000100: data <= 21'h001ea5; 
        10'b0010000101: data <= 21'h0021ff; 
        10'b0010000110: data <= 21'h001d3f; 
        10'b0010000111: data <= 21'h0013a4; 
        10'b0010001000: data <= 21'h0002c9; 
        10'b0010001001: data <= 21'h000537; 
        10'b0010001010: data <= 21'h0000b9; 
        10'b0010001011: data <= 21'h1fffff; 
        10'b0010001100: data <= 21'h0000c9; 
        10'b0010001101: data <= 21'h000260; 
        10'b0010001110: data <= 21'h00015b; 
        10'b0010001111: data <= 21'h1ffe31; 
        10'b0010010000: data <= 21'h1ffcc1; 
        10'b0010010001: data <= 21'h1fffa5; 
        10'b0010010010: data <= 21'h1ffd48; 
        10'b0010010011: data <= 21'h1ffa9e; 
        10'b0010010100: data <= 21'h000408; 
        10'b0010010101: data <= 21'h1fface; 
        10'b0010010110: data <= 21'h0001e0; 
        10'b0010010111: data <= 21'h1fee29; 
        10'b0010011000: data <= 21'h1ff68e; 
        10'b0010011001: data <= 21'h1ff97a; 
        10'b0010011010: data <= 21'h1ffd9a; 
        10'b0010011011: data <= 21'h1ff793; 
        10'b0010011100: data <= 21'h1ff793; 
        10'b0010011101: data <= 21'h00019f; 
        10'b0010011110: data <= 21'h000b76; 
        10'b0010011111: data <= 21'h00157c; 
        10'b0010100000: data <= 21'h0012a4; 
        10'b0010100001: data <= 21'h0010aa; 
        10'b0010100010: data <= 21'h000d25; 
        10'b0010100011: data <= 21'h000905; 
        10'b0010100100: data <= 21'h1ffef4; 
        10'b0010100101: data <= 21'h000074; 
        10'b0010100110: data <= 21'h1ffb78; 
        10'b0010100111: data <= 21'h000448; 
        10'b0010101000: data <= 21'h1fff6a; 
        10'b0010101001: data <= 21'h0003da; 
        10'b0010101010: data <= 21'h000398; 
        10'b0010101011: data <= 21'h1ffb5c; 
        10'b0010101100: data <= 21'h0001a5; 
        10'b0010101101: data <= 21'h1fff44; 
        10'b0010101110: data <= 21'h00017c; 
        10'b0010101111: data <= 21'h00001d; 
        10'b0010110000: data <= 21'h1ff95f; 
        10'b0010110001: data <= 21'h1ff7ec; 
        10'b0010110010: data <= 21'h1feb74; 
        10'b0010110011: data <= 21'h1fe524; 
        10'b0010110100: data <= 21'h1ff064; 
        10'b0010110101: data <= 21'h1fe160; 
        10'b0010110110: data <= 21'h1ff27d; 
        10'b0010110111: data <= 21'h1ff614; 
        10'b0010111000: data <= 21'h1ff1df; 
        10'b0010111001: data <= 21'h1ff384; 
        10'b0010111010: data <= 21'h1ffc88; 
        10'b0010111011: data <= 21'h1ff7a0; 
        10'b0010111100: data <= 21'h1ff26d; 
        10'b0010111101: data <= 21'h1ff310; 
        10'b0010111110: data <= 21'h1febe2; 
        10'b0010111111: data <= 21'h1ff2e1; 
        10'b0011000000: data <= 21'h1ff51d; 
        10'b0011000001: data <= 21'h1ff486; 
        10'b0011000010: data <= 21'h1ffe4a; 
        10'b0011000011: data <= 21'h0003bd; 
        10'b0011000100: data <= 21'h00017c; 
        10'b0011000101: data <= 21'h000239; 
        10'b0011000110: data <= 21'h000022; 
        10'b0011000111: data <= 21'h1fff44; 
        10'b0011001000: data <= 21'h000040; 
        10'b0011001001: data <= 21'h1ffc05; 
        10'b0011001010: data <= 21'h1ff7ee; 
        10'b0011001011: data <= 21'h1ffeb4; 
        10'b0011001100: data <= 21'h1ff48c; 
        10'b0011001101: data <= 21'h1ff1c7; 
        10'b0011001110: data <= 21'h1feb4c; 
        10'b0011001111: data <= 21'h1fefba; 
        10'b0011010000: data <= 21'h1fe2c3; 
        10'b0011010001: data <= 21'h1fdf3b; 
        10'b0011010010: data <= 21'h1feed1; 
        10'b0011010011: data <= 21'h1fefb3; 
        10'b0011010100: data <= 21'h1fe674; 
        10'b0011010101: data <= 21'h1fe7d1; 
        10'b0011010110: data <= 21'h1fe203; 
        10'b0011010111: data <= 21'h1fd751; 
        10'b0011011000: data <= 21'h1fd67b; 
        10'b0011011001: data <= 21'h1fdd47; 
        10'b0011011010: data <= 21'h1fdbad; 
        10'b0011011011: data <= 21'h1fe350; 
        10'b0011011100: data <= 21'h1ff509; 
        10'b0011011101: data <= 21'h1ff614; 
        10'b0011011110: data <= 21'h1ffc16; 
        10'b0011011111: data <= 21'h1ffd03; 
        10'b0011100000: data <= 21'h1ffe8f; 
        10'b0011100001: data <= 21'h1ffec7; 
        10'b0011100010: data <= 21'h000463; 
        10'b0011100011: data <= 21'h1ffa64; 
        10'b0011100100: data <= 21'h1ffb55; 
        10'b0011100101: data <= 21'h1ff9ca; 
        10'b0011100110: data <= 21'h1ff068; 
        10'b0011100111: data <= 21'h1ffc94; 
        10'b0011101000: data <= 21'h1ffa3e; 
        10'b0011101001: data <= 21'h1fefb1; 
        10'b0011101010: data <= 21'h1fecf5; 
        10'b0011101011: data <= 21'h1fea2c; 
        10'b0011101100: data <= 21'h1fe5b9; 
        10'b0011101101: data <= 21'h1fe187; 
        10'b0011101110: data <= 21'h1fe24f; 
        10'b0011101111: data <= 21'h1fe047; 
        10'b0011110000: data <= 21'h1fda64; 
        10'b0011110001: data <= 21'h1fd4ad; 
        10'b0011110010: data <= 21'h1fc2c7; 
        10'b0011110011: data <= 21'h1fc704; 
        10'b0011110100: data <= 21'h1fcd0c; 
        10'b0011110101: data <= 21'h1fcd8b; 
        10'b0011110110: data <= 21'h1fdcbd; 
        10'b0011110111: data <= 21'h1fe0f2; 
        10'b0011111000: data <= 21'h1fec9d; 
        10'b0011111001: data <= 21'h1ff3c9; 
        10'b0011111010: data <= 21'h1ff73c; 
        10'b0011111011: data <= 21'h00014c; 
        10'b0011111100: data <= 21'h1fff5e; 
        10'b0011111101: data <= 21'h1ffc96; 
        10'b0011111110: data <= 21'h1ffe0b; 
        10'b0011111111: data <= 21'h1ffc1d; 
        10'b0100000000: data <= 21'h00001e; 
        10'b0100000001: data <= 21'h1ffc6c; 
        10'b0100000010: data <= 21'h1ffa8f; 
        10'b0100000011: data <= 21'h1ffcda; 
        10'b0100000100: data <= 21'h0003ba; 
        10'b0100000101: data <= 21'h1ff628; 
        10'b0100000110: data <= 21'h1fed63; 
        10'b0100000111: data <= 21'h1ff1b9; 
        10'b0100001000: data <= 21'h1ff6ce; 
        10'b0100001001: data <= 21'h1feea9; 
        10'b0100001010: data <= 21'h1ff01e; 
        10'b0100001011: data <= 21'h1fdd40; 
        10'b0100001100: data <= 21'h1fd783; 
        10'b0100001101: data <= 21'h1fc559; 
        10'b0100001110: data <= 21'h1fc170; 
        10'b0100001111: data <= 21'h1fcce8; 
        10'b0100010000: data <= 21'h1fd617; 
        10'b0100010001: data <= 21'h1fdeaa; 
        10'b0100010010: data <= 21'h1fd963; 
        10'b0100010011: data <= 21'h1fe72f; 
        10'b0100010100: data <= 21'h1fed11; 
        10'b0100010101: data <= 21'h1ff1f3; 
        10'b0100010110: data <= 21'h1ffa38; 
        10'b0100010111: data <= 21'h00030a; 
        10'b0100011000: data <= 21'h1ffd0f; 
        10'b0100011001: data <= 21'h0003d6; 
        10'b0100011010: data <= 21'h000299; 
        10'b0100011011: data <= 21'h1ffb80; 
        10'b0100011100: data <= 21'h1ff973; 
        10'b0100011101: data <= 21'h0001aa; 
        10'b0100011110: data <= 21'h000566; 
        10'b0100011111: data <= 21'h000530; 
        10'b0100100000: data <= 21'h001300; 
        10'b0100100001: data <= 21'h1fff9b; 
        10'b0100100010: data <= 21'h0003c7; 
        10'b0100100011: data <= 21'h000193; 
        10'b0100100100: data <= 21'h1ff482; 
        10'b0100100101: data <= 21'h1ff830; 
        10'b0100100110: data <= 21'h1feedb; 
        10'b0100100111: data <= 21'h1fdc08; 
        10'b0100101000: data <= 21'h1fdb6d; 
        10'b0100101001: data <= 21'h1fd51d; 
        10'b0100101010: data <= 21'h1fd359; 
        10'b0100101011: data <= 21'h1fdc59; 
        10'b0100101100: data <= 21'h1fe7cb; 
        10'b0100101101: data <= 21'h1feeaa; 
        10'b0100101110: data <= 21'h1fe930; 
        10'b0100101111: data <= 21'h1ffd9d; 
        10'b0100110000: data <= 21'h1ff12a; 
        10'b0100110001: data <= 21'h1ff5b0; 
        10'b0100110010: data <= 21'h1ffcf0; 
        10'b0100110011: data <= 21'h1ffe85; 
        10'b0100110100: data <= 21'h1ffd9d; 
        10'b0100110101: data <= 21'h00018f; 
        10'b0100110110: data <= 21'h1ffd62; 
        10'b0100110111: data <= 21'h1fffa0; 
        10'b0100111000: data <= 21'h1ffd67; 
        10'b0100111001: data <= 21'h0000ad; 
        10'b0100111010: data <= 21'h1ffe97; 
        10'b0100111011: data <= 21'h000fe5; 
        10'b0100111100: data <= 21'h000b5f; 
        10'b0100111101: data <= 21'h000578; 
        10'b0100111110: data <= 21'h0006e0; 
        10'b0100111111: data <= 21'h0004dd; 
        10'b0101000000: data <= 21'h0004e0; 
        10'b0101000001: data <= 21'h0000c8; 
        10'b0101000010: data <= 21'h1ff7b7; 
        10'b0101000011: data <= 21'h1fe379; 
        10'b0101000100: data <= 21'h1fe53f; 
        10'b0101000101: data <= 21'h1fe93b; 
        10'b0101000110: data <= 21'h1fe922; 
        10'b0101000111: data <= 21'h1fee33; 
        10'b0101001000: data <= 21'h1ff7b0; 
        10'b0101001001: data <= 21'h000334; 
        10'b0101001010: data <= 21'h000ae9; 
        10'b0101001011: data <= 21'h0010fa; 
        10'b0101001100: data <= 21'h1ffff5; 
        10'b0101001101: data <= 21'h1ff6f8; 
        10'b0101001110: data <= 21'h1ffc3b; 
        10'b0101001111: data <= 21'h1ffe9f; 
        10'b0101010000: data <= 21'h1ffd9a; 
        10'b0101010001: data <= 21'h1ffeb8; 
        10'b0101010010: data <= 21'h1ffc1b; 
        10'b0101010011: data <= 21'h1ffe23; 
        10'b0101010100: data <= 21'h000245; 
        10'b0101010101: data <= 21'h000771; 
        10'b0101010110: data <= 21'h000b5e; 
        10'b0101010111: data <= 21'h000ee8; 
        10'b0101011000: data <= 21'h0006e9; 
        10'b0101011001: data <= 21'h0009af; 
        10'b0101011010: data <= 21'h0006d6; 
        10'b0101011011: data <= 21'h0011f7; 
        10'b0101011100: data <= 21'h001149; 
        10'b0101011101: data <= 21'h000c5e; 
        10'b0101011110: data <= 21'h1ff566; 
        10'b0101011111: data <= 21'h1fecdc; 
        10'b0101100000: data <= 21'h1fff32; 
        10'b0101100001: data <= 21'h1ffe3c; 
        10'b0101100010: data <= 21'h1fed44; 
        10'b0101100011: data <= 21'h1fee0c; 
        10'b0101100100: data <= 21'h1ffdc5; 
        10'b0101100101: data <= 21'h000a24; 
        10'b0101100110: data <= 21'h001880; 
        10'b0101100111: data <= 21'h002b78; 
        10'b0101101000: data <= 21'h001761; 
        10'b0101101001: data <= 21'h1ff955; 
        10'b0101101010: data <= 21'h1ff858; 
        10'b0101101011: data <= 21'h1ffdb0; 
        10'b0101101100: data <= 21'h1ffdb9; 
        10'b0101101101: data <= 21'h00040a; 
        10'b0101101110: data <= 21'h000316; 
        10'b0101101111: data <= 21'h1ffb9c; 
        10'b0101110000: data <= 21'h1ff9ff; 
        10'b0101110001: data <= 21'h00026b; 
        10'b0101110010: data <= 21'h0012dd; 
        10'b0101110011: data <= 21'h000a27; 
        10'b0101110100: data <= 21'h0008b9; 
        10'b0101110101: data <= 21'h000450; 
        10'b0101110110: data <= 21'h001250; 
        10'b0101110111: data <= 21'h000f48; 
        10'b0101111000: data <= 21'h000e05; 
        10'b0101111001: data <= 21'h00027a; 
        10'b0101111010: data <= 21'h1ffd68; 
        10'b0101111011: data <= 21'h1fff8e; 
        10'b0101111100: data <= 21'h00016b; 
        10'b0101111101: data <= 21'h1ffbe1; 
        10'b0101111110: data <= 21'h1fefb1; 
        10'b0101111111: data <= 21'h1ffddb; 
        10'b0110000000: data <= 21'h1ff828; 
        10'b0110000001: data <= 21'h000d0a; 
        10'b0110000010: data <= 21'h0021ec; 
        10'b0110000011: data <= 21'h0035be; 
        10'b0110000100: data <= 21'h001d08; 
        10'b0110000101: data <= 21'h1ffdaf; 
        10'b0110000110: data <= 21'h000017; 
        10'b0110000111: data <= 21'h0002a3; 
        10'b0110001000: data <= 21'h1ffe12; 
        10'b0110001001: data <= 21'h00006d; 
        10'b0110001010: data <= 21'h00030c; 
        10'b0110001011: data <= 21'h000029; 
        10'b0110001100: data <= 21'h1ff9a7; 
        10'b0110001101: data <= 21'h0006c2; 
        10'b0110001110: data <= 21'h00114d; 
        10'b0110001111: data <= 21'h000ee9; 
        10'b0110010000: data <= 21'h001486; 
        10'b0110010001: data <= 21'h001339; 
        10'b0110010010: data <= 21'h0014ce; 
        10'b0110010011: data <= 21'h001686; 
        10'b0110010100: data <= 21'h000796; 
        10'b0110010101: data <= 21'h1ff503; 
        10'b0110010110: data <= 21'h0000bb; 
        10'b0110010111: data <= 21'h00092e; 
        10'b0110011000: data <= 21'h000458; 
        10'b0110011001: data <= 21'h1ff8db; 
        10'b0110011010: data <= 21'h1ff90f; 
        10'b0110011011: data <= 21'h1fff01; 
        10'b0110011100: data <= 21'h000eb8; 
        10'b0110011101: data <= 21'h000e8d; 
        10'b0110011110: data <= 21'h002669; 
        10'b0110011111: data <= 21'h002cb2; 
        10'b0110100000: data <= 21'h001d4e; 
        10'b0110100001: data <= 21'h1fff97; 
        10'b0110100010: data <= 21'h1ff79d; 
        10'b0110100011: data <= 21'h1ffbdf; 
        10'b0110100100: data <= 21'h000323; 
        10'b0110100101: data <= 21'h1ffe68; 
        10'b0110100110: data <= 21'h00009d; 
        10'b0110100111: data <= 21'h1ffc8a; 
        10'b0110101000: data <= 21'h1ff3e0; 
        10'b0110101001: data <= 21'h1ffe79; 
        10'b0110101010: data <= 21'h00120a; 
        10'b0110101011: data <= 21'h0017fa; 
        10'b0110101100: data <= 21'h000f70; 
        10'b0110101101: data <= 21'h00183c; 
        10'b0110101110: data <= 21'h001e8b; 
        10'b0110101111: data <= 21'h002544; 
        10'b0110110000: data <= 21'h0009bc; 
        10'b0110110001: data <= 21'h1ffd4c; 
        10'b0110110010: data <= 21'h000e61; 
        10'b0110110011: data <= 21'h000d3a; 
        10'b0110110100: data <= 21'h00020c; 
        10'b0110110101: data <= 21'h1ff939; 
        10'b0110110110: data <= 21'h00015e; 
        10'b0110110111: data <= 21'h00076c; 
        10'b0110111000: data <= 21'h001138; 
        10'b0110111001: data <= 21'h0017a3; 
        10'b0110111010: data <= 21'h0015b8; 
        10'b0110111011: data <= 21'h001ae9; 
        10'b0110111100: data <= 21'h000e5c; 
        10'b0110111101: data <= 21'h1ff8a3; 
        10'b0110111110: data <= 21'h1ffb6b; 
        10'b0110111111: data <= 21'h1ffb50; 
        10'b0111000000: data <= 21'h0000d6; 
        10'b0111000001: data <= 21'h1ffc94; 
        10'b0111000010: data <= 21'h1ffc73; 
        10'b0111000011: data <= 21'h1ffc13; 
        10'b0111000100: data <= 21'h1feff9; 
        10'b0111000101: data <= 21'h1ff74e; 
        10'b0111000110: data <= 21'h001ab9; 
        10'b0111000111: data <= 21'h001b4d; 
        10'b0111001000: data <= 21'h001211; 
        10'b0111001001: data <= 21'h001bdf; 
        10'b0111001010: data <= 21'h002f46; 
        10'b0111001011: data <= 21'h002ee3; 
        10'b0111001100: data <= 21'h000e4d; 
        10'b0111001101: data <= 21'h000880; 
        10'b0111001110: data <= 21'h001461; 
        10'b0111001111: data <= 21'h000ac0; 
        10'b0111010000: data <= 21'h1ffa60; 
        10'b0111010001: data <= 21'h1ff4db; 
        10'b0111010010: data <= 21'h0003db; 
        10'b0111010011: data <= 21'h000be9; 
        10'b0111010100: data <= 21'h00058a; 
        10'b0111010101: data <= 21'h00002a; 
        10'b0111010110: data <= 21'h000b20; 
        10'b0111010111: data <= 21'h0006aa; 
        10'b0111011000: data <= 21'h1ffcc3; 
        10'b0111011001: data <= 21'h1ff756; 
        10'b0111011010: data <= 21'h1ffab0; 
        10'b0111011011: data <= 21'h1fff46; 
        10'b0111011100: data <= 21'h0000c9; 
        10'b0111011101: data <= 21'h0002a2; 
        10'b0111011110: data <= 21'h0003a1; 
        10'b0111011111: data <= 21'h1fff5d; 
        10'b0111100000: data <= 21'h1fe924; 
        10'b0111100001: data <= 21'h1ff40b; 
        10'b0111100010: data <= 21'h000b2c; 
        10'b0111100011: data <= 21'h00153b; 
        10'b0111100100: data <= 21'h001829; 
        10'b0111100101: data <= 21'h001e79; 
        10'b0111100110: data <= 21'h003497; 
        10'b0111100111: data <= 21'h003571; 
        10'b0111101000: data <= 21'h001b9d; 
        10'b0111101001: data <= 21'h000f8d; 
        10'b0111101010: data <= 21'h000fbe; 
        10'b0111101011: data <= 21'h0009f0; 
        10'b0111101100: data <= 21'h1ffffe; 
        10'b0111101101: data <= 21'h0002df; 
        10'b0111101110: data <= 21'h0015e7; 
        10'b0111101111: data <= 21'h000790; 
        10'b0111110000: data <= 21'h000323; 
        10'b0111110001: data <= 21'h1ffa6a; 
        10'b0111110010: data <= 21'h000502; 
        10'b0111110011: data <= 21'h1ffeef; 
        10'b0111110100: data <= 21'h1ff9c7; 
        10'b0111110101: data <= 21'h1ff3e1; 
        10'b0111110110: data <= 21'h1ffe43; 
        10'b0111110111: data <= 21'h0001fa; 
        10'b0111111000: data <= 21'h1ffe36; 
        10'b0111111001: data <= 21'h1ffd87; 
        10'b0111111010: data <= 21'h1fffee; 
        10'b0111111011: data <= 21'h1ff954; 
        10'b0111111100: data <= 21'h1fea8e; 
        10'b0111111101: data <= 21'h1feb11; 
        10'b0111111110: data <= 21'h1ff5dd; 
        10'b0111111111: data <= 21'h000e9a; 
        10'b1000000000: data <= 21'h001766; 
        10'b1000000001: data <= 21'h001545; 
        10'b1000000010: data <= 21'h0024d4; 
        10'b1000000011: data <= 21'h002d6d; 
        10'b1000000100: data <= 21'h003587; 
        10'b1000000101: data <= 21'h0018dd; 
        10'b1000000110: data <= 21'h0006ba; 
        10'b1000000111: data <= 21'h000dd6; 
        10'b1000001000: data <= 21'h0017e1; 
        10'b1000001001: data <= 21'h000f7e; 
        10'b1000001010: data <= 21'h00134b; 
        10'b1000001011: data <= 21'h000a28; 
        10'b1000001100: data <= 21'h00014f; 
        10'b1000001101: data <= 21'h000363; 
        10'b1000001110: data <= 21'h0003bf; 
        10'b1000001111: data <= 21'h1ffde1; 
        10'b1000010000: data <= 21'h1ff85d; 
        10'b1000010001: data <= 21'h1ffa5d; 
        10'b1000010010: data <= 21'h1ffba3; 
        10'b1000010011: data <= 21'h1ffb5c; 
        10'b1000010100: data <= 21'h000125; 
        10'b1000010101: data <= 21'h1ffcc3; 
        10'b1000010110: data <= 21'h00020c; 
        10'b1000010111: data <= 21'h1ff789; 
        10'b1000011000: data <= 21'h1ff21c; 
        10'b1000011001: data <= 21'h1fe9b8; 
        10'b1000011010: data <= 21'h1feeb1; 
        10'b1000011011: data <= 21'h000139; 
        10'b1000011100: data <= 21'h000f31; 
        10'b1000011101: data <= 21'h0017dc; 
        10'b1000011110: data <= 21'h001fc6; 
        10'b1000011111: data <= 21'h0032a4; 
        10'b1000100000: data <= 21'h0038fa; 
        10'b1000100001: data <= 21'h001d60; 
        10'b1000100010: data <= 21'h001a3e; 
        10'b1000100011: data <= 21'h001b6f; 
        10'b1000100100: data <= 21'h001387; 
        10'b1000100101: data <= 21'h00100d; 
        10'b1000100110: data <= 21'h00190b; 
        10'b1000100111: data <= 21'h00110f; 
        10'b1000101000: data <= 21'h000b0a; 
        10'b1000101001: data <= 21'h000260; 
        10'b1000101010: data <= 21'h1ffc02; 
        10'b1000101011: data <= 21'h1ffb11; 
        10'b1000101100: data <= 21'h1ffad6; 
        10'b1000101101: data <= 21'h1fff2b; 
        10'b1000101110: data <= 21'h1ffd86; 
        10'b1000101111: data <= 21'h0003a5; 
        10'b1000110000: data <= 21'h1ffdc2; 
        10'b1000110001: data <= 21'h1ffcbe; 
        10'b1000110010: data <= 21'h1ffedc; 
        10'b1000110011: data <= 21'h1ffc29; 
        10'b1000110100: data <= 21'h1fee3a; 
        10'b1000110101: data <= 21'h1feac0; 
        10'b1000110110: data <= 21'h1fed99; 
        10'b1000110111: data <= 21'h1ff87b; 
        10'b1000111000: data <= 21'h000507; 
        10'b1000111001: data <= 21'h000ff9; 
        10'b1000111010: data <= 21'h001a4e; 
        10'b1000111011: data <= 21'h001188; 
        10'b1000111100: data <= 21'h002285; 
        10'b1000111101: data <= 21'h002963; 
        10'b1000111110: data <= 21'h003120; 
        10'b1000111111: data <= 21'h0029d2; 
        10'b1001000000: data <= 21'h0016ac; 
        10'b1001000001: data <= 21'h000e80; 
        10'b1001000010: data <= 21'h001c28; 
        10'b1001000011: data <= 21'h0013da; 
        10'b1001000100: data <= 21'h000d77; 
        10'b1001000101: data <= 21'h1ffd3c; 
        10'b1001000110: data <= 21'h1ff591; 
        10'b1001000111: data <= 21'h0000ae; 
        10'b1001001000: data <= 21'h1ffd79; 
        10'b1001001001: data <= 21'h1ffebd; 
        10'b1001001010: data <= 21'h1ffcd7; 
        10'b1001001011: data <= 21'h0000ab; 
        10'b1001001100: data <= 21'h1fff98; 
        10'b1001001101: data <= 21'h00006a; 
        10'b1001001110: data <= 21'h000155; 
        10'b1001001111: data <= 21'h1ffea5; 
        10'b1001010000: data <= 21'h1ff944; 
        10'b1001010001: data <= 21'h1ff15e; 
        10'b1001010010: data <= 21'h1fe726; 
        10'b1001010011: data <= 21'h1ff4c0; 
        10'b1001010100: data <= 21'h1ff943; 
        10'b1001010101: data <= 21'h000c05; 
        10'b1001010110: data <= 21'h0015d4; 
        10'b1001010111: data <= 21'h001f0c; 
        10'b1001011000: data <= 21'h0027ef; 
        10'b1001011001: data <= 21'h00288e; 
        10'b1001011010: data <= 21'h00220b; 
        10'b1001011011: data <= 21'h001d59; 
        10'b1001011100: data <= 21'h001250; 
        10'b1001011101: data <= 21'h00190b; 
        10'b1001011110: data <= 21'h001759; 
        10'b1001011111: data <= 21'h000eec; 
        10'b1001100000: data <= 21'h0001fc; 
        10'b1001100001: data <= 21'h1ff818; 
        10'b1001100010: data <= 21'h1ff4ec; 
        10'b1001100011: data <= 21'h1ff98f; 
        10'b1001100100: data <= 21'h000060; 
        10'b1001100101: data <= 21'h1ffbd4; 
        10'b1001100110: data <= 21'h1fff19; 
        10'b1001100111: data <= 21'h1ffdaf; 
        10'b1001101000: data <= 21'h1ffdaa; 
        10'b1001101001: data <= 21'h1fff9a; 
        10'b1001101010: data <= 21'h0003fb; 
        10'b1001101011: data <= 21'h000114; 
        10'b1001101100: data <= 21'h1ffda6; 
        10'b1001101101: data <= 21'h1ff340; 
        10'b1001101110: data <= 21'h1ff0dc; 
        10'b1001101111: data <= 21'h1febb0; 
        10'b1001110000: data <= 21'h1ff274; 
        10'b1001110001: data <= 21'h1ff9da; 
        10'b1001110010: data <= 21'h1ffaf2; 
        10'b1001110011: data <= 21'h000274; 
        10'b1001110100: data <= 21'h000bad; 
        10'b1001110101: data <= 21'h00050e; 
        10'b1001110110: data <= 21'h000441; 
        10'b1001110111: data <= 21'h000c9a; 
        10'b1001111000: data <= 21'h000962; 
        10'b1001111001: data <= 21'h000015; 
        10'b1001111010: data <= 21'h1ffcdd; 
        10'b1001111011: data <= 21'h1ff1ea; 
        10'b1001111100: data <= 21'h1ff273; 
        10'b1001111101: data <= 21'h1ff4ba; 
        10'b1001111110: data <= 21'h1ff576; 
        10'b1001111111: data <= 21'h1ffefc; 
        10'b1010000000: data <= 21'h1ffe28; 
        10'b1010000001: data <= 21'h1ffc13; 
        10'b1010000010: data <= 21'h00044d; 
        10'b1010000011: data <= 21'h0001a8; 
        10'b1010000100: data <= 21'h000374; 
        10'b1010000101: data <= 21'h1ffea4; 
        10'b1010000110: data <= 21'h1ffe12; 
        10'b1010000111: data <= 21'h000066; 
        10'b1010001000: data <= 21'h000137; 
        10'b1010001001: data <= 21'h1ffabb; 
        10'b1010001010: data <= 21'h1ff7c3; 
        10'b1010001011: data <= 21'h1fedea; 
        10'b1010001100: data <= 21'h1fe922; 
        10'b1010001101: data <= 21'h1fdf1a; 
        10'b1010001110: data <= 21'h1fdf43; 
        10'b1010001111: data <= 21'h1fd9d9; 
        10'b1010010000: data <= 21'h1fe87d; 
        10'b1010010001: data <= 21'h1fed7a; 
        10'b1010010010: data <= 21'h1ff18f; 
        10'b1010010011: data <= 21'h1fea86; 
        10'b1010010100: data <= 21'h1fe3c7; 
        10'b1010010101: data <= 21'h1fdffe; 
        10'b1010010110: data <= 21'h1fe6c5; 
        10'b1010010111: data <= 21'h1ff47f; 
        10'b1010011000: data <= 21'h1ff44b; 
        10'b1010011001: data <= 21'h1ff5c0; 
        10'b1010011010: data <= 21'h1ffc58; 
        10'b1010011011: data <= 21'h000082; 
        10'b1010011100: data <= 21'h1ffbbb; 
        10'b1010011101: data <= 21'h1ffc7b; 
        10'b1010011110: data <= 21'h1ffe7f; 
        10'b1010011111: data <= 21'h1fff91; 
        10'b1010100000: data <= 21'h000279; 
        10'b1010100001: data <= 21'h0001fe; 
        10'b1010100010: data <= 21'h00015c; 
        10'b1010100011: data <= 21'h1ffbf1; 
        10'b1010100100: data <= 21'h1ffcc7; 
        10'b1010100101: data <= 21'h1ffe7c; 
        10'b1010100110: data <= 21'h1ffc1b; 
        10'b1010100111: data <= 21'h1ff9b2; 
        10'b1010101000: data <= 21'h1ffb03; 
        10'b1010101001: data <= 21'h1ff807; 
        10'b1010101010: data <= 21'h1ff40e; 
        10'b1010101011: data <= 21'h1ff0e2; 
        10'b1010101100: data <= 21'h1fee6c; 
        10'b1010101101: data <= 21'h1feecd; 
        10'b1010101110: data <= 21'h1febec; 
        10'b1010101111: data <= 21'h1febf1; 
        10'b1010110000: data <= 21'h1feb06; 
        10'b1010110001: data <= 21'h1feffe; 
        10'b1010110010: data <= 21'h1ffa72; 
        10'b1010110011: data <= 21'h1ffad5; 
        10'b1010110100: data <= 21'h1ffe32; 
        10'b1010110101: data <= 21'h1ffd25; 
        10'b1010110110: data <= 21'h00021f; 
        10'b1010110111: data <= 21'h1fff12; 
        10'b1010111000: data <= 21'h1ffbd0; 
        10'b1010111001: data <= 21'h1ffeae; 
        10'b1010111010: data <= 21'h1ffce2; 
        10'b1010111011: data <= 21'h1ffcf6; 
        10'b1010111100: data <= 21'h0003e9; 
        10'b1010111101: data <= 21'h1ffc5d; 
        10'b1010111110: data <= 21'h000112; 
        10'b1010111111: data <= 21'h1ffe24; 
        10'b1011000000: data <= 21'h1ffd26; 
        10'b1011000001: data <= 21'h1fff76; 
        10'b1011000010: data <= 21'h00029a; 
        10'b1011000011: data <= 21'h1fffcb; 
        10'b1011000100: data <= 21'h1ffb90; 
        10'b1011000101: data <= 21'h00019c; 
        10'b1011000110: data <= 21'h1ffbac; 
        10'b1011000111: data <= 21'h1fff55; 
        10'b1011001000: data <= 21'h000037; 
        10'b1011001001: data <= 21'h1ffb6b; 
        10'b1011001010: data <= 21'h1ffd7a; 
        10'b1011001011: data <= 21'h1ffe75; 
        10'b1011001100: data <= 21'h1fff96; 
        10'b1011001101: data <= 21'h1ffc02; 
        10'b1011001110: data <= 21'h1ffda9; 
        10'b1011001111: data <= 21'h1ffb97; 
        10'b1011010000: data <= 21'h1ffc86; 
        10'b1011010001: data <= 21'h00008d; 
        10'b1011010010: data <= 21'h1ffe55; 
        10'b1011010011: data <= 21'h00032d; 
        10'b1011010100: data <= 21'h00047e; 
        10'b1011010101: data <= 21'h0003f8; 
        10'b1011010110: data <= 21'h00002e; 
        10'b1011010111: data <= 21'h0002fa; 
        10'b1011011000: data <= 21'h000437; 
        10'b1011011001: data <= 21'h1fffce; 
        10'b1011011010: data <= 21'h0000c5; 
        10'b1011011011: data <= 21'h1fff32; 
        10'b1011011100: data <= 21'h1ffda0; 
        10'b1011011101: data <= 21'h00038e; 
        10'b1011011110: data <= 21'h0002ad; 
        10'b1011011111: data <= 21'h1ffdb2; 
        10'b1011100000: data <= 21'h1ffea0; 
        10'b1011100001: data <= 21'h000202; 
        10'b1011100010: data <= 21'h1ffe56; 
        10'b1011100011: data <= 21'h0000e2; 
        10'b1011100100: data <= 21'h1ffe3f; 
        10'b1011100101: data <= 21'h00029e; 
        10'b1011100110: data <= 21'h0002c1; 
        10'b1011100111: data <= 21'h1ffc70; 
        10'b1011101000: data <= 21'h1ffd4a; 
        10'b1011101001: data <= 21'h00039a; 
        10'b1011101010: data <= 21'h0002d4; 
        10'b1011101011: data <= 21'h1ffe9e; 
        10'b1011101100: data <= 21'h000289; 
        10'b1011101101: data <= 21'h1fff0a; 
        10'b1011101110: data <= 21'h1ffefe; 
        10'b1011101111: data <= 21'h000193; 
        10'b1011110000: data <= 21'h0001ce; 
        10'b1011110001: data <= 21'h1fff1e; 
        10'b1011110010: data <= 21'h1ffde2; 
        10'b1011110011: data <= 21'h1ffec9; 
        10'b1011110100: data <= 21'h000412; 
        10'b1011110101: data <= 21'h1fffcc; 
        10'b1011110110: data <= 21'h00024c; 
        10'b1011110111: data <= 21'h1ffdaa; 
        10'b1011111000: data <= 21'h00016c; 
        10'b1011111001: data <= 21'h1fffe3; 
        10'b1011111010: data <= 21'h0003d4; 
        10'b1011111011: data <= 21'h00008b; 
        10'b1011111100: data <= 21'h1fff7e; 
        10'b1011111101: data <= 21'h1ffb7f; 
        10'b1011111110: data <= 21'h1ffcf3; 
        10'b1011111111: data <= 21'h000163; 
        10'b1100000000: data <= 21'h1ffbee; 
        10'b1100000001: data <= 21'h1ffc99; 
        10'b1100000010: data <= 21'h1ffd6b; 
        10'b1100000011: data <= 21'h1ffbd8; 
        10'b1100000100: data <= 21'h1ffd2e; 
        10'b1100000101: data <= 21'h1ffe9c; 
        10'b1100000110: data <= 21'h1ffc46; 
        10'b1100000111: data <= 21'h1ffd30; 
        10'b1100001000: data <= 21'h1ffd91; 
        10'b1100001001: data <= 21'h1ffe04; 
        10'b1100001010: data <= 21'h0003c5; 
        10'b1100001011: data <= 21'h1ffc52; 
        10'b1100001100: data <= 21'h1ffd99; 
        10'b1100001101: data <= 21'h1ffc71; 
        10'b1100001110: data <= 21'h1ffd7f; 
        10'b1100001111: data <= 21'h0000b2; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 16) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 22'h3ffd28; 
        10'b0000000001: data <= 22'h0005cf; 
        10'b0000000010: data <= 22'h3ff970; 
        10'b0000000011: data <= 22'h3fff7f; 
        10'b0000000100: data <= 22'h3fffc8; 
        10'b0000000101: data <= 22'h3fff1c; 
        10'b0000000110: data <= 22'h00030d; 
        10'b0000000111: data <= 22'h000937; 
        10'b0000001000: data <= 22'h3ff9f3; 
        10'b0000001001: data <= 22'h3ffbfc; 
        10'b0000001010: data <= 22'h3ffc3d; 
        10'b0000001011: data <= 22'h3ffa38; 
        10'b0000001100: data <= 22'h0002fc; 
        10'b0000001101: data <= 22'h00086b; 
        10'b0000001110: data <= 22'h0004bb; 
        10'b0000001111: data <= 22'h3ff84d; 
        10'b0000010000: data <= 22'h3ffef1; 
        10'b0000010001: data <= 22'h000937; 
        10'b0000010010: data <= 22'h000190; 
        10'b0000010011: data <= 22'h3fff2f; 
        10'b0000010100: data <= 22'h3ff8e9; 
        10'b0000010101: data <= 22'h3ffb44; 
        10'b0000010110: data <= 22'h00022c; 
        10'b0000010111: data <= 22'h000814; 
        10'b0000011000: data <= 22'h00045b; 
        10'b0000011001: data <= 22'h000550; 
        10'b0000011010: data <= 22'h3ff8cc; 
        10'b0000011011: data <= 22'h3ff919; 
        10'b0000011100: data <= 22'h0005ee; 
        10'b0000011101: data <= 22'h0004b3; 
        10'b0000011110: data <= 22'h0005f9; 
        10'b0000011111: data <= 22'h3ffe7a; 
        10'b0000100000: data <= 22'h3ff7ec; 
        10'b0000100001: data <= 22'h3ffb2e; 
        10'b0000100010: data <= 22'h00041f; 
        10'b0000100011: data <= 22'h000d6a; 
        10'b0000100100: data <= 22'h000919; 
        10'b0000100101: data <= 22'h0002bb; 
        10'b0000100110: data <= 22'h000b01; 
        10'b0000100111: data <= 22'h000bc0; 
        10'b0000101000: data <= 22'h000c85; 
        10'b0000101001: data <= 22'h000bcb; 
        10'b0000101010: data <= 22'h00076d; 
        10'b0000101011: data <= 22'h0007f2; 
        10'b0000101100: data <= 22'h3ff784; 
        10'b0000101101: data <= 22'h000790; 
        10'b0000101110: data <= 22'h000a41; 
        10'b0000101111: data <= 22'h0005d7; 
        10'b0000110000: data <= 22'h3ffe5a; 
        10'b0000110001: data <= 22'h3ffaca; 
        10'b0000110010: data <= 22'h000ae3; 
        10'b0000110011: data <= 22'h000837; 
        10'b0000110100: data <= 22'h3ffc9f; 
        10'b0000110101: data <= 22'h00092c; 
        10'b0000110110: data <= 22'h3ffe6b; 
        10'b0000110111: data <= 22'h0006c9; 
        10'b0000111000: data <= 22'h3ffaa7; 
        10'b0000111001: data <= 22'h3ff990; 
        10'b0000111010: data <= 22'h3ff7e9; 
        10'b0000111011: data <= 22'h3fff35; 
        10'b0000111100: data <= 22'h00048f; 
        10'b0000111101: data <= 22'h0002d0; 
        10'b0000111110: data <= 22'h0004aa; 
        10'b0000111111: data <= 22'h000d1f; 
        10'b0001000000: data <= 22'h000955; 
        10'b0001000001: data <= 22'h0013e2; 
        10'b0001000010: data <= 22'h001904; 
        10'b0001000011: data <= 22'h001c45; 
        10'b0001000100: data <= 22'h001c55; 
        10'b0001000101: data <= 22'h001dc4; 
        10'b0001000110: data <= 22'h000f16; 
        10'b0001000111: data <= 22'h000ab2; 
        10'b0001001000: data <= 22'h0018d8; 
        10'b0001001001: data <= 22'h000af6; 
        10'b0001001010: data <= 22'h000aaa; 
        10'b0001001011: data <= 22'h000bad; 
        10'b0001001100: data <= 22'h000b6b; 
        10'b0001001101: data <= 22'h0005c8; 
        10'b0001001110: data <= 22'h00079c; 
        10'b0001001111: data <= 22'h00016c; 
        10'b0001010000: data <= 22'h000430; 
        10'b0001010001: data <= 22'h3ffd9d; 
        10'b0001010010: data <= 22'h3ff794; 
        10'b0001010011: data <= 22'h000294; 
        10'b0001010100: data <= 22'h3ff8da; 
        10'b0001010101: data <= 22'h0000d8; 
        10'b0001010110: data <= 22'h0006bd; 
        10'b0001010111: data <= 22'h0003e4; 
        10'b0001011000: data <= 22'h0008d7; 
        10'b0001011001: data <= 22'h3ff84f; 
        10'b0001011010: data <= 22'h000996; 
        10'b0001011011: data <= 22'h000a82; 
        10'b0001011100: data <= 22'h000c82; 
        10'b0001011101: data <= 22'h001959; 
        10'b0001011110: data <= 22'h001675; 
        10'b0001011111: data <= 22'h001c1f; 
        10'b0001100000: data <= 22'h001b71; 
        10'b0001100001: data <= 22'h001a6a; 
        10'b0001100010: data <= 22'h0026dc; 
        10'b0001100011: data <= 22'h0024a8; 
        10'b0001100100: data <= 22'h0016ca; 
        10'b0001100101: data <= 22'h001cc5; 
        10'b0001100110: data <= 22'h002e39; 
        10'b0001100111: data <= 22'h002e18; 
        10'b0001101000: data <= 22'h00312b; 
        10'b0001101001: data <= 22'h002b8d; 
        10'b0001101010: data <= 22'h002c19; 
        10'b0001101011: data <= 22'h00199d; 
        10'b0001101100: data <= 22'h0016bc; 
        10'b0001101101: data <= 22'h00058f; 
        10'b0001101110: data <= 22'h3ffc18; 
        10'b0001101111: data <= 22'h000507; 
        10'b0001110000: data <= 22'h000153; 
        10'b0001110001: data <= 22'h3ffe52; 
        10'b0001110010: data <= 22'h3fff68; 
        10'b0001110011: data <= 22'h0007d0; 
        10'b0001110100: data <= 22'h0006b9; 
        10'b0001110101: data <= 22'h000274; 
        10'b0001110110: data <= 22'h00027e; 
        10'b0001110111: data <= 22'h000fb4; 
        10'b0001111000: data <= 22'h3ffe3f; 
        10'b0001111001: data <= 22'h3ffcb8; 
        10'b0001111010: data <= 22'h000f31; 
        10'b0001111011: data <= 22'h0005b8; 
        10'b0001111100: data <= 22'h00070b; 
        10'b0001111101: data <= 22'h00028b; 
        10'b0001111110: data <= 22'h0005fb; 
        10'b0001111111: data <= 22'h0008fe; 
        10'b0010000000: data <= 22'h001ecf; 
        10'b0010000001: data <= 22'h001e82; 
        10'b0010000010: data <= 22'h002fc6; 
        10'b0010000011: data <= 22'h003092; 
        10'b0010000100: data <= 22'h003d4a; 
        10'b0010000101: data <= 22'h0043ff; 
        10'b0010000110: data <= 22'h003a7f; 
        10'b0010000111: data <= 22'h002748; 
        10'b0010001000: data <= 22'h000591; 
        10'b0010001001: data <= 22'h000a6d; 
        10'b0010001010: data <= 22'h000173; 
        10'b0010001011: data <= 22'h3ffffe; 
        10'b0010001100: data <= 22'h000193; 
        10'b0010001101: data <= 22'h0004c0; 
        10'b0010001110: data <= 22'h0002b5; 
        10'b0010001111: data <= 22'h3ffc63; 
        10'b0010010000: data <= 22'h3ff982; 
        10'b0010010001: data <= 22'h3fff49; 
        10'b0010010010: data <= 22'h3ffa90; 
        10'b0010010011: data <= 22'h3ff53c; 
        10'b0010010100: data <= 22'h000811; 
        10'b0010010101: data <= 22'h3ff59c; 
        10'b0010010110: data <= 22'h0003c0; 
        10'b0010010111: data <= 22'h3fdc52; 
        10'b0010011000: data <= 22'h3fed1c; 
        10'b0010011001: data <= 22'h3ff2f4; 
        10'b0010011010: data <= 22'h3ffb34; 
        10'b0010011011: data <= 22'h3fef26; 
        10'b0010011100: data <= 22'h3fef27; 
        10'b0010011101: data <= 22'h00033e; 
        10'b0010011110: data <= 22'h0016ec; 
        10'b0010011111: data <= 22'h002af7; 
        10'b0010100000: data <= 22'h002548; 
        10'b0010100001: data <= 22'h002153; 
        10'b0010100010: data <= 22'h001a4b; 
        10'b0010100011: data <= 22'h00120a; 
        10'b0010100100: data <= 22'h3ffde8; 
        10'b0010100101: data <= 22'h0000e8; 
        10'b0010100110: data <= 22'h3ff6f0; 
        10'b0010100111: data <= 22'h00088f; 
        10'b0010101000: data <= 22'h3ffed3; 
        10'b0010101001: data <= 22'h0007b5; 
        10'b0010101010: data <= 22'h000730; 
        10'b0010101011: data <= 22'h3ff6b9; 
        10'b0010101100: data <= 22'h000349; 
        10'b0010101101: data <= 22'h3ffe89; 
        10'b0010101110: data <= 22'h0002f9; 
        10'b0010101111: data <= 22'h000039; 
        10'b0010110000: data <= 22'h3ff2bf; 
        10'b0010110001: data <= 22'h3fefd9; 
        10'b0010110010: data <= 22'h3fd6e9; 
        10'b0010110011: data <= 22'h3fca48; 
        10'b0010110100: data <= 22'h3fe0c9; 
        10'b0010110101: data <= 22'h3fc2c1; 
        10'b0010110110: data <= 22'h3fe4fa; 
        10'b0010110111: data <= 22'h3fec29; 
        10'b0010111000: data <= 22'h3fe3bf; 
        10'b0010111001: data <= 22'h3fe708; 
        10'b0010111010: data <= 22'h3ff911; 
        10'b0010111011: data <= 22'h3fef40; 
        10'b0010111100: data <= 22'h3fe4da; 
        10'b0010111101: data <= 22'h3fe61f; 
        10'b0010111110: data <= 22'h3fd7c4; 
        10'b0010111111: data <= 22'h3fe5c2; 
        10'b0011000000: data <= 22'h3fea3a; 
        10'b0011000001: data <= 22'h3fe90c; 
        10'b0011000010: data <= 22'h3ffc93; 
        10'b0011000011: data <= 22'h00077a; 
        10'b0011000100: data <= 22'h0002f8; 
        10'b0011000101: data <= 22'h000472; 
        10'b0011000110: data <= 22'h000045; 
        10'b0011000111: data <= 22'h3ffe87; 
        10'b0011001000: data <= 22'h000080; 
        10'b0011001001: data <= 22'h3ff809; 
        10'b0011001010: data <= 22'h3fefdc; 
        10'b0011001011: data <= 22'h3ffd67; 
        10'b0011001100: data <= 22'h3fe919; 
        10'b0011001101: data <= 22'h3fe38d; 
        10'b0011001110: data <= 22'h3fd699; 
        10'b0011001111: data <= 22'h3fdf75; 
        10'b0011010000: data <= 22'h3fc585; 
        10'b0011010001: data <= 22'h3fbe77; 
        10'b0011010010: data <= 22'h3fdda3; 
        10'b0011010011: data <= 22'h3fdf66; 
        10'b0011010100: data <= 22'h3fcce9; 
        10'b0011010101: data <= 22'h3fcfa3; 
        10'b0011010110: data <= 22'h3fc407; 
        10'b0011010111: data <= 22'h3faea3; 
        10'b0011011000: data <= 22'h3facf7; 
        10'b0011011001: data <= 22'h3fba8d; 
        10'b0011011010: data <= 22'h3fb75b; 
        10'b0011011011: data <= 22'h3fc69f; 
        10'b0011011100: data <= 22'h3fea12; 
        10'b0011011101: data <= 22'h3fec29; 
        10'b0011011110: data <= 22'h3ff82c; 
        10'b0011011111: data <= 22'h3ffa06; 
        10'b0011100000: data <= 22'h3ffd1d; 
        10'b0011100001: data <= 22'h3ffd8d; 
        10'b0011100010: data <= 22'h0008c7; 
        10'b0011100011: data <= 22'h3ff4c7; 
        10'b0011100100: data <= 22'h3ff6ab; 
        10'b0011100101: data <= 22'h3ff393; 
        10'b0011100110: data <= 22'h3fe0d0; 
        10'b0011100111: data <= 22'h3ff928; 
        10'b0011101000: data <= 22'h3ff47d; 
        10'b0011101001: data <= 22'h3fdf63; 
        10'b0011101010: data <= 22'h3fd9e9; 
        10'b0011101011: data <= 22'h3fd457; 
        10'b0011101100: data <= 22'h3fcb72; 
        10'b0011101101: data <= 22'h3fc30d; 
        10'b0011101110: data <= 22'h3fc49d; 
        10'b0011101111: data <= 22'h3fc08f; 
        10'b0011110000: data <= 22'h3fb4c9; 
        10'b0011110001: data <= 22'h3fa95b; 
        10'b0011110010: data <= 22'h3f858f; 
        10'b0011110011: data <= 22'h3f8e07; 
        10'b0011110100: data <= 22'h3f9a18; 
        10'b0011110101: data <= 22'h3f9b16; 
        10'b0011110110: data <= 22'h3fb97a; 
        10'b0011110111: data <= 22'h3fc1e3; 
        10'b0011111000: data <= 22'h3fd93a; 
        10'b0011111001: data <= 22'h3fe793; 
        10'b0011111010: data <= 22'h3fee78; 
        10'b0011111011: data <= 22'h000299; 
        10'b0011111100: data <= 22'h3ffebc; 
        10'b0011111101: data <= 22'h3ff92d; 
        10'b0011111110: data <= 22'h3ffc16; 
        10'b0011111111: data <= 22'h3ff83b; 
        10'b0100000000: data <= 22'h00003b; 
        10'b0100000001: data <= 22'h3ff8d8; 
        10'b0100000010: data <= 22'h3ff51f; 
        10'b0100000011: data <= 22'h3ff9b3; 
        10'b0100000100: data <= 22'h000774; 
        10'b0100000101: data <= 22'h3fec51; 
        10'b0100000110: data <= 22'h3fdac5; 
        10'b0100000111: data <= 22'h3fe373; 
        10'b0100001000: data <= 22'h3fed9d; 
        10'b0100001001: data <= 22'h3fdd52; 
        10'b0100001010: data <= 22'h3fe03b; 
        10'b0100001011: data <= 22'h3fba80; 
        10'b0100001100: data <= 22'h3faf06; 
        10'b0100001101: data <= 22'h3f8ab2; 
        10'b0100001110: data <= 22'h3f82df; 
        10'b0100001111: data <= 22'h3f99d0; 
        10'b0100010000: data <= 22'h3fac2e; 
        10'b0100010001: data <= 22'h3fbd53; 
        10'b0100010010: data <= 22'h3fb2c7; 
        10'b0100010011: data <= 22'h3fce5d; 
        10'b0100010100: data <= 22'h3fda22; 
        10'b0100010101: data <= 22'h3fe3e6; 
        10'b0100010110: data <= 22'h3ff470; 
        10'b0100010111: data <= 22'h000613; 
        10'b0100011000: data <= 22'h3ffa1e; 
        10'b0100011001: data <= 22'h0007ad; 
        10'b0100011010: data <= 22'h000532; 
        10'b0100011011: data <= 22'h3ff6ff; 
        10'b0100011100: data <= 22'h3ff2e6; 
        10'b0100011101: data <= 22'h000353; 
        10'b0100011110: data <= 22'h000acd; 
        10'b0100011111: data <= 22'h000a61; 
        10'b0100100000: data <= 22'h002600; 
        10'b0100100001: data <= 22'h3fff36; 
        10'b0100100010: data <= 22'h00078e; 
        10'b0100100011: data <= 22'h000325; 
        10'b0100100100: data <= 22'h3fe904; 
        10'b0100100101: data <= 22'h3ff060; 
        10'b0100100110: data <= 22'h3fddb5; 
        10'b0100100111: data <= 22'h3fb810; 
        10'b0100101000: data <= 22'h3fb6da; 
        10'b0100101001: data <= 22'h3faa3b; 
        10'b0100101010: data <= 22'h3fa6b2; 
        10'b0100101011: data <= 22'h3fb8b1; 
        10'b0100101100: data <= 22'h3fcf96; 
        10'b0100101101: data <= 22'h3fdd54; 
        10'b0100101110: data <= 22'h3fd261; 
        10'b0100101111: data <= 22'h3ffb39; 
        10'b0100110000: data <= 22'h3fe253; 
        10'b0100110001: data <= 22'h3feb60; 
        10'b0100110010: data <= 22'h3ff9df; 
        10'b0100110011: data <= 22'h3ffd09; 
        10'b0100110100: data <= 22'h3ffb3a; 
        10'b0100110101: data <= 22'h00031d; 
        10'b0100110110: data <= 22'h3ffac4; 
        10'b0100110111: data <= 22'h3fff40; 
        10'b0100111000: data <= 22'h3fface; 
        10'b0100111001: data <= 22'h00015a; 
        10'b0100111010: data <= 22'h3ffd2f; 
        10'b0100111011: data <= 22'h001fca; 
        10'b0100111100: data <= 22'h0016bf; 
        10'b0100111101: data <= 22'h000af1; 
        10'b0100111110: data <= 22'h000dc1; 
        10'b0100111111: data <= 22'h0009bb; 
        10'b0101000000: data <= 22'h0009c0; 
        10'b0101000001: data <= 22'h000190; 
        10'b0101000010: data <= 22'h3fef6f; 
        10'b0101000011: data <= 22'h3fc6f3; 
        10'b0101000100: data <= 22'h3fca7e; 
        10'b0101000101: data <= 22'h3fd276; 
        10'b0101000110: data <= 22'h3fd244; 
        10'b0101000111: data <= 22'h3fdc66; 
        10'b0101001000: data <= 22'h3fef5f; 
        10'b0101001001: data <= 22'h000668; 
        10'b0101001010: data <= 22'h0015d3; 
        10'b0101001011: data <= 22'h0021f3; 
        10'b0101001100: data <= 22'h3fffeb; 
        10'b0101001101: data <= 22'h3fedf1; 
        10'b0101001110: data <= 22'h3ff876; 
        10'b0101001111: data <= 22'h3ffd3e; 
        10'b0101010000: data <= 22'h3ffb35; 
        10'b0101010001: data <= 22'h3ffd6f; 
        10'b0101010010: data <= 22'h3ff836; 
        10'b0101010011: data <= 22'h3ffc47; 
        10'b0101010100: data <= 22'h000489; 
        10'b0101010101: data <= 22'h000ee2; 
        10'b0101010110: data <= 22'h0016bb; 
        10'b0101010111: data <= 22'h001dd0; 
        10'b0101011000: data <= 22'h000dd3; 
        10'b0101011001: data <= 22'h00135d; 
        10'b0101011010: data <= 22'h000dab; 
        10'b0101011011: data <= 22'h0023ed; 
        10'b0101011100: data <= 22'h002292; 
        10'b0101011101: data <= 22'h0018bd; 
        10'b0101011110: data <= 22'h3feacd; 
        10'b0101011111: data <= 22'h3fd9b8; 
        10'b0101100000: data <= 22'h3ffe65; 
        10'b0101100001: data <= 22'h3ffc77; 
        10'b0101100010: data <= 22'h3fda87; 
        10'b0101100011: data <= 22'h3fdc17; 
        10'b0101100100: data <= 22'h3ffb8b; 
        10'b0101100101: data <= 22'h001448; 
        10'b0101100110: data <= 22'h003100; 
        10'b0101100111: data <= 22'h0056f0; 
        10'b0101101000: data <= 22'h002ec3; 
        10'b0101101001: data <= 22'h3ff2a9; 
        10'b0101101010: data <= 22'h3ff0af; 
        10'b0101101011: data <= 22'h3ffb60; 
        10'b0101101100: data <= 22'h3ffb72; 
        10'b0101101101: data <= 22'h000814; 
        10'b0101101110: data <= 22'h00062c; 
        10'b0101101111: data <= 22'h3ff737; 
        10'b0101110000: data <= 22'h3ff3fe; 
        10'b0101110001: data <= 22'h0004d7; 
        10'b0101110010: data <= 22'h0025bb; 
        10'b0101110011: data <= 22'h00144d; 
        10'b0101110100: data <= 22'h001173; 
        10'b0101110101: data <= 22'h0008a0; 
        10'b0101110110: data <= 22'h00249f; 
        10'b0101110111: data <= 22'h001e90; 
        10'b0101111000: data <= 22'h001c0a; 
        10'b0101111001: data <= 22'h0004f3; 
        10'b0101111010: data <= 22'h3ffad1; 
        10'b0101111011: data <= 22'h3fff1b; 
        10'b0101111100: data <= 22'h0002d7; 
        10'b0101111101: data <= 22'h3ff7c2; 
        10'b0101111110: data <= 22'h3fdf62; 
        10'b0101111111: data <= 22'h3ffbb6; 
        10'b0110000000: data <= 22'h3ff04f; 
        10'b0110000001: data <= 22'h001a14; 
        10'b0110000010: data <= 22'h0043d8; 
        10'b0110000011: data <= 22'h006b7c; 
        10'b0110000100: data <= 22'h003a11; 
        10'b0110000101: data <= 22'h3ffb5d; 
        10'b0110000110: data <= 22'h00002d; 
        10'b0110000111: data <= 22'h000545; 
        10'b0110001000: data <= 22'h3ffc24; 
        10'b0110001001: data <= 22'h0000d9; 
        10'b0110001010: data <= 22'h000618; 
        10'b0110001011: data <= 22'h000052; 
        10'b0110001100: data <= 22'h3ff34d; 
        10'b0110001101: data <= 22'h000d85; 
        10'b0110001110: data <= 22'h00229a; 
        10'b0110001111: data <= 22'h001dd2; 
        10'b0110010000: data <= 22'h00290c; 
        10'b0110010001: data <= 22'h002672; 
        10'b0110010010: data <= 22'h00299c; 
        10'b0110010011: data <= 22'h002d0c; 
        10'b0110010100: data <= 22'h000f2b; 
        10'b0110010101: data <= 22'h3fea06; 
        10'b0110010110: data <= 22'h000176; 
        10'b0110010111: data <= 22'h00125b; 
        10'b0110011000: data <= 22'h0008b1; 
        10'b0110011001: data <= 22'h3ff1b6; 
        10'b0110011010: data <= 22'h3ff21e; 
        10'b0110011011: data <= 22'h3ffe01; 
        10'b0110011100: data <= 22'h001d70; 
        10'b0110011101: data <= 22'h001d1b; 
        10'b0110011110: data <= 22'h004cd1; 
        10'b0110011111: data <= 22'h005964; 
        10'b0110100000: data <= 22'h003a9b; 
        10'b0110100001: data <= 22'h3fff2f; 
        10'b0110100010: data <= 22'h3fef39; 
        10'b0110100011: data <= 22'h3ff7be; 
        10'b0110100100: data <= 22'h000646; 
        10'b0110100101: data <= 22'h3ffcd1; 
        10'b0110100110: data <= 22'h00013a; 
        10'b0110100111: data <= 22'h3ff913; 
        10'b0110101000: data <= 22'h3fe7c0; 
        10'b0110101001: data <= 22'h3ffcf1; 
        10'b0110101010: data <= 22'h002413; 
        10'b0110101011: data <= 22'h002ff4; 
        10'b0110101100: data <= 22'h001ee0; 
        10'b0110101101: data <= 22'h003077; 
        10'b0110101110: data <= 22'h003d15; 
        10'b0110101111: data <= 22'h004a88; 
        10'b0110110000: data <= 22'h001379; 
        10'b0110110001: data <= 22'h3ffa99; 
        10'b0110110010: data <= 22'h001cc2; 
        10'b0110110011: data <= 22'h001a73; 
        10'b0110110100: data <= 22'h000418; 
        10'b0110110101: data <= 22'h3ff273; 
        10'b0110110110: data <= 22'h0002bb; 
        10'b0110110111: data <= 22'h000ed7; 
        10'b0110111000: data <= 22'h002270; 
        10'b0110111001: data <= 22'h002f45; 
        10'b0110111010: data <= 22'h002b6f; 
        10'b0110111011: data <= 22'h0035d2; 
        10'b0110111100: data <= 22'h001cb8; 
        10'b0110111101: data <= 22'h3ff146; 
        10'b0110111110: data <= 22'h3ff6d7; 
        10'b0110111111: data <= 22'h3ff6a0; 
        10'b0111000000: data <= 22'h0001ab; 
        10'b0111000001: data <= 22'h3ff927; 
        10'b0111000010: data <= 22'h3ff8e6; 
        10'b0111000011: data <= 22'h3ff825; 
        10'b0111000100: data <= 22'h3fdff2; 
        10'b0111000101: data <= 22'h3fee9c; 
        10'b0111000110: data <= 22'h003571; 
        10'b0111000111: data <= 22'h00369b; 
        10'b0111001000: data <= 22'h002421; 
        10'b0111001001: data <= 22'h0037be; 
        10'b0111001010: data <= 22'h005e8b; 
        10'b0111001011: data <= 22'h005dc6; 
        10'b0111001100: data <= 22'h001c9a; 
        10'b0111001101: data <= 22'h001101; 
        10'b0111001110: data <= 22'h0028c1; 
        10'b0111001111: data <= 22'h001581; 
        10'b0111010000: data <= 22'h3ff4c1; 
        10'b0111010001: data <= 22'h3fe9b5; 
        10'b0111010010: data <= 22'h0007b5; 
        10'b0111010011: data <= 22'h0017d1; 
        10'b0111010100: data <= 22'h000b15; 
        10'b0111010101: data <= 22'h000053; 
        10'b0111010110: data <= 22'h001640; 
        10'b0111010111: data <= 22'h000d54; 
        10'b0111011000: data <= 22'h3ff987; 
        10'b0111011001: data <= 22'h3feeac; 
        10'b0111011010: data <= 22'h3ff55f; 
        10'b0111011011: data <= 22'h3ffe8c; 
        10'b0111011100: data <= 22'h000193; 
        10'b0111011101: data <= 22'h000544; 
        10'b0111011110: data <= 22'h000743; 
        10'b0111011111: data <= 22'h3ffeba; 
        10'b0111100000: data <= 22'h3fd248; 
        10'b0111100001: data <= 22'h3fe816; 
        10'b0111100010: data <= 22'h001659; 
        10'b0111100011: data <= 22'h002a77; 
        10'b0111100100: data <= 22'h003052; 
        10'b0111100101: data <= 22'h003cf1; 
        10'b0111100110: data <= 22'h00692e; 
        10'b0111100111: data <= 22'h006ae3; 
        10'b0111101000: data <= 22'h00373a; 
        10'b0111101001: data <= 22'h001f1a; 
        10'b0111101010: data <= 22'h001f7b; 
        10'b0111101011: data <= 22'h0013df; 
        10'b0111101100: data <= 22'h3ffffd; 
        10'b0111101101: data <= 22'h0005be; 
        10'b0111101110: data <= 22'h002bcd; 
        10'b0111101111: data <= 22'h000f1f; 
        10'b0111110000: data <= 22'h000645; 
        10'b0111110001: data <= 22'h3ff4d4; 
        10'b0111110010: data <= 22'h000a05; 
        10'b0111110011: data <= 22'h3ffddd; 
        10'b0111110100: data <= 22'h3ff38e; 
        10'b0111110101: data <= 22'h3fe7c2; 
        10'b0111110110: data <= 22'h3ffc86; 
        10'b0111110111: data <= 22'h0003f4; 
        10'b0111111000: data <= 22'h3ffc6d; 
        10'b0111111001: data <= 22'h3ffb0f; 
        10'b0111111010: data <= 22'h3fffdd; 
        10'b0111111011: data <= 22'h3ff2a9; 
        10'b0111111100: data <= 22'h3fd51c; 
        10'b0111111101: data <= 22'h3fd621; 
        10'b0111111110: data <= 22'h3febb9; 
        10'b0111111111: data <= 22'h001d35; 
        10'b1000000000: data <= 22'h002ecc; 
        10'b1000000001: data <= 22'h002a89; 
        10'b1000000010: data <= 22'h0049a8; 
        10'b1000000011: data <= 22'h005ad9; 
        10'b1000000100: data <= 22'h006b0d; 
        10'b1000000101: data <= 22'h0031b9; 
        10'b1000000110: data <= 22'h000d73; 
        10'b1000000111: data <= 22'h001bac; 
        10'b1000001000: data <= 22'h002fc3; 
        10'b1000001001: data <= 22'h001efc; 
        10'b1000001010: data <= 22'h002697; 
        10'b1000001011: data <= 22'h00144f; 
        10'b1000001100: data <= 22'h00029e; 
        10'b1000001101: data <= 22'h0006c6; 
        10'b1000001110: data <= 22'h00077e; 
        10'b1000001111: data <= 22'h3ffbc2; 
        10'b1000010000: data <= 22'h3ff0ba; 
        10'b1000010001: data <= 22'h3ff4ba; 
        10'b1000010010: data <= 22'h3ff746; 
        10'b1000010011: data <= 22'h3ff6b7; 
        10'b1000010100: data <= 22'h00024b; 
        10'b1000010101: data <= 22'h3ff985; 
        10'b1000010110: data <= 22'h000418; 
        10'b1000010111: data <= 22'h3fef12; 
        10'b1000011000: data <= 22'h3fe439; 
        10'b1000011001: data <= 22'h3fd370; 
        10'b1000011010: data <= 22'h3fdd62; 
        10'b1000011011: data <= 22'h000273; 
        10'b1000011100: data <= 22'h001e61; 
        10'b1000011101: data <= 22'h002fb8; 
        10'b1000011110: data <= 22'h003f8c; 
        10'b1000011111: data <= 22'h006547; 
        10'b1000100000: data <= 22'h0071f4; 
        10'b1000100001: data <= 22'h003abf; 
        10'b1000100010: data <= 22'h00347b; 
        10'b1000100011: data <= 22'h0036dd; 
        10'b1000100100: data <= 22'h00270f; 
        10'b1000100101: data <= 22'h00201b; 
        10'b1000100110: data <= 22'h003216; 
        10'b1000100111: data <= 22'h00221e; 
        10'b1000101000: data <= 22'h001615; 
        10'b1000101001: data <= 22'h0004bf; 
        10'b1000101010: data <= 22'h3ff804; 
        10'b1000101011: data <= 22'h3ff623; 
        10'b1000101100: data <= 22'h3ff5ab; 
        10'b1000101101: data <= 22'h3ffe57; 
        10'b1000101110: data <= 22'h3ffb0c; 
        10'b1000101111: data <= 22'h00074b; 
        10'b1000110000: data <= 22'h3ffb85; 
        10'b1000110001: data <= 22'h3ff97c; 
        10'b1000110010: data <= 22'h3ffdb8; 
        10'b1000110011: data <= 22'h3ff853; 
        10'b1000110100: data <= 22'h3fdc75; 
        10'b1000110101: data <= 22'h3fd580; 
        10'b1000110110: data <= 22'h3fdb32; 
        10'b1000110111: data <= 22'h3ff0f6; 
        10'b1000111000: data <= 22'h000a0d; 
        10'b1000111001: data <= 22'h001ff1; 
        10'b1000111010: data <= 22'h00349b; 
        10'b1000111011: data <= 22'h002310; 
        10'b1000111100: data <= 22'h00450a; 
        10'b1000111101: data <= 22'h0052c5; 
        10'b1000111110: data <= 22'h00623f; 
        10'b1000111111: data <= 22'h0053a5; 
        10'b1001000000: data <= 22'h002d57; 
        10'b1001000001: data <= 22'h001d01; 
        10'b1001000010: data <= 22'h00384f; 
        10'b1001000011: data <= 22'h0027b5; 
        10'b1001000100: data <= 22'h001aef; 
        10'b1001000101: data <= 22'h3ffa78; 
        10'b1001000110: data <= 22'h3feb21; 
        10'b1001000111: data <= 22'h00015c; 
        10'b1001001000: data <= 22'h3ffaf3; 
        10'b1001001001: data <= 22'h3ffd7a; 
        10'b1001001010: data <= 22'h3ff9ae; 
        10'b1001001011: data <= 22'h000156; 
        10'b1001001100: data <= 22'h3fff2f; 
        10'b1001001101: data <= 22'h0000d4; 
        10'b1001001110: data <= 22'h0002aa; 
        10'b1001001111: data <= 22'h3ffd49; 
        10'b1001010000: data <= 22'h3ff288; 
        10'b1001010001: data <= 22'h3fe2bc; 
        10'b1001010010: data <= 22'h3fce4d; 
        10'b1001010011: data <= 22'h3fe980; 
        10'b1001010100: data <= 22'h3ff286; 
        10'b1001010101: data <= 22'h00180b; 
        10'b1001010110: data <= 22'h002ba8; 
        10'b1001010111: data <= 22'h003e19; 
        10'b1001011000: data <= 22'h004fde; 
        10'b1001011001: data <= 22'h00511c; 
        10'b1001011010: data <= 22'h004416; 
        10'b1001011011: data <= 22'h003ab1; 
        10'b1001011100: data <= 22'h0024a0; 
        10'b1001011101: data <= 22'h003216; 
        10'b1001011110: data <= 22'h002eb1; 
        10'b1001011111: data <= 22'h001dd9; 
        10'b1001100000: data <= 22'h0003f8; 
        10'b1001100001: data <= 22'h3ff02f; 
        10'b1001100010: data <= 22'h3fe9d8; 
        10'b1001100011: data <= 22'h3ff31e; 
        10'b1001100100: data <= 22'h0000c0; 
        10'b1001100101: data <= 22'h3ff7a9; 
        10'b1001100110: data <= 22'h3ffe33; 
        10'b1001100111: data <= 22'h3ffb5e; 
        10'b1001101000: data <= 22'h3ffb55; 
        10'b1001101001: data <= 22'h3fff33; 
        10'b1001101010: data <= 22'h0007f6; 
        10'b1001101011: data <= 22'h000228; 
        10'b1001101100: data <= 22'h3ffb4c; 
        10'b1001101101: data <= 22'h3fe680; 
        10'b1001101110: data <= 22'h3fe1b9; 
        10'b1001101111: data <= 22'h3fd760; 
        10'b1001110000: data <= 22'h3fe4e9; 
        10'b1001110001: data <= 22'h3ff3b3; 
        10'b1001110010: data <= 22'h3ff5e5; 
        10'b1001110011: data <= 22'h0004e7; 
        10'b1001110100: data <= 22'h00175a; 
        10'b1001110101: data <= 22'h000a1c; 
        10'b1001110110: data <= 22'h000883; 
        10'b1001110111: data <= 22'h001935; 
        10'b1001111000: data <= 22'h0012c3; 
        10'b1001111001: data <= 22'h000029; 
        10'b1001111010: data <= 22'h3ff9ba; 
        10'b1001111011: data <= 22'h3fe3d4; 
        10'b1001111100: data <= 22'h3fe4e6; 
        10'b1001111101: data <= 22'h3fe973; 
        10'b1001111110: data <= 22'h3feaed; 
        10'b1001111111: data <= 22'h3ffdf7; 
        10'b1010000000: data <= 22'h3ffc4f; 
        10'b1010000001: data <= 22'h3ff825; 
        10'b1010000010: data <= 22'h000899; 
        10'b1010000011: data <= 22'h000350; 
        10'b1010000100: data <= 22'h0006e7; 
        10'b1010000101: data <= 22'h3ffd47; 
        10'b1010000110: data <= 22'h3ffc25; 
        10'b1010000111: data <= 22'h0000cb; 
        10'b1010001000: data <= 22'h00026d; 
        10'b1010001001: data <= 22'h3ff576; 
        10'b1010001010: data <= 22'h3fef85; 
        10'b1010001011: data <= 22'h3fdbd4; 
        10'b1010001100: data <= 22'h3fd244; 
        10'b1010001101: data <= 22'h3fbe34; 
        10'b1010001110: data <= 22'h3fbe87; 
        10'b1010001111: data <= 22'h3fb3b2; 
        10'b1010010000: data <= 22'h3fd0fa; 
        10'b1010010001: data <= 22'h3fdaf3; 
        10'b1010010010: data <= 22'h3fe31e; 
        10'b1010010011: data <= 22'h3fd50d; 
        10'b1010010100: data <= 22'h3fc78e; 
        10'b1010010101: data <= 22'h3fbffd; 
        10'b1010010110: data <= 22'h3fcd8a; 
        10'b1010010111: data <= 22'h3fe8fe; 
        10'b1010011000: data <= 22'h3fe896; 
        10'b1010011001: data <= 22'h3feb80; 
        10'b1010011010: data <= 22'h3ff8b1; 
        10'b1010011011: data <= 22'h000104; 
        10'b1010011100: data <= 22'h3ff777; 
        10'b1010011101: data <= 22'h3ff8f5; 
        10'b1010011110: data <= 22'h3ffcfe; 
        10'b1010011111: data <= 22'h3fff21; 
        10'b1010100000: data <= 22'h0004f2; 
        10'b1010100001: data <= 22'h0003fc; 
        10'b1010100010: data <= 22'h0002b8; 
        10'b1010100011: data <= 22'h3ff7e2; 
        10'b1010100100: data <= 22'h3ff98e; 
        10'b1010100101: data <= 22'h3ffcf8; 
        10'b1010100110: data <= 22'h3ff836; 
        10'b1010100111: data <= 22'h3ff363; 
        10'b1010101000: data <= 22'h3ff607; 
        10'b1010101001: data <= 22'h3ff00e; 
        10'b1010101010: data <= 22'h3fe81c; 
        10'b1010101011: data <= 22'h3fe1c4; 
        10'b1010101100: data <= 22'h3fdcd8; 
        10'b1010101101: data <= 22'h3fdd99; 
        10'b1010101110: data <= 22'h3fd7d8; 
        10'b1010101111: data <= 22'h3fd7e2; 
        10'b1010110000: data <= 22'h3fd60d; 
        10'b1010110001: data <= 22'h3fdffc; 
        10'b1010110010: data <= 22'h3ff4e3; 
        10'b1010110011: data <= 22'h3ff5aa; 
        10'b1010110100: data <= 22'h3ffc64; 
        10'b1010110101: data <= 22'h3ffa4a; 
        10'b1010110110: data <= 22'h00043e; 
        10'b1010110111: data <= 22'h3ffe24; 
        10'b1010111000: data <= 22'h3ff7a0; 
        10'b1010111001: data <= 22'h3ffd5c; 
        10'b1010111010: data <= 22'h3ff9c3; 
        10'b1010111011: data <= 22'h3ff9ec; 
        10'b1010111100: data <= 22'h0007d2; 
        10'b1010111101: data <= 22'h3ff8b9; 
        10'b1010111110: data <= 22'h000224; 
        10'b1010111111: data <= 22'h3ffc49; 
        10'b1011000000: data <= 22'h3ffa4c; 
        10'b1011000001: data <= 22'h3ffeed; 
        10'b1011000010: data <= 22'h000534; 
        10'b1011000011: data <= 22'h3fff96; 
        10'b1011000100: data <= 22'h3ff720; 
        10'b1011000101: data <= 22'h000337; 
        10'b1011000110: data <= 22'h3ff758; 
        10'b1011000111: data <= 22'h3ffeaa; 
        10'b1011001000: data <= 22'h00006f; 
        10'b1011001001: data <= 22'h3ff6d6; 
        10'b1011001010: data <= 22'h3ffaf3; 
        10'b1011001011: data <= 22'h3ffcea; 
        10'b1011001100: data <= 22'h3fff2b; 
        10'b1011001101: data <= 22'h3ff803; 
        10'b1011001110: data <= 22'h3ffb52; 
        10'b1011001111: data <= 22'h3ff72e; 
        10'b1011010000: data <= 22'h3ff90d; 
        10'b1011010001: data <= 22'h00011a; 
        10'b1011010010: data <= 22'h3ffcaa; 
        10'b1011010011: data <= 22'h00065a; 
        10'b1011010100: data <= 22'h0008fc; 
        10'b1011010101: data <= 22'h0007ef; 
        10'b1011010110: data <= 22'h00005d; 
        10'b1011010111: data <= 22'h0005f5; 
        10'b1011011000: data <= 22'h00086e; 
        10'b1011011001: data <= 22'h3fff9b; 
        10'b1011011010: data <= 22'h00018a; 
        10'b1011011011: data <= 22'h3ffe64; 
        10'b1011011100: data <= 22'h3ffb41; 
        10'b1011011101: data <= 22'h00071b; 
        10'b1011011110: data <= 22'h000559; 
        10'b1011011111: data <= 22'h3ffb63; 
        10'b1011100000: data <= 22'h3ffd3f; 
        10'b1011100001: data <= 22'h000404; 
        10'b1011100010: data <= 22'h3ffcab; 
        10'b1011100011: data <= 22'h0001c4; 
        10'b1011100100: data <= 22'h3ffc7e; 
        10'b1011100101: data <= 22'h00053b; 
        10'b1011100110: data <= 22'h000581; 
        10'b1011100111: data <= 22'h3ff8e0; 
        10'b1011101000: data <= 22'h3ffa93; 
        10'b1011101001: data <= 22'h000733; 
        10'b1011101010: data <= 22'h0005a8; 
        10'b1011101011: data <= 22'h3ffd3b; 
        10'b1011101100: data <= 22'h000512; 
        10'b1011101101: data <= 22'h3ffe15; 
        10'b1011101110: data <= 22'h3ffdfc; 
        10'b1011101111: data <= 22'h000326; 
        10'b1011110000: data <= 22'h00039b; 
        10'b1011110001: data <= 22'h3ffe3d; 
        10'b1011110010: data <= 22'h3ffbc4; 
        10'b1011110011: data <= 22'h3ffd92; 
        10'b1011110100: data <= 22'h000825; 
        10'b1011110101: data <= 22'h3fff98; 
        10'b1011110110: data <= 22'h000499; 
        10'b1011110111: data <= 22'h3ffb55; 
        10'b1011111000: data <= 22'h0002d9; 
        10'b1011111001: data <= 22'h3fffc5; 
        10'b1011111010: data <= 22'h0007a7; 
        10'b1011111011: data <= 22'h000117; 
        10'b1011111100: data <= 22'h3ffefc; 
        10'b1011111101: data <= 22'h3ff6fd; 
        10'b1011111110: data <= 22'h3ff9e6; 
        10'b1011111111: data <= 22'h0002c6; 
        10'b1100000000: data <= 22'h3ff7db; 
        10'b1100000001: data <= 22'h3ff931; 
        10'b1100000010: data <= 22'h3ffad7; 
        10'b1100000011: data <= 22'h3ff7b1; 
        10'b1100000100: data <= 22'h3ffa5d; 
        10'b1100000101: data <= 22'h3ffd37; 
        10'b1100000110: data <= 22'h3ff88c; 
        10'b1100000111: data <= 22'h3ffa60; 
        10'b1100001000: data <= 22'h3ffb23; 
        10'b1100001001: data <= 22'h3ffc08; 
        10'b1100001010: data <= 22'h00078a; 
        10'b1100001011: data <= 22'h3ff8a4; 
        10'b1100001100: data <= 22'h3ffb32; 
        10'b1100001101: data <= 22'h3ff8e2; 
        10'b1100001110: data <= 22'h3ffaff; 
        10'b1100001111: data <= 22'h000163; 
      endcase 
    end 
  end 
endgenerate 
assign dout = data; 
endmodule
