`timescale 1ns / 1ps 
 
////////////////////////////////////////////////////////////////////////////////// 
// WEIGHT MEMORY (ROM) 
////////////////////////////////////////////////////////////////////////////////// 
module ROM_weights_4 #( 
    parameter int WGHT_INT = 6, // integer part 
    parameter int WGHT_FRC = 16 // fractional part 
)( 
    input logic clk, // clock 
    input logic [9:0] address,
    output [WGHT_INT + WGHT_FRC-1:0] dout 
); 

(* rom_style = "block" *) reg [WGHT_INT + WGHT_FRC-1:0] data;
generate 
  if (WGHT_FRC == 1) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 7'h00; 
        10'b0000000001: data <= 7'h00; 
        10'b0000000010: data <= 7'h00; 
        10'b0000000011: data <= 7'h00; 
        10'b0000000100: data <= 7'h00; 
        10'b0000000101: data <= 7'h00; 
        10'b0000000110: data <= 7'h00; 
        10'b0000000111: data <= 7'h00; 
        10'b0000001000: data <= 7'h00; 
        10'b0000001001: data <= 7'h00; 
        10'b0000001010: data <= 7'h00; 
        10'b0000001011: data <= 7'h00; 
        10'b0000001100: data <= 7'h00; 
        10'b0000001101: data <= 7'h00; 
        10'b0000001110: data <= 7'h00; 
        10'b0000001111: data <= 7'h00; 
        10'b0000010000: data <= 7'h00; 
        10'b0000010001: data <= 7'h00; 
        10'b0000010010: data <= 7'h00; 
        10'b0000010011: data <= 7'h00; 
        10'b0000010100: data <= 7'h00; 
        10'b0000010101: data <= 7'h00; 
        10'b0000010110: data <= 7'h00; 
        10'b0000010111: data <= 7'h00; 
        10'b0000011000: data <= 7'h00; 
        10'b0000011001: data <= 7'h00; 
        10'b0000011010: data <= 7'h00; 
        10'b0000011011: data <= 7'h00; 
        10'b0000011100: data <= 7'h00; 
        10'b0000011101: data <= 7'h00; 
        10'b0000011110: data <= 7'h00; 
        10'b0000011111: data <= 7'h00; 
        10'b0000100000: data <= 7'h00; 
        10'b0000100001: data <= 7'h00; 
        10'b0000100010: data <= 7'h00; 
        10'b0000100011: data <= 7'h00; 
        10'b0000100100: data <= 7'h00; 
        10'b0000100101: data <= 7'h00; 
        10'b0000100110: data <= 7'h00; 
        10'b0000100111: data <= 7'h00; 
        10'b0000101000: data <= 7'h00; 
        10'b0000101001: data <= 7'h00; 
        10'b0000101010: data <= 7'h00; 
        10'b0000101011: data <= 7'h00; 
        10'b0000101100: data <= 7'h00; 
        10'b0000101101: data <= 7'h00; 
        10'b0000101110: data <= 7'h00; 
        10'b0000101111: data <= 7'h00; 
        10'b0000110000: data <= 7'h00; 
        10'b0000110001: data <= 7'h00; 
        10'b0000110010: data <= 7'h00; 
        10'b0000110011: data <= 7'h00; 
        10'b0000110100: data <= 7'h00; 
        10'b0000110101: data <= 7'h00; 
        10'b0000110110: data <= 7'h00; 
        10'b0000110111: data <= 7'h00; 
        10'b0000111000: data <= 7'h00; 
        10'b0000111001: data <= 7'h00; 
        10'b0000111010: data <= 7'h00; 
        10'b0000111011: data <= 7'h00; 
        10'b0000111100: data <= 7'h00; 
        10'b0000111101: data <= 7'h00; 
        10'b0000111110: data <= 7'h00; 
        10'b0000111111: data <= 7'h00; 
        10'b0001000000: data <= 7'h00; 
        10'b0001000001: data <= 7'h00; 
        10'b0001000010: data <= 7'h00; 
        10'b0001000011: data <= 7'h00; 
        10'b0001000100: data <= 7'h00; 
        10'b0001000101: data <= 7'h00; 
        10'b0001000110: data <= 7'h00; 
        10'b0001000111: data <= 7'h00; 
        10'b0001001000: data <= 7'h00; 
        10'b0001001001: data <= 7'h00; 
        10'b0001001010: data <= 7'h00; 
        10'b0001001011: data <= 7'h00; 
        10'b0001001100: data <= 7'h00; 
        10'b0001001101: data <= 7'h00; 
        10'b0001001110: data <= 7'h00; 
        10'b0001001111: data <= 7'h00; 
        10'b0001010000: data <= 7'h00; 
        10'b0001010001: data <= 7'h00; 
        10'b0001010010: data <= 7'h00; 
        10'b0001010011: data <= 7'h00; 
        10'b0001010100: data <= 7'h00; 
        10'b0001010101: data <= 7'h00; 
        10'b0001010110: data <= 7'h00; 
        10'b0001010111: data <= 7'h00; 
        10'b0001011000: data <= 7'h00; 
        10'b0001011001: data <= 7'h00; 
        10'b0001011010: data <= 7'h00; 
        10'b0001011011: data <= 7'h00; 
        10'b0001011100: data <= 7'h00; 
        10'b0001011101: data <= 7'h00; 
        10'b0001011110: data <= 7'h00; 
        10'b0001011111: data <= 7'h00; 
        10'b0001100000: data <= 7'h00; 
        10'b0001100001: data <= 7'h00; 
        10'b0001100010: data <= 7'h00; 
        10'b0001100011: data <= 7'h00; 
        10'b0001100100: data <= 7'h00; 
        10'b0001100101: data <= 7'h00; 
        10'b0001100110: data <= 7'h00; 
        10'b0001100111: data <= 7'h00; 
        10'b0001101000: data <= 7'h00; 
        10'b0001101001: data <= 7'h00; 
        10'b0001101010: data <= 7'h00; 
        10'b0001101011: data <= 7'h00; 
        10'b0001101100: data <= 7'h00; 
        10'b0001101101: data <= 7'h00; 
        10'b0001101110: data <= 7'h00; 
        10'b0001101111: data <= 7'h00; 
        10'b0001110000: data <= 7'h00; 
        10'b0001110001: data <= 7'h00; 
        10'b0001110010: data <= 7'h00; 
        10'b0001110011: data <= 7'h00; 
        10'b0001110100: data <= 7'h00; 
        10'b0001110101: data <= 7'h00; 
        10'b0001110110: data <= 7'h00; 
        10'b0001110111: data <= 7'h00; 
        10'b0001111000: data <= 7'h00; 
        10'b0001111001: data <= 7'h00; 
        10'b0001111010: data <= 7'h00; 
        10'b0001111011: data <= 7'h00; 
        10'b0001111100: data <= 7'h7f; 
        10'b0001111101: data <= 7'h00; 
        10'b0001111110: data <= 7'h7f; 
        10'b0001111111: data <= 7'h00; 
        10'b0010000000: data <= 7'h00; 
        10'b0010000001: data <= 7'h00; 
        10'b0010000010: data <= 7'h00; 
        10'b0010000011: data <= 7'h00; 
        10'b0010000100: data <= 7'h00; 
        10'b0010000101: data <= 7'h00; 
        10'b0010000110: data <= 7'h00; 
        10'b0010000111: data <= 7'h00; 
        10'b0010001000: data <= 7'h00; 
        10'b0010001001: data <= 7'h00; 
        10'b0010001010: data <= 7'h00; 
        10'b0010001011: data <= 7'h00; 
        10'b0010001100: data <= 7'h00; 
        10'b0010001101: data <= 7'h00; 
        10'b0010001110: data <= 7'h00; 
        10'b0010001111: data <= 7'h00; 
        10'b0010010000: data <= 7'h00; 
        10'b0010010001: data <= 7'h00; 
        10'b0010010010: data <= 7'h00; 
        10'b0010010011: data <= 7'h00; 
        10'b0010010100: data <= 7'h00; 
        10'b0010010101: data <= 7'h00; 
        10'b0010010110: data <= 7'h00; 
        10'b0010010111: data <= 7'h00; 
        10'b0010011000: data <= 7'h00; 
        10'b0010011001: data <= 7'h00; 
        10'b0010011010: data <= 7'h00; 
        10'b0010011011: data <= 7'h00; 
        10'b0010011100: data <= 7'h00; 
        10'b0010011101: data <= 7'h00; 
        10'b0010011110: data <= 7'h00; 
        10'b0010011111: data <= 7'h00; 
        10'b0010100000: data <= 7'h00; 
        10'b0010100001: data <= 7'h00; 
        10'b0010100010: data <= 7'h00; 
        10'b0010100011: data <= 7'h00; 
        10'b0010100100: data <= 7'h00; 
        10'b0010100101: data <= 7'h00; 
        10'b0010100110: data <= 7'h00; 
        10'b0010100111: data <= 7'h00; 
        10'b0010101000: data <= 7'h00; 
        10'b0010101001: data <= 7'h00; 
        10'b0010101010: data <= 7'h00; 
        10'b0010101011: data <= 7'h00; 
        10'b0010101100: data <= 7'h00; 
        10'b0010101101: data <= 7'h00; 
        10'b0010101110: data <= 7'h00; 
        10'b0010101111: data <= 7'h00; 
        10'b0010110000: data <= 7'h00; 
        10'b0010110001: data <= 7'h00; 
        10'b0010110010: data <= 7'h00; 
        10'b0010110011: data <= 7'h00; 
        10'b0010110100: data <= 7'h7f; 
        10'b0010110101: data <= 7'h7f; 
        10'b0010110110: data <= 7'h7f; 
        10'b0010110111: data <= 7'h7f; 
        10'b0010111000: data <= 7'h7f; 
        10'b0010111001: data <= 7'h00; 
        10'b0010111010: data <= 7'h00; 
        10'b0010111011: data <= 7'h00; 
        10'b0010111100: data <= 7'h00; 
        10'b0010111101: data <= 7'h00; 
        10'b0010111110: data <= 7'h01; 
        10'b0010111111: data <= 7'h01; 
        10'b0011000000: data <= 7'h00; 
        10'b0011000001: data <= 7'h00; 
        10'b0011000010: data <= 7'h00; 
        10'b0011000011: data <= 7'h00; 
        10'b0011000100: data <= 7'h00; 
        10'b0011000101: data <= 7'h00; 
        10'b0011000110: data <= 7'h00; 
        10'b0011000111: data <= 7'h00; 
        10'b0011001000: data <= 7'h00; 
        10'b0011001001: data <= 7'h00; 
        10'b0011001010: data <= 7'h00; 
        10'b0011001011: data <= 7'h00; 
        10'b0011001100: data <= 7'h00; 
        10'b0011001101: data <= 7'h00; 
        10'b0011001110: data <= 7'h00; 
        10'b0011001111: data <= 7'h7f; 
        10'b0011010000: data <= 7'h7f; 
        10'b0011010001: data <= 7'h7f; 
        10'b0011010010: data <= 7'h7f; 
        10'b0011010011: data <= 7'h7f; 
        10'b0011010100: data <= 7'h7f; 
        10'b0011010101: data <= 7'h00; 
        10'b0011010110: data <= 7'h00; 
        10'b0011010111: data <= 7'h00; 
        10'b0011011000: data <= 7'h00; 
        10'b0011011001: data <= 7'h00; 
        10'b0011011010: data <= 7'h00; 
        10'b0011011011: data <= 7'h00; 
        10'b0011011100: data <= 7'h00; 
        10'b0011011101: data <= 7'h00; 
        10'b0011011110: data <= 7'h00; 
        10'b0011011111: data <= 7'h00; 
        10'b0011100000: data <= 7'h00; 
        10'b0011100001: data <= 7'h00; 
        10'b0011100010: data <= 7'h00; 
        10'b0011100011: data <= 7'h00; 
        10'b0011100100: data <= 7'h00; 
        10'b0011100101: data <= 7'h00; 
        10'b0011100110: data <= 7'h00; 
        10'b0011100111: data <= 7'h00; 
        10'b0011101000: data <= 7'h00; 
        10'b0011101001: data <= 7'h00; 
        10'b0011101010: data <= 7'h00; 
        10'b0011101011: data <= 7'h00; 
        10'b0011101100: data <= 7'h7f; 
        10'b0011101101: data <= 7'h00; 
        10'b0011101110: data <= 7'h7f; 
        10'b0011101111: data <= 7'h7f; 
        10'b0011110000: data <= 7'h7f; 
        10'b0011110001: data <= 7'h00; 
        10'b0011110010: data <= 7'h00; 
        10'b0011110011: data <= 7'h00; 
        10'b0011110100: data <= 7'h00; 
        10'b0011110101: data <= 7'h00; 
        10'b0011110110: data <= 7'h00; 
        10'b0011110111: data <= 7'h00; 
        10'b0011111000: data <= 7'h00; 
        10'b0011111001: data <= 7'h00; 
        10'b0011111010: data <= 7'h00; 
        10'b0011111011: data <= 7'h00; 
        10'b0011111100: data <= 7'h00; 
        10'b0011111101: data <= 7'h00; 
        10'b0011111110: data <= 7'h00; 
        10'b0011111111: data <= 7'h00; 
        10'b0100000000: data <= 7'h00; 
        10'b0100000001: data <= 7'h00; 
        10'b0100000010: data <= 7'h00; 
        10'b0100000011: data <= 7'h00; 
        10'b0100000100: data <= 7'h00; 
        10'b0100000101: data <= 7'h00; 
        10'b0100000110: data <= 7'h00; 
        10'b0100000111: data <= 7'h00; 
        10'b0100001000: data <= 7'h00; 
        10'b0100001001: data <= 7'h00; 
        10'b0100001010: data <= 7'h7f; 
        10'b0100001011: data <= 7'h7f; 
        10'b0100001100: data <= 7'h00; 
        10'b0100001101: data <= 7'h00; 
        10'b0100001110: data <= 7'h00; 
        10'b0100001111: data <= 7'h00; 
        10'b0100010000: data <= 7'h00; 
        10'b0100010001: data <= 7'h00; 
        10'b0100010010: data <= 7'h00; 
        10'b0100010011: data <= 7'h00; 
        10'b0100010100: data <= 7'h00; 
        10'b0100010101: data <= 7'h00; 
        10'b0100010110: data <= 7'h00; 
        10'b0100010111: data <= 7'h00; 
        10'b0100011000: data <= 7'h00; 
        10'b0100011001: data <= 7'h00; 
        10'b0100011010: data <= 7'h00; 
        10'b0100011011: data <= 7'h00; 
        10'b0100011100: data <= 7'h00; 
        10'b0100011101: data <= 7'h00; 
        10'b0100011110: data <= 7'h00; 
        10'b0100011111: data <= 7'h00; 
        10'b0100100000: data <= 7'h00; 
        10'b0100100001: data <= 7'h00; 
        10'b0100100010: data <= 7'h00; 
        10'b0100100011: data <= 7'h00; 
        10'b0100100100: data <= 7'h00; 
        10'b0100100101: data <= 7'h00; 
        10'b0100100110: data <= 7'h7f; 
        10'b0100100111: data <= 7'h00; 
        10'b0100101000: data <= 7'h00; 
        10'b0100101001: data <= 7'h00; 
        10'b0100101010: data <= 7'h00; 
        10'b0100101011: data <= 7'h00; 
        10'b0100101100: data <= 7'h00; 
        10'b0100101101: data <= 7'h00; 
        10'b0100101110: data <= 7'h00; 
        10'b0100101111: data <= 7'h00; 
        10'b0100110000: data <= 7'h00; 
        10'b0100110001: data <= 7'h00; 
        10'b0100110010: data <= 7'h00; 
        10'b0100110011: data <= 7'h00; 
        10'b0100110100: data <= 7'h00; 
        10'b0100110101: data <= 7'h00; 
        10'b0100110110: data <= 7'h00; 
        10'b0100110111: data <= 7'h00; 
        10'b0100111000: data <= 7'h00; 
        10'b0100111001: data <= 7'h00; 
        10'b0100111010: data <= 7'h00; 
        10'b0100111011: data <= 7'h00; 
        10'b0100111100: data <= 7'h00; 
        10'b0100111101: data <= 7'h00; 
        10'b0100111110: data <= 7'h01; 
        10'b0100111111: data <= 7'h00; 
        10'b0101000000: data <= 7'h00; 
        10'b0101000001: data <= 7'h7f; 
        10'b0101000010: data <= 7'h7f; 
        10'b0101000011: data <= 7'h00; 
        10'b0101000100: data <= 7'h00; 
        10'b0101000101: data <= 7'h00; 
        10'b0101000110: data <= 7'h00; 
        10'b0101000111: data <= 7'h00; 
        10'b0101001000: data <= 7'h00; 
        10'b0101001001: data <= 7'h00; 
        10'b0101001010: data <= 7'h00; 
        10'b0101001011: data <= 7'h00; 
        10'b0101001100: data <= 7'h00; 
        10'b0101001101: data <= 7'h00; 
        10'b0101001110: data <= 7'h00; 
        10'b0101001111: data <= 7'h00; 
        10'b0101010000: data <= 7'h00; 
        10'b0101010001: data <= 7'h00; 
        10'b0101010010: data <= 7'h00; 
        10'b0101010011: data <= 7'h00; 
        10'b0101010100: data <= 7'h00; 
        10'b0101010101: data <= 7'h00; 
        10'b0101010110: data <= 7'h00; 
        10'b0101010111: data <= 7'h00; 
        10'b0101011000: data <= 7'h01; 
        10'b0101011001: data <= 7'h01; 
        10'b0101011010: data <= 7'h01; 
        10'b0101011011: data <= 7'h01; 
        10'b0101011100: data <= 7'h01; 
        10'b0101011101: data <= 7'h00; 
        10'b0101011110: data <= 7'h00; 
        10'b0101011111: data <= 7'h00; 
        10'b0101100000: data <= 7'h01; 
        10'b0101100001: data <= 7'h00; 
        10'b0101100010: data <= 7'h00; 
        10'b0101100011: data <= 7'h00; 
        10'b0101100100: data <= 7'h00; 
        10'b0101100101: data <= 7'h00; 
        10'b0101100110: data <= 7'h00; 
        10'b0101100111: data <= 7'h00; 
        10'b0101101000: data <= 7'h00; 
        10'b0101101001: data <= 7'h00; 
        10'b0101101010: data <= 7'h00; 
        10'b0101101011: data <= 7'h00; 
        10'b0101101100: data <= 7'h00; 
        10'b0101101101: data <= 7'h00; 
        10'b0101101110: data <= 7'h00; 
        10'b0101101111: data <= 7'h00; 
        10'b0101110000: data <= 7'h00; 
        10'b0101110001: data <= 7'h00; 
        10'b0101110010: data <= 7'h01; 
        10'b0101110011: data <= 7'h01; 
        10'b0101110100: data <= 7'h01; 
        10'b0101110101: data <= 7'h01; 
        10'b0101110110: data <= 7'h01; 
        10'b0101110111: data <= 7'h01; 
        10'b0101111000: data <= 7'h01; 
        10'b0101111001: data <= 7'h00; 
        10'b0101111010: data <= 7'h00; 
        10'b0101111011: data <= 7'h00; 
        10'b0101111100: data <= 7'h00; 
        10'b0101111101: data <= 7'h01; 
        10'b0101111110: data <= 7'h00; 
        10'b0101111111: data <= 7'h00; 
        10'b0110000000: data <= 7'h00; 
        10'b0110000001: data <= 7'h00; 
        10'b0110000010: data <= 7'h00; 
        10'b0110000011: data <= 7'h00; 
        10'b0110000100: data <= 7'h00; 
        10'b0110000101: data <= 7'h00; 
        10'b0110000110: data <= 7'h00; 
        10'b0110000111: data <= 7'h00; 
        10'b0110001000: data <= 7'h00; 
        10'b0110001001: data <= 7'h00; 
        10'b0110001010: data <= 7'h00; 
        10'b0110001011: data <= 7'h00; 
        10'b0110001100: data <= 7'h00; 
        10'b0110001101: data <= 7'h01; 
        10'b0110001110: data <= 7'h01; 
        10'b0110001111: data <= 7'h01; 
        10'b0110010000: data <= 7'h01; 
        10'b0110010001: data <= 7'h01; 
        10'b0110010010: data <= 7'h01; 
        10'b0110010011: data <= 7'h01; 
        10'b0110010100: data <= 7'h01; 
        10'b0110010101: data <= 7'h00; 
        10'b0110010110: data <= 7'h00; 
        10'b0110010111: data <= 7'h00; 
        10'b0110011000: data <= 7'h01; 
        10'b0110011001: data <= 7'h01; 
        10'b0110011010: data <= 7'h01; 
        10'b0110011011: data <= 7'h01; 
        10'b0110011100: data <= 7'h00; 
        10'b0110011101: data <= 7'h00; 
        10'b0110011110: data <= 7'h00; 
        10'b0110011111: data <= 7'h00; 
        10'b0110100000: data <= 7'h00; 
        10'b0110100001: data <= 7'h00; 
        10'b0110100010: data <= 7'h00; 
        10'b0110100011: data <= 7'h00; 
        10'b0110100100: data <= 7'h00; 
        10'b0110100101: data <= 7'h00; 
        10'b0110100110: data <= 7'h00; 
        10'b0110100111: data <= 7'h00; 
        10'b0110101000: data <= 7'h00; 
        10'b0110101001: data <= 7'h00; 
        10'b0110101010: data <= 7'h00; 
        10'b0110101011: data <= 7'h00; 
        10'b0110101100: data <= 7'h01; 
        10'b0110101101: data <= 7'h01; 
        10'b0110101110: data <= 7'h00; 
        10'b0110101111: data <= 7'h00; 
        10'b0110110000: data <= 7'h00; 
        10'b0110110001: data <= 7'h00; 
        10'b0110110010: data <= 7'h00; 
        10'b0110110011: data <= 7'h00; 
        10'b0110110100: data <= 7'h01; 
        10'b0110110101: data <= 7'h01; 
        10'b0110110110: data <= 7'h00; 
        10'b0110110111: data <= 7'h00; 
        10'b0110111000: data <= 7'h00; 
        10'b0110111001: data <= 7'h00; 
        10'b0110111010: data <= 7'h00; 
        10'b0110111011: data <= 7'h00; 
        10'b0110111100: data <= 7'h00; 
        10'b0110111101: data <= 7'h00; 
        10'b0110111110: data <= 7'h00; 
        10'b0110111111: data <= 7'h00; 
        10'b0111000000: data <= 7'h00; 
        10'b0111000001: data <= 7'h00; 
        10'b0111000010: data <= 7'h00; 
        10'b0111000011: data <= 7'h00; 
        10'b0111000100: data <= 7'h00; 
        10'b0111000101: data <= 7'h00; 
        10'b0111000110: data <= 7'h00; 
        10'b0111000111: data <= 7'h00; 
        10'b0111001000: data <= 7'h01; 
        10'b0111001001: data <= 7'h00; 
        10'b0111001010: data <= 7'h00; 
        10'b0111001011: data <= 7'h00; 
        10'b0111001100: data <= 7'h00; 
        10'b0111001101: data <= 7'h00; 
        10'b0111001110: data <= 7'h01; 
        10'b0111001111: data <= 7'h01; 
        10'b0111010000: data <= 7'h01; 
        10'b0111010001: data <= 7'h01; 
        10'b0111010010: data <= 7'h00; 
        10'b0111010011: data <= 7'h00; 
        10'b0111010100: data <= 7'h00; 
        10'b0111010101: data <= 7'h00; 
        10'b0111010110: data <= 7'h00; 
        10'b0111010111: data <= 7'h00; 
        10'b0111011000: data <= 7'h00; 
        10'b0111011001: data <= 7'h00; 
        10'b0111011010: data <= 7'h00; 
        10'b0111011011: data <= 7'h00; 
        10'b0111011100: data <= 7'h00; 
        10'b0111011101: data <= 7'h00; 
        10'b0111011110: data <= 7'h00; 
        10'b0111011111: data <= 7'h00; 
        10'b0111100000: data <= 7'h00; 
        10'b0111100001: data <= 7'h00; 
        10'b0111100010: data <= 7'h00; 
        10'b0111100011: data <= 7'h00; 
        10'b0111100100: data <= 7'h01; 
        10'b0111100101: data <= 7'h01; 
        10'b0111100110: data <= 7'h00; 
        10'b0111100111: data <= 7'h00; 
        10'b0111101000: data <= 7'h00; 
        10'b0111101001: data <= 7'h01; 
        10'b0111101010: data <= 7'h01; 
        10'b0111101011: data <= 7'h01; 
        10'b0111101100: data <= 7'h01; 
        10'b0111101101: data <= 7'h00; 
        10'b0111101110: data <= 7'h00; 
        10'b0111101111: data <= 7'h00; 
        10'b0111110000: data <= 7'h00; 
        10'b0111110001: data <= 7'h00; 
        10'b0111110010: data <= 7'h00; 
        10'b0111110011: data <= 7'h00; 
        10'b0111110100: data <= 7'h00; 
        10'b0111110101: data <= 7'h00; 
        10'b0111110110: data <= 7'h00; 
        10'b0111110111: data <= 7'h00; 
        10'b0111111000: data <= 7'h00; 
        10'b0111111001: data <= 7'h00; 
        10'b0111111010: data <= 7'h00; 
        10'b0111111011: data <= 7'h00; 
        10'b0111111100: data <= 7'h00; 
        10'b0111111101: data <= 7'h00; 
        10'b0111111110: data <= 7'h00; 
        10'b0111111111: data <= 7'h00; 
        10'b1000000000: data <= 7'h00; 
        10'b1000000001: data <= 7'h00; 
        10'b1000000010: data <= 7'h00; 
        10'b1000000011: data <= 7'h00; 
        10'b1000000100: data <= 7'h00; 
        10'b1000000101: data <= 7'h00; 
        10'b1000000110: data <= 7'h00; 
        10'b1000000111: data <= 7'h00; 
        10'b1000001000: data <= 7'h00; 
        10'b1000001001: data <= 7'h00; 
        10'b1000001010: data <= 7'h00; 
        10'b1000001011: data <= 7'h00; 
        10'b1000001100: data <= 7'h00; 
        10'b1000001101: data <= 7'h00; 
        10'b1000001110: data <= 7'h00; 
        10'b1000001111: data <= 7'h00; 
        10'b1000010000: data <= 7'h00; 
        10'b1000010001: data <= 7'h00; 
        10'b1000010010: data <= 7'h00; 
        10'b1000010011: data <= 7'h00; 
        10'b1000010100: data <= 7'h00; 
        10'b1000010101: data <= 7'h00; 
        10'b1000010110: data <= 7'h00; 
        10'b1000010111: data <= 7'h00; 
        10'b1000011000: data <= 7'h00; 
        10'b1000011001: data <= 7'h00; 
        10'b1000011010: data <= 7'h00; 
        10'b1000011011: data <= 7'h00; 
        10'b1000011100: data <= 7'h7f; 
        10'b1000011101: data <= 7'h7f; 
        10'b1000011110: data <= 7'h7f; 
        10'b1000011111: data <= 7'h7f; 
        10'b1000100000: data <= 7'h7f; 
        10'b1000100001: data <= 7'h00; 
        10'b1000100010: data <= 7'h00; 
        10'b1000100011: data <= 7'h00; 
        10'b1000100100: data <= 7'h00; 
        10'b1000100101: data <= 7'h00; 
        10'b1000100110: data <= 7'h00; 
        10'b1000100111: data <= 7'h00; 
        10'b1000101000: data <= 7'h00; 
        10'b1000101001: data <= 7'h00; 
        10'b1000101010: data <= 7'h00; 
        10'b1000101011: data <= 7'h00; 
        10'b1000101100: data <= 7'h00; 
        10'b1000101101: data <= 7'h00; 
        10'b1000101110: data <= 7'h00; 
        10'b1000101111: data <= 7'h00; 
        10'b1000110000: data <= 7'h00; 
        10'b1000110001: data <= 7'h00; 
        10'b1000110010: data <= 7'h00; 
        10'b1000110011: data <= 7'h00; 
        10'b1000110100: data <= 7'h00; 
        10'b1000110101: data <= 7'h00; 
        10'b1000110110: data <= 7'h00; 
        10'b1000110111: data <= 7'h7f; 
        10'b1000111000: data <= 7'h7f; 
        10'b1000111001: data <= 7'h7f; 
        10'b1000111010: data <= 7'h7f; 
        10'b1000111011: data <= 7'h7f; 
        10'b1000111100: data <= 7'h00; 
        10'b1000111101: data <= 7'h7f; 
        10'b1000111110: data <= 7'h00; 
        10'b1000111111: data <= 7'h00; 
        10'b1001000000: data <= 7'h00; 
        10'b1001000001: data <= 7'h00; 
        10'b1001000010: data <= 7'h00; 
        10'b1001000011: data <= 7'h00; 
        10'b1001000100: data <= 7'h00; 
        10'b1001000101: data <= 7'h00; 
        10'b1001000110: data <= 7'h00; 
        10'b1001000111: data <= 7'h00; 
        10'b1001001000: data <= 7'h00; 
        10'b1001001001: data <= 7'h00; 
        10'b1001001010: data <= 7'h00; 
        10'b1001001011: data <= 7'h00; 
        10'b1001001100: data <= 7'h00; 
        10'b1001001101: data <= 7'h00; 
        10'b1001001110: data <= 7'h00; 
        10'b1001001111: data <= 7'h00; 
        10'b1001010000: data <= 7'h00; 
        10'b1001010001: data <= 7'h00; 
        10'b1001010010: data <= 7'h00; 
        10'b1001010011: data <= 7'h7f; 
        10'b1001010100: data <= 7'h00; 
        10'b1001010101: data <= 7'h7f; 
        10'b1001010110: data <= 7'h00; 
        10'b1001010111: data <= 7'h00; 
        10'b1001011000: data <= 7'h00; 
        10'b1001011001: data <= 7'h00; 
        10'b1001011010: data <= 7'h00; 
        10'b1001011011: data <= 7'h00; 
        10'b1001011100: data <= 7'h00; 
        10'b1001011101: data <= 7'h00; 
        10'b1001011110: data <= 7'h00; 
        10'b1001011111: data <= 7'h00; 
        10'b1001100000: data <= 7'h00; 
        10'b1001100001: data <= 7'h00; 
        10'b1001100010: data <= 7'h00; 
        10'b1001100011: data <= 7'h00; 
        10'b1001100100: data <= 7'h00; 
        10'b1001100101: data <= 7'h00; 
        10'b1001100110: data <= 7'h00; 
        10'b1001100111: data <= 7'h00; 
        10'b1001101000: data <= 7'h00; 
        10'b1001101001: data <= 7'h00; 
        10'b1001101010: data <= 7'h00; 
        10'b1001101011: data <= 7'h00; 
        10'b1001101100: data <= 7'h00; 
        10'b1001101101: data <= 7'h00; 
        10'b1001101110: data <= 7'h00; 
        10'b1001101111: data <= 7'h00; 
        10'b1001110000: data <= 7'h00; 
        10'b1001110001: data <= 7'h00; 
        10'b1001110010: data <= 7'h00; 
        10'b1001110011: data <= 7'h00; 
        10'b1001110100: data <= 7'h00; 
        10'b1001110101: data <= 7'h00; 
        10'b1001110110: data <= 7'h00; 
        10'b1001110111: data <= 7'h00; 
        10'b1001111000: data <= 7'h00; 
        10'b1001111001: data <= 7'h00; 
        10'b1001111010: data <= 7'h00; 
        10'b1001111011: data <= 7'h00; 
        10'b1001111100: data <= 7'h00; 
        10'b1001111101: data <= 7'h00; 
        10'b1001111110: data <= 7'h00; 
        10'b1001111111: data <= 7'h00; 
        10'b1010000000: data <= 7'h00; 
        10'b1010000001: data <= 7'h00; 
        10'b1010000010: data <= 7'h00; 
        10'b1010000011: data <= 7'h00; 
        10'b1010000100: data <= 7'h00; 
        10'b1010000101: data <= 7'h00; 
        10'b1010000110: data <= 7'h00; 
        10'b1010000111: data <= 7'h00; 
        10'b1010001000: data <= 7'h00; 
        10'b1010001001: data <= 7'h00; 
        10'b1010001010: data <= 7'h00; 
        10'b1010001011: data <= 7'h00; 
        10'b1010001100: data <= 7'h00; 
        10'b1010001101: data <= 7'h00; 
        10'b1010001110: data <= 7'h00; 
        10'b1010001111: data <= 7'h00; 
        10'b1010010000: data <= 7'h00; 
        10'b1010010001: data <= 7'h00; 
        10'b1010010010: data <= 7'h00; 
        10'b1010010011: data <= 7'h00; 
        10'b1010010100: data <= 7'h00; 
        10'b1010010101: data <= 7'h00; 
        10'b1010010110: data <= 7'h00; 
        10'b1010010111: data <= 7'h00; 
        10'b1010011000: data <= 7'h00; 
        10'b1010011001: data <= 7'h00; 
        10'b1010011010: data <= 7'h00; 
        10'b1010011011: data <= 7'h00; 
        10'b1010011100: data <= 7'h00; 
        10'b1010011101: data <= 7'h00; 
        10'b1010011110: data <= 7'h00; 
        10'b1010011111: data <= 7'h00; 
        10'b1010100000: data <= 7'h00; 
        10'b1010100001: data <= 7'h00; 
        10'b1010100010: data <= 7'h00; 
        10'b1010100011: data <= 7'h00; 
        10'b1010100100: data <= 7'h00; 
        10'b1010100101: data <= 7'h00; 
        10'b1010100110: data <= 7'h00; 
        10'b1010100111: data <= 7'h00; 
        10'b1010101000: data <= 7'h00; 
        10'b1010101001: data <= 7'h00; 
        10'b1010101010: data <= 7'h00; 
        10'b1010101011: data <= 7'h00; 
        10'b1010101100: data <= 7'h00; 
        10'b1010101101: data <= 7'h00; 
        10'b1010101110: data <= 7'h00; 
        10'b1010101111: data <= 7'h00; 
        10'b1010110000: data <= 7'h00; 
        10'b1010110001: data <= 7'h00; 
        10'b1010110010: data <= 7'h00; 
        10'b1010110011: data <= 7'h00; 
        10'b1010110100: data <= 7'h00; 
        10'b1010110101: data <= 7'h00; 
        10'b1010110110: data <= 7'h00; 
        10'b1010110111: data <= 7'h00; 
        10'b1010111000: data <= 7'h00; 
        10'b1010111001: data <= 7'h00; 
        10'b1010111010: data <= 7'h00; 
        10'b1010111011: data <= 7'h00; 
        10'b1010111100: data <= 7'h00; 
        10'b1010111101: data <= 7'h00; 
        10'b1010111110: data <= 7'h00; 
        10'b1010111111: data <= 7'h00; 
        10'b1011000000: data <= 7'h00; 
        10'b1011000001: data <= 7'h00; 
        10'b1011000010: data <= 7'h00; 
        10'b1011000011: data <= 7'h00; 
        10'b1011000100: data <= 7'h00; 
        10'b1011000101: data <= 7'h00; 
        10'b1011000110: data <= 7'h00; 
        10'b1011000111: data <= 7'h00; 
        10'b1011001000: data <= 7'h00; 
        10'b1011001001: data <= 7'h00; 
        10'b1011001010: data <= 7'h00; 
        10'b1011001011: data <= 7'h00; 
        10'b1011001100: data <= 7'h00; 
        10'b1011001101: data <= 7'h00; 
        10'b1011001110: data <= 7'h00; 
        10'b1011001111: data <= 7'h00; 
        10'b1011010000: data <= 7'h00; 
        10'b1011010001: data <= 7'h00; 
        10'b1011010010: data <= 7'h00; 
        10'b1011010011: data <= 7'h00; 
        10'b1011010100: data <= 7'h00; 
        10'b1011010101: data <= 7'h00; 
        10'b1011010110: data <= 7'h00; 
        10'b1011010111: data <= 7'h00; 
        10'b1011011000: data <= 7'h00; 
        10'b1011011001: data <= 7'h00; 
        10'b1011011010: data <= 7'h00; 
        10'b1011011011: data <= 7'h00; 
        10'b1011011100: data <= 7'h00; 
        10'b1011011101: data <= 7'h00; 
        10'b1011011110: data <= 7'h00; 
        10'b1011011111: data <= 7'h00; 
        10'b1011100000: data <= 7'h00; 
        10'b1011100001: data <= 7'h00; 
        10'b1011100010: data <= 7'h00; 
        10'b1011100011: data <= 7'h00; 
        10'b1011100100: data <= 7'h00; 
        10'b1011100101: data <= 7'h00; 
        10'b1011100110: data <= 7'h00; 
        10'b1011100111: data <= 7'h00; 
        10'b1011101000: data <= 7'h00; 
        10'b1011101001: data <= 7'h00; 
        10'b1011101010: data <= 7'h00; 
        10'b1011101011: data <= 7'h00; 
        10'b1011101100: data <= 7'h00; 
        10'b1011101101: data <= 7'h00; 
        10'b1011101110: data <= 7'h00; 
        10'b1011101111: data <= 7'h00; 
        10'b1011110000: data <= 7'h00; 
        10'b1011110001: data <= 7'h00; 
        10'b1011110010: data <= 7'h00; 
        10'b1011110011: data <= 7'h00; 
        10'b1011110100: data <= 7'h00; 
        10'b1011110101: data <= 7'h00; 
        10'b1011110110: data <= 7'h00; 
        10'b1011110111: data <= 7'h00; 
        10'b1011111000: data <= 7'h00; 
        10'b1011111001: data <= 7'h00; 
        10'b1011111010: data <= 7'h00; 
        10'b1011111011: data <= 7'h00; 
        10'b1011111100: data <= 7'h00; 
        10'b1011111101: data <= 7'h00; 
        10'b1011111110: data <= 7'h00; 
        10'b1011111111: data <= 7'h00; 
        10'b1100000000: data <= 7'h00; 
        10'b1100000001: data <= 7'h00; 
        10'b1100000010: data <= 7'h00; 
        10'b1100000011: data <= 7'h00; 
        10'b1100000100: data <= 7'h00; 
        10'b1100000101: data <= 7'h00; 
        10'b1100000110: data <= 7'h00; 
        10'b1100000111: data <= 7'h00; 
        10'b1100001000: data <= 7'h00; 
        10'b1100001001: data <= 7'h00; 
        10'b1100001010: data <= 7'h00; 
        10'b1100001011: data <= 7'h00; 
        10'b1100001100: data <= 7'h00; 
        10'b1100001101: data <= 7'h00; 
        10'b1100001110: data <= 7'h00; 
        10'b1100001111: data <= 7'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 2) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 8'h00; 
        10'b0000000001: data <= 8'h00; 
        10'b0000000010: data <= 8'h00; 
        10'b0000000011: data <= 8'h00; 
        10'b0000000100: data <= 8'h00; 
        10'b0000000101: data <= 8'h00; 
        10'b0000000110: data <= 8'h00; 
        10'b0000000111: data <= 8'h00; 
        10'b0000001000: data <= 8'h00; 
        10'b0000001001: data <= 8'h00; 
        10'b0000001010: data <= 8'h00; 
        10'b0000001011: data <= 8'h00; 
        10'b0000001100: data <= 8'h00; 
        10'b0000001101: data <= 8'h00; 
        10'b0000001110: data <= 8'h00; 
        10'b0000001111: data <= 8'h00; 
        10'b0000010000: data <= 8'h00; 
        10'b0000010001: data <= 8'h00; 
        10'b0000010010: data <= 8'h00; 
        10'b0000010011: data <= 8'h00; 
        10'b0000010100: data <= 8'h00; 
        10'b0000010101: data <= 8'h00; 
        10'b0000010110: data <= 8'h00; 
        10'b0000010111: data <= 8'h00; 
        10'b0000011000: data <= 8'h00; 
        10'b0000011001: data <= 8'h00; 
        10'b0000011010: data <= 8'h00; 
        10'b0000011011: data <= 8'h00; 
        10'b0000011100: data <= 8'h00; 
        10'b0000011101: data <= 8'h00; 
        10'b0000011110: data <= 8'h00; 
        10'b0000011111: data <= 8'h00; 
        10'b0000100000: data <= 8'h00; 
        10'b0000100001: data <= 8'h00; 
        10'b0000100010: data <= 8'h00; 
        10'b0000100011: data <= 8'h00; 
        10'b0000100100: data <= 8'h00; 
        10'b0000100101: data <= 8'h00; 
        10'b0000100110: data <= 8'h00; 
        10'b0000100111: data <= 8'h00; 
        10'b0000101000: data <= 8'h00; 
        10'b0000101001: data <= 8'h00; 
        10'b0000101010: data <= 8'h00; 
        10'b0000101011: data <= 8'h00; 
        10'b0000101100: data <= 8'h00; 
        10'b0000101101: data <= 8'h00; 
        10'b0000101110: data <= 8'h00; 
        10'b0000101111: data <= 8'h00; 
        10'b0000110000: data <= 8'h00; 
        10'b0000110001: data <= 8'h00; 
        10'b0000110010: data <= 8'h00; 
        10'b0000110011: data <= 8'h00; 
        10'b0000110100: data <= 8'h00; 
        10'b0000110101: data <= 8'h00; 
        10'b0000110110: data <= 8'h00; 
        10'b0000110111: data <= 8'h00; 
        10'b0000111000: data <= 8'h00; 
        10'b0000111001: data <= 8'h00; 
        10'b0000111010: data <= 8'h00; 
        10'b0000111011: data <= 8'h00; 
        10'b0000111100: data <= 8'h00; 
        10'b0000111101: data <= 8'h00; 
        10'b0000111110: data <= 8'h00; 
        10'b0000111111: data <= 8'h00; 
        10'b0001000000: data <= 8'h00; 
        10'b0001000001: data <= 8'h00; 
        10'b0001000010: data <= 8'h00; 
        10'b0001000011: data <= 8'h00; 
        10'b0001000100: data <= 8'hff; 
        10'b0001000101: data <= 8'h00; 
        10'b0001000110: data <= 8'h00; 
        10'b0001000111: data <= 8'h00; 
        10'b0001001000: data <= 8'h00; 
        10'b0001001001: data <= 8'h00; 
        10'b0001001010: data <= 8'h00; 
        10'b0001001011: data <= 8'h00; 
        10'b0001001100: data <= 8'h00; 
        10'b0001001101: data <= 8'h00; 
        10'b0001001110: data <= 8'h00; 
        10'b0001001111: data <= 8'h00; 
        10'b0001010000: data <= 8'h00; 
        10'b0001010001: data <= 8'h00; 
        10'b0001010010: data <= 8'h00; 
        10'b0001010011: data <= 8'h00; 
        10'b0001010100: data <= 8'h00; 
        10'b0001010101: data <= 8'h00; 
        10'b0001010110: data <= 8'h00; 
        10'b0001010111: data <= 8'h00; 
        10'b0001011000: data <= 8'h00; 
        10'b0001011001: data <= 8'h00; 
        10'b0001011010: data <= 8'h00; 
        10'b0001011011: data <= 8'h00; 
        10'b0001011100: data <= 8'h00; 
        10'b0001011101: data <= 8'h00; 
        10'b0001011110: data <= 8'h00; 
        10'b0001011111: data <= 8'hff; 
        10'b0001100000: data <= 8'hff; 
        10'b0001100001: data <= 8'hff; 
        10'b0001100010: data <= 8'hff; 
        10'b0001100011: data <= 8'hff; 
        10'b0001100100: data <= 8'hff; 
        10'b0001100101: data <= 8'h00; 
        10'b0001100110: data <= 8'h00; 
        10'b0001100111: data <= 8'h00; 
        10'b0001101000: data <= 8'h00; 
        10'b0001101001: data <= 8'h00; 
        10'b0001101010: data <= 8'h00; 
        10'b0001101011: data <= 8'h00; 
        10'b0001101100: data <= 8'h00; 
        10'b0001101101: data <= 8'h00; 
        10'b0001101110: data <= 8'h00; 
        10'b0001101111: data <= 8'h00; 
        10'b0001110000: data <= 8'h00; 
        10'b0001110001: data <= 8'h00; 
        10'b0001110010: data <= 8'h00; 
        10'b0001110011: data <= 8'h00; 
        10'b0001110100: data <= 8'h00; 
        10'b0001110101: data <= 8'h00; 
        10'b0001110110: data <= 8'h00; 
        10'b0001110111: data <= 8'h00; 
        10'b0001111000: data <= 8'h00; 
        10'b0001111001: data <= 8'h00; 
        10'b0001111010: data <= 8'hff; 
        10'b0001111011: data <= 8'hff; 
        10'b0001111100: data <= 8'hff; 
        10'b0001111101: data <= 8'hff; 
        10'b0001111110: data <= 8'hff; 
        10'b0001111111: data <= 8'hff; 
        10'b0010000000: data <= 8'h00; 
        10'b0010000001: data <= 8'h00; 
        10'b0010000010: data <= 8'h00; 
        10'b0010000011: data <= 8'h00; 
        10'b0010000100: data <= 8'h00; 
        10'b0010000101: data <= 8'h00; 
        10'b0010000110: data <= 8'h00; 
        10'b0010000111: data <= 8'h00; 
        10'b0010001000: data <= 8'h00; 
        10'b0010001001: data <= 8'h00; 
        10'b0010001010: data <= 8'h00; 
        10'b0010001011: data <= 8'h00; 
        10'b0010001100: data <= 8'h00; 
        10'b0010001101: data <= 8'h00; 
        10'b0010001110: data <= 8'h00; 
        10'b0010001111: data <= 8'h00; 
        10'b0010010000: data <= 8'h00; 
        10'b0010010001: data <= 8'h00; 
        10'b0010010010: data <= 8'h00; 
        10'b0010010011: data <= 8'h00; 
        10'b0010010100: data <= 8'h00; 
        10'b0010010101: data <= 8'h00; 
        10'b0010010110: data <= 8'hff; 
        10'b0010010111: data <= 8'h00; 
        10'b0010011000: data <= 8'hff; 
        10'b0010011001: data <= 8'hff; 
        10'b0010011010: data <= 8'hff; 
        10'b0010011011: data <= 8'h00; 
        10'b0010011100: data <= 8'h00; 
        10'b0010011101: data <= 8'h00; 
        10'b0010011110: data <= 8'h00; 
        10'b0010011111: data <= 8'h00; 
        10'b0010100000: data <= 8'h00; 
        10'b0010100001: data <= 8'h00; 
        10'b0010100010: data <= 8'h01; 
        10'b0010100011: data <= 8'h01; 
        10'b0010100100: data <= 8'h00; 
        10'b0010100101: data <= 8'h00; 
        10'b0010100110: data <= 8'h00; 
        10'b0010100111: data <= 8'h00; 
        10'b0010101000: data <= 8'h00; 
        10'b0010101001: data <= 8'h00; 
        10'b0010101010: data <= 8'h00; 
        10'b0010101011: data <= 8'h00; 
        10'b0010101100: data <= 8'h00; 
        10'b0010101101: data <= 8'h00; 
        10'b0010101110: data <= 8'h00; 
        10'b0010101111: data <= 8'h00; 
        10'b0010110000: data <= 8'h00; 
        10'b0010110001: data <= 8'h00; 
        10'b0010110010: data <= 8'h00; 
        10'b0010110011: data <= 8'hff; 
        10'b0010110100: data <= 8'hff; 
        10'b0010110101: data <= 8'hff; 
        10'b0010110110: data <= 8'hff; 
        10'b0010110111: data <= 8'hff; 
        10'b0010111000: data <= 8'hff; 
        10'b0010111001: data <= 8'hff; 
        10'b0010111010: data <= 8'hff; 
        10'b0010111011: data <= 8'h00; 
        10'b0010111100: data <= 8'h00; 
        10'b0010111101: data <= 8'h00; 
        10'b0010111110: data <= 8'h01; 
        10'b0010111111: data <= 8'h01; 
        10'b0011000000: data <= 8'h00; 
        10'b0011000001: data <= 8'h00; 
        10'b0011000010: data <= 8'h00; 
        10'b0011000011: data <= 8'h00; 
        10'b0011000100: data <= 8'h00; 
        10'b0011000101: data <= 8'h00; 
        10'b0011000110: data <= 8'h00; 
        10'b0011000111: data <= 8'h00; 
        10'b0011001000: data <= 8'h00; 
        10'b0011001001: data <= 8'h00; 
        10'b0011001010: data <= 8'h00; 
        10'b0011001011: data <= 8'h00; 
        10'b0011001100: data <= 8'h00; 
        10'b0011001101: data <= 8'h00; 
        10'b0011001110: data <= 8'hff; 
        10'b0011001111: data <= 8'hff; 
        10'b0011010000: data <= 8'hfe; 
        10'b0011010001: data <= 8'hff; 
        10'b0011010010: data <= 8'hff; 
        10'b0011010011: data <= 8'hff; 
        10'b0011010100: data <= 8'hff; 
        10'b0011010101: data <= 8'hff; 
        10'b0011010110: data <= 8'hff; 
        10'b0011010111: data <= 8'hff; 
        10'b0011011000: data <= 8'hff; 
        10'b0011011001: data <= 8'h00; 
        10'b0011011010: data <= 8'h01; 
        10'b0011011011: data <= 8'h01; 
        10'b0011011100: data <= 8'h00; 
        10'b0011011101: data <= 8'h00; 
        10'b0011011110: data <= 8'h00; 
        10'b0011011111: data <= 8'h00; 
        10'b0011100000: data <= 8'h00; 
        10'b0011100001: data <= 8'h00; 
        10'b0011100010: data <= 8'h00; 
        10'b0011100011: data <= 8'h00; 
        10'b0011100100: data <= 8'h00; 
        10'b0011100101: data <= 8'h00; 
        10'b0011100110: data <= 8'h00; 
        10'b0011100111: data <= 8'h00; 
        10'b0011101000: data <= 8'hff; 
        10'b0011101001: data <= 8'h00; 
        10'b0011101010: data <= 8'h00; 
        10'b0011101011: data <= 8'hff; 
        10'b0011101100: data <= 8'hff; 
        10'b0011101101: data <= 8'hff; 
        10'b0011101110: data <= 8'hfe; 
        10'b0011101111: data <= 8'hfe; 
        10'b0011110000: data <= 8'hff; 
        10'b0011110001: data <= 8'hff; 
        10'b0011110010: data <= 8'hff; 
        10'b0011110011: data <= 8'h00; 
        10'b0011110100: data <= 8'h00; 
        10'b0011110101: data <= 8'h00; 
        10'b0011110110: data <= 8'h00; 
        10'b0011110111: data <= 8'h00; 
        10'b0011111000: data <= 8'h00; 
        10'b0011111001: data <= 8'h00; 
        10'b0011111010: data <= 8'h00; 
        10'b0011111011: data <= 8'h00; 
        10'b0011111100: data <= 8'h00; 
        10'b0011111101: data <= 8'h00; 
        10'b0011111110: data <= 8'h00; 
        10'b0011111111: data <= 8'h00; 
        10'b0100000000: data <= 8'h00; 
        10'b0100000001: data <= 8'h00; 
        10'b0100000010: data <= 8'h00; 
        10'b0100000011: data <= 8'h00; 
        10'b0100000100: data <= 8'h00; 
        10'b0100000101: data <= 8'h00; 
        10'b0100000110: data <= 8'h00; 
        10'b0100000111: data <= 8'h00; 
        10'b0100001000: data <= 8'h00; 
        10'b0100001001: data <= 8'hff; 
        10'b0100001010: data <= 8'hfe; 
        10'b0100001011: data <= 8'hfe; 
        10'b0100001100: data <= 8'h00; 
        10'b0100001101: data <= 8'h00; 
        10'b0100001110: data <= 8'h00; 
        10'b0100001111: data <= 8'h00; 
        10'b0100010000: data <= 8'h00; 
        10'b0100010001: data <= 8'h00; 
        10'b0100010010: data <= 8'h00; 
        10'b0100010011: data <= 8'h00; 
        10'b0100010100: data <= 8'h00; 
        10'b0100010101: data <= 8'h00; 
        10'b0100010110: data <= 8'h00; 
        10'b0100010111: data <= 8'h00; 
        10'b0100011000: data <= 8'h00; 
        10'b0100011001: data <= 8'h00; 
        10'b0100011010: data <= 8'h00; 
        10'b0100011011: data <= 8'h00; 
        10'b0100011100: data <= 8'h00; 
        10'b0100011101: data <= 8'h00; 
        10'b0100011110: data <= 8'hff; 
        10'b0100011111: data <= 8'h00; 
        10'b0100100000: data <= 8'h00; 
        10'b0100100001: data <= 8'h01; 
        10'b0100100010: data <= 8'h00; 
        10'b0100100011: data <= 8'h00; 
        10'b0100100100: data <= 8'h00; 
        10'b0100100101: data <= 8'hff; 
        10'b0100100110: data <= 8'hfd; 
        10'b0100100111: data <= 8'hff; 
        10'b0100101000: data <= 8'h00; 
        10'b0100101001: data <= 8'h00; 
        10'b0100101010: data <= 8'h00; 
        10'b0100101011: data <= 8'h00; 
        10'b0100101100: data <= 8'h00; 
        10'b0100101101: data <= 8'h00; 
        10'b0100101110: data <= 8'h00; 
        10'b0100101111: data <= 8'hff; 
        10'b0100110000: data <= 8'h00; 
        10'b0100110001: data <= 8'h00; 
        10'b0100110010: data <= 8'h00; 
        10'b0100110011: data <= 8'h00; 
        10'b0100110100: data <= 8'h00; 
        10'b0100110101: data <= 8'h00; 
        10'b0100110110: data <= 8'h00; 
        10'b0100110111: data <= 8'h00; 
        10'b0100111000: data <= 8'h00; 
        10'b0100111001: data <= 8'h00; 
        10'b0100111010: data <= 8'h00; 
        10'b0100111011: data <= 8'h00; 
        10'b0100111100: data <= 8'h01; 
        10'b0100111101: data <= 8'h01; 
        10'b0100111110: data <= 8'h01; 
        10'b0100111111: data <= 8'h01; 
        10'b0101000000: data <= 8'h01; 
        10'b0101000001: data <= 8'hff; 
        10'b0101000010: data <= 8'hfe; 
        10'b0101000011: data <= 8'h00; 
        10'b0101000100: data <= 8'h01; 
        10'b0101000101: data <= 8'h00; 
        10'b0101000110: data <= 8'h00; 
        10'b0101000111: data <= 8'h00; 
        10'b0101001000: data <= 8'hff; 
        10'b0101001001: data <= 8'h00; 
        10'b0101001010: data <= 8'h00; 
        10'b0101001011: data <= 8'h00; 
        10'b0101001100: data <= 8'h00; 
        10'b0101001101: data <= 8'h00; 
        10'b0101001110: data <= 8'h00; 
        10'b0101001111: data <= 8'h00; 
        10'b0101010000: data <= 8'h00; 
        10'b0101010001: data <= 8'h00; 
        10'b0101010010: data <= 8'h00; 
        10'b0101010011: data <= 8'h00; 
        10'b0101010100: data <= 8'h00; 
        10'b0101010101: data <= 8'h00; 
        10'b0101010110: data <= 8'h01; 
        10'b0101010111: data <= 8'h01; 
        10'b0101011000: data <= 8'h01; 
        10'b0101011001: data <= 8'h01; 
        10'b0101011010: data <= 8'h02; 
        10'b0101011011: data <= 8'h02; 
        10'b0101011100: data <= 8'h02; 
        10'b0101011101: data <= 8'h00; 
        10'b0101011110: data <= 8'hff; 
        10'b0101011111: data <= 8'h01; 
        10'b0101100000: data <= 8'h01; 
        10'b0101100001: data <= 8'h00; 
        10'b0101100010: data <= 8'h00; 
        10'b0101100011: data <= 8'h00; 
        10'b0101100100: data <= 8'h00; 
        10'b0101100101: data <= 8'h00; 
        10'b0101100110: data <= 8'h00; 
        10'b0101100111: data <= 8'h00; 
        10'b0101101000: data <= 8'h00; 
        10'b0101101001: data <= 8'h00; 
        10'b0101101010: data <= 8'h00; 
        10'b0101101011: data <= 8'h00; 
        10'b0101101100: data <= 8'h00; 
        10'b0101101101: data <= 8'h00; 
        10'b0101101110: data <= 8'h00; 
        10'b0101101111: data <= 8'h00; 
        10'b0101110000: data <= 8'h00; 
        10'b0101110001: data <= 8'h01; 
        10'b0101110010: data <= 8'h01; 
        10'b0101110011: data <= 8'h01; 
        10'b0101110100: data <= 8'h02; 
        10'b0101110101: data <= 8'h01; 
        10'b0101110110: data <= 8'h02; 
        10'b0101110111: data <= 8'h03; 
        10'b0101111000: data <= 8'h02; 
        10'b0101111001: data <= 8'h00; 
        10'b0101111010: data <= 8'h00; 
        10'b0101111011: data <= 8'h01; 
        10'b0101111100: data <= 8'h01; 
        10'b0101111101: data <= 8'h01; 
        10'b0101111110: data <= 8'h01; 
        10'b0101111111: data <= 8'h00; 
        10'b0110000000: data <= 8'h01; 
        10'b0110000001: data <= 8'h01; 
        10'b0110000010: data <= 8'h00; 
        10'b0110000011: data <= 8'h00; 
        10'b0110000100: data <= 8'h00; 
        10'b0110000101: data <= 8'h00; 
        10'b0110000110: data <= 8'h00; 
        10'b0110000111: data <= 8'h00; 
        10'b0110001000: data <= 8'h00; 
        10'b0110001001: data <= 8'h00; 
        10'b0110001010: data <= 8'h00; 
        10'b0110001011: data <= 8'h00; 
        10'b0110001100: data <= 8'h01; 
        10'b0110001101: data <= 8'h01; 
        10'b0110001110: data <= 8'h01; 
        10'b0110001111: data <= 8'h02; 
        10'b0110010000: data <= 8'h01; 
        10'b0110010001: data <= 8'h01; 
        10'b0110010010: data <= 8'h01; 
        10'b0110010011: data <= 8'h02; 
        10'b0110010100: data <= 8'h01; 
        10'b0110010101: data <= 8'h00; 
        10'b0110010110: data <= 8'h00; 
        10'b0110010111: data <= 8'h00; 
        10'b0110011000: data <= 8'h01; 
        10'b0110011001: data <= 8'h02; 
        10'b0110011010: data <= 8'h01; 
        10'b0110011011: data <= 8'h01; 
        10'b0110011100: data <= 8'h01; 
        10'b0110011101: data <= 8'h00; 
        10'b0110011110: data <= 8'h00; 
        10'b0110011111: data <= 8'h00; 
        10'b0110100000: data <= 8'h00; 
        10'b0110100001: data <= 8'h00; 
        10'b0110100010: data <= 8'h00; 
        10'b0110100011: data <= 8'h00; 
        10'b0110100100: data <= 8'h00; 
        10'b0110100101: data <= 8'h00; 
        10'b0110100110: data <= 8'h00; 
        10'b0110100111: data <= 8'h00; 
        10'b0110101000: data <= 8'h00; 
        10'b0110101001: data <= 8'h01; 
        10'b0110101010: data <= 8'h01; 
        10'b0110101011: data <= 8'h01; 
        10'b0110101100: data <= 8'h01; 
        10'b0110101101: data <= 8'h01; 
        10'b0110101110: data <= 8'h01; 
        10'b0110101111: data <= 8'h01; 
        10'b0110110000: data <= 8'h01; 
        10'b0110110001: data <= 8'h00; 
        10'b0110110010: data <= 8'h01; 
        10'b0110110011: data <= 8'h01; 
        10'b0110110100: data <= 8'h02; 
        10'b0110110101: data <= 8'h01; 
        10'b0110110110: data <= 8'h01; 
        10'b0110110111: data <= 8'h01; 
        10'b0110111000: data <= 8'h00; 
        10'b0110111001: data <= 8'h00; 
        10'b0110111010: data <= 8'h00; 
        10'b0110111011: data <= 8'h00; 
        10'b0110111100: data <= 8'h00; 
        10'b0110111101: data <= 8'h00; 
        10'b0110111110: data <= 8'h00; 
        10'b0110111111: data <= 8'h00; 
        10'b0111000000: data <= 8'h00; 
        10'b0111000001: data <= 8'h00; 
        10'b0111000010: data <= 8'h00; 
        10'b0111000011: data <= 8'h00; 
        10'b0111000100: data <= 8'h00; 
        10'b0111000101: data <= 8'h00; 
        10'b0111000110: data <= 8'h01; 
        10'b0111000111: data <= 8'h01; 
        10'b0111001000: data <= 8'h01; 
        10'b0111001001: data <= 8'h01; 
        10'b0111001010: data <= 8'h00; 
        10'b0111001011: data <= 8'h00; 
        10'b0111001100: data <= 8'h00; 
        10'b0111001101: data <= 8'h00; 
        10'b0111001110: data <= 8'h01; 
        10'b0111001111: data <= 8'h02; 
        10'b0111010000: data <= 8'h02; 
        10'b0111010001: data <= 8'h01; 
        10'b0111010010: data <= 8'h01; 
        10'b0111010011: data <= 8'h00; 
        10'b0111010100: data <= 8'h00; 
        10'b0111010101: data <= 8'h01; 
        10'b0111010110: data <= 8'h00; 
        10'b0111010111: data <= 8'h00; 
        10'b0111011000: data <= 8'h00; 
        10'b0111011001: data <= 8'h00; 
        10'b0111011010: data <= 8'h00; 
        10'b0111011011: data <= 8'h00; 
        10'b0111011100: data <= 8'h00; 
        10'b0111011101: data <= 8'h00; 
        10'b0111011110: data <= 8'h00; 
        10'b0111011111: data <= 8'h00; 
        10'b0111100000: data <= 8'h00; 
        10'b0111100001: data <= 8'h00; 
        10'b0111100010: data <= 8'h00; 
        10'b0111100011: data <= 8'h01; 
        10'b0111100100: data <= 8'h01; 
        10'b0111100101: data <= 8'h01; 
        10'b0111100110: data <= 8'h00; 
        10'b0111100111: data <= 8'h00; 
        10'b0111101000: data <= 8'h01; 
        10'b0111101001: data <= 8'h01; 
        10'b0111101010: data <= 8'h02; 
        10'b0111101011: data <= 8'h02; 
        10'b0111101100: data <= 8'h01; 
        10'b0111101101: data <= 8'h00; 
        10'b0111101110: data <= 8'h00; 
        10'b0111101111: data <= 8'h00; 
        10'b0111110000: data <= 8'h00; 
        10'b0111110001: data <= 8'h00; 
        10'b0111110010: data <= 8'h00; 
        10'b0111110011: data <= 8'h00; 
        10'b0111110100: data <= 8'h00; 
        10'b0111110101: data <= 8'h00; 
        10'b0111110110: data <= 8'h00; 
        10'b0111110111: data <= 8'h00; 
        10'b0111111000: data <= 8'h00; 
        10'b0111111001: data <= 8'h00; 
        10'b0111111010: data <= 8'h00; 
        10'b0111111011: data <= 8'h00; 
        10'b0111111100: data <= 8'h00; 
        10'b0111111101: data <= 8'h00; 
        10'b0111111110: data <= 8'h00; 
        10'b0111111111: data <= 8'h00; 
        10'b1000000000: data <= 8'h00; 
        10'b1000000001: data <= 8'h00; 
        10'b1000000010: data <= 8'h00; 
        10'b1000000011: data <= 8'h00; 
        10'b1000000100: data <= 8'h00; 
        10'b1000000101: data <= 8'h01; 
        10'b1000000110: data <= 8'h01; 
        10'b1000000111: data <= 8'h01; 
        10'b1000001000: data <= 8'h00; 
        10'b1000001001: data <= 8'hff; 
        10'b1000001010: data <= 8'hff; 
        10'b1000001011: data <= 8'hff; 
        10'b1000001100: data <= 8'hff; 
        10'b1000001101: data <= 8'hff; 
        10'b1000001110: data <= 8'hff; 
        10'b1000001111: data <= 8'hff; 
        10'b1000010000: data <= 8'h00; 
        10'b1000010001: data <= 8'h00; 
        10'b1000010010: data <= 8'h00; 
        10'b1000010011: data <= 8'h00; 
        10'b1000010100: data <= 8'h00; 
        10'b1000010101: data <= 8'h00; 
        10'b1000010110: data <= 8'h00; 
        10'b1000010111: data <= 8'h00; 
        10'b1000011000: data <= 8'h00; 
        10'b1000011001: data <= 8'h00; 
        10'b1000011010: data <= 8'hff; 
        10'b1000011011: data <= 8'hff; 
        10'b1000011100: data <= 8'hff; 
        10'b1000011101: data <= 8'hff; 
        10'b1000011110: data <= 8'hff; 
        10'b1000011111: data <= 8'hff; 
        10'b1000100000: data <= 8'hff; 
        10'b1000100001: data <= 8'hff; 
        10'b1000100010: data <= 8'h00; 
        10'b1000100011: data <= 8'h00; 
        10'b1000100100: data <= 8'hff; 
        10'b1000100101: data <= 8'h00; 
        10'b1000100110: data <= 8'hff; 
        10'b1000100111: data <= 8'hff; 
        10'b1000101000: data <= 8'hff; 
        10'b1000101001: data <= 8'hff; 
        10'b1000101010: data <= 8'hff; 
        10'b1000101011: data <= 8'hff; 
        10'b1000101100: data <= 8'h00; 
        10'b1000101101: data <= 8'h00; 
        10'b1000101110: data <= 8'h00; 
        10'b1000101111: data <= 8'h00; 
        10'b1000110000: data <= 8'h00; 
        10'b1000110001: data <= 8'h00; 
        10'b1000110010: data <= 8'h00; 
        10'b1000110011: data <= 8'h00; 
        10'b1000110100: data <= 8'h00; 
        10'b1000110101: data <= 8'hff; 
        10'b1000110110: data <= 8'hff; 
        10'b1000110111: data <= 8'hff; 
        10'b1000111000: data <= 8'hfe; 
        10'b1000111001: data <= 8'hfe; 
        10'b1000111010: data <= 8'hfe; 
        10'b1000111011: data <= 8'hff; 
        10'b1000111100: data <= 8'hff; 
        10'b1000111101: data <= 8'hff; 
        10'b1000111110: data <= 8'hff; 
        10'b1000111111: data <= 8'h00; 
        10'b1001000000: data <= 8'h00; 
        10'b1001000001: data <= 8'h00; 
        10'b1001000010: data <= 8'h00; 
        10'b1001000011: data <= 8'hff; 
        10'b1001000100: data <= 8'h00; 
        10'b1001000101: data <= 8'h00; 
        10'b1001000110: data <= 8'hff; 
        10'b1001000111: data <= 8'h00; 
        10'b1001001000: data <= 8'h00; 
        10'b1001001001: data <= 8'h00; 
        10'b1001001010: data <= 8'h00; 
        10'b1001001011: data <= 8'h00; 
        10'b1001001100: data <= 8'h00; 
        10'b1001001101: data <= 8'h00; 
        10'b1001001110: data <= 8'h00; 
        10'b1001001111: data <= 8'h00; 
        10'b1001010000: data <= 8'h00; 
        10'b1001010001: data <= 8'h00; 
        10'b1001010010: data <= 8'hff; 
        10'b1001010011: data <= 8'hff; 
        10'b1001010100: data <= 8'hff; 
        10'b1001010101: data <= 8'hff; 
        10'b1001010110: data <= 8'hff; 
        10'b1001010111: data <= 8'hff; 
        10'b1001011000: data <= 8'hff; 
        10'b1001011001: data <= 8'hff; 
        10'b1001011010: data <= 8'hff; 
        10'b1001011011: data <= 8'h00; 
        10'b1001011100: data <= 8'h00; 
        10'b1001011101: data <= 8'h00; 
        10'b1001011110: data <= 8'h00; 
        10'b1001011111: data <= 8'h00; 
        10'b1001100000: data <= 8'h00; 
        10'b1001100001: data <= 8'h00; 
        10'b1001100010: data <= 8'h00; 
        10'b1001100011: data <= 8'h00; 
        10'b1001100100: data <= 8'h00; 
        10'b1001100101: data <= 8'h00; 
        10'b1001100110: data <= 8'h00; 
        10'b1001100111: data <= 8'h00; 
        10'b1001101000: data <= 8'h00; 
        10'b1001101001: data <= 8'h00; 
        10'b1001101010: data <= 8'h00; 
        10'b1001101011: data <= 8'h00; 
        10'b1001101100: data <= 8'h00; 
        10'b1001101101: data <= 8'h00; 
        10'b1001101110: data <= 8'h00; 
        10'b1001101111: data <= 8'hff; 
        10'b1001110000: data <= 8'hff; 
        10'b1001110001: data <= 8'h00; 
        10'b1001110010: data <= 8'h00; 
        10'b1001110011: data <= 8'h00; 
        10'b1001110100: data <= 8'h00; 
        10'b1001110101: data <= 8'h00; 
        10'b1001110110: data <= 8'h00; 
        10'b1001110111: data <= 8'h00; 
        10'b1001111000: data <= 8'h00; 
        10'b1001111001: data <= 8'h00; 
        10'b1001111010: data <= 8'h00; 
        10'b1001111011: data <= 8'h01; 
        10'b1001111100: data <= 8'h00; 
        10'b1001111101: data <= 8'h00; 
        10'b1001111110: data <= 8'h00; 
        10'b1001111111: data <= 8'h00; 
        10'b1010000000: data <= 8'h00; 
        10'b1010000001: data <= 8'h00; 
        10'b1010000010: data <= 8'h00; 
        10'b1010000011: data <= 8'h00; 
        10'b1010000100: data <= 8'h00; 
        10'b1010000101: data <= 8'h00; 
        10'b1010000110: data <= 8'h00; 
        10'b1010000111: data <= 8'h00; 
        10'b1010001000: data <= 8'h00; 
        10'b1010001001: data <= 8'h00; 
        10'b1010001010: data <= 8'h00; 
        10'b1010001011: data <= 8'h00; 
        10'b1010001100: data <= 8'h00; 
        10'b1010001101: data <= 8'h00; 
        10'b1010001110: data <= 8'h00; 
        10'b1010001111: data <= 8'h00; 
        10'b1010010000: data <= 8'h00; 
        10'b1010010001: data <= 8'h00; 
        10'b1010010010: data <= 8'h00; 
        10'b1010010011: data <= 8'h00; 
        10'b1010010100: data <= 8'h00; 
        10'b1010010101: data <= 8'h00; 
        10'b1010010110: data <= 8'h01; 
        10'b1010010111: data <= 8'h01; 
        10'b1010011000: data <= 8'h00; 
        10'b1010011001: data <= 8'h00; 
        10'b1010011010: data <= 8'h00; 
        10'b1010011011: data <= 8'h00; 
        10'b1010011100: data <= 8'h00; 
        10'b1010011101: data <= 8'h00; 
        10'b1010011110: data <= 8'h00; 
        10'b1010011111: data <= 8'h00; 
        10'b1010100000: data <= 8'h00; 
        10'b1010100001: data <= 8'h00; 
        10'b1010100010: data <= 8'h00; 
        10'b1010100011: data <= 8'h00; 
        10'b1010100100: data <= 8'h00; 
        10'b1010100101: data <= 8'h00; 
        10'b1010100110: data <= 8'h00; 
        10'b1010100111: data <= 8'h00; 
        10'b1010101000: data <= 8'h00; 
        10'b1010101001: data <= 8'h00; 
        10'b1010101010: data <= 8'h00; 
        10'b1010101011: data <= 8'h00; 
        10'b1010101100: data <= 8'h00; 
        10'b1010101101: data <= 8'h00; 
        10'b1010101110: data <= 8'h00; 
        10'b1010101111: data <= 8'h00; 
        10'b1010110000: data <= 8'h00; 
        10'b1010110001: data <= 8'h00; 
        10'b1010110010: data <= 8'h00; 
        10'b1010110011: data <= 8'h00; 
        10'b1010110100: data <= 8'h00; 
        10'b1010110101: data <= 8'h00; 
        10'b1010110110: data <= 8'h00; 
        10'b1010110111: data <= 8'h00; 
        10'b1010111000: data <= 8'h00; 
        10'b1010111001: data <= 8'h00; 
        10'b1010111010: data <= 8'h00; 
        10'b1010111011: data <= 8'h00; 
        10'b1010111100: data <= 8'h00; 
        10'b1010111101: data <= 8'h00; 
        10'b1010111110: data <= 8'h00; 
        10'b1010111111: data <= 8'h00; 
        10'b1011000000: data <= 8'h00; 
        10'b1011000001: data <= 8'h00; 
        10'b1011000010: data <= 8'h00; 
        10'b1011000011: data <= 8'h00; 
        10'b1011000100: data <= 8'h00; 
        10'b1011000101: data <= 8'h00; 
        10'b1011000110: data <= 8'hff; 
        10'b1011000111: data <= 8'hff; 
        10'b1011001000: data <= 8'hff; 
        10'b1011001001: data <= 8'hff; 
        10'b1011001010: data <= 8'hff; 
        10'b1011001011: data <= 8'hff; 
        10'b1011001100: data <= 8'hff; 
        10'b1011001101: data <= 8'hff; 
        10'b1011001110: data <= 8'hff; 
        10'b1011001111: data <= 8'h00; 
        10'b1011010000: data <= 8'h00; 
        10'b1011010001: data <= 8'h00; 
        10'b1011010010: data <= 8'h00; 
        10'b1011010011: data <= 8'h00; 
        10'b1011010100: data <= 8'h00; 
        10'b1011010101: data <= 8'h00; 
        10'b1011010110: data <= 8'h00; 
        10'b1011010111: data <= 8'h00; 
        10'b1011011000: data <= 8'h00; 
        10'b1011011001: data <= 8'h00; 
        10'b1011011010: data <= 8'h00; 
        10'b1011011011: data <= 8'h00; 
        10'b1011011100: data <= 8'h00; 
        10'b1011011101: data <= 8'h00; 
        10'b1011011110: data <= 8'h00; 
        10'b1011011111: data <= 8'h00; 
        10'b1011100000: data <= 8'h00; 
        10'b1011100001: data <= 8'h00; 
        10'b1011100010: data <= 8'hff; 
        10'b1011100011: data <= 8'h00; 
        10'b1011100100: data <= 8'hff; 
        10'b1011100101: data <= 8'hff; 
        10'b1011100110: data <= 8'hff; 
        10'b1011100111: data <= 8'hff; 
        10'b1011101000: data <= 8'hff; 
        10'b1011101001: data <= 8'hff; 
        10'b1011101010: data <= 8'hff; 
        10'b1011101011: data <= 8'h00; 
        10'b1011101100: data <= 8'h00; 
        10'b1011101101: data <= 8'h00; 
        10'b1011101110: data <= 8'h00; 
        10'b1011101111: data <= 8'h00; 
        10'b1011110000: data <= 8'h00; 
        10'b1011110001: data <= 8'h00; 
        10'b1011110010: data <= 8'h00; 
        10'b1011110011: data <= 8'h00; 
        10'b1011110100: data <= 8'h00; 
        10'b1011110101: data <= 8'h00; 
        10'b1011110110: data <= 8'h00; 
        10'b1011110111: data <= 8'h00; 
        10'b1011111000: data <= 8'h00; 
        10'b1011111001: data <= 8'h00; 
        10'b1011111010: data <= 8'h00; 
        10'b1011111011: data <= 8'h00; 
        10'b1011111100: data <= 8'h00; 
        10'b1011111101: data <= 8'h00; 
        10'b1011111110: data <= 8'h00; 
        10'b1011111111: data <= 8'h00; 
        10'b1100000000: data <= 8'h00; 
        10'b1100000001: data <= 8'h00; 
        10'b1100000010: data <= 8'h00; 
        10'b1100000011: data <= 8'h00; 
        10'b1100000100: data <= 8'h00; 
        10'b1100000101: data <= 8'h00; 
        10'b1100000110: data <= 8'h00; 
        10'b1100000111: data <= 8'h00; 
        10'b1100001000: data <= 8'h00; 
        10'b1100001001: data <= 8'h00; 
        10'b1100001010: data <= 8'h00; 
        10'b1100001011: data <= 8'h00; 
        10'b1100001100: data <= 8'h00; 
        10'b1100001101: data <= 8'h00; 
        10'b1100001110: data <= 8'h00; 
        10'b1100001111: data <= 8'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 3) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 9'h000; 
        10'b0000000001: data <= 9'h000; 
        10'b0000000010: data <= 9'h000; 
        10'b0000000011: data <= 9'h000; 
        10'b0000000100: data <= 9'h000; 
        10'b0000000101: data <= 9'h000; 
        10'b0000000110: data <= 9'h000; 
        10'b0000000111: data <= 9'h000; 
        10'b0000001000: data <= 9'h000; 
        10'b0000001001: data <= 9'h000; 
        10'b0000001010: data <= 9'h000; 
        10'b0000001011: data <= 9'h000; 
        10'b0000001100: data <= 9'h000; 
        10'b0000001101: data <= 9'h000; 
        10'b0000001110: data <= 9'h000; 
        10'b0000001111: data <= 9'h000; 
        10'b0000010000: data <= 9'h000; 
        10'b0000010001: data <= 9'h000; 
        10'b0000010010: data <= 9'h000; 
        10'b0000010011: data <= 9'h000; 
        10'b0000010100: data <= 9'h000; 
        10'b0000010101: data <= 9'h000; 
        10'b0000010110: data <= 9'h000; 
        10'b0000010111: data <= 9'h000; 
        10'b0000011000: data <= 9'h000; 
        10'b0000011001: data <= 9'h000; 
        10'b0000011010: data <= 9'h000; 
        10'b0000011011: data <= 9'h000; 
        10'b0000011100: data <= 9'h000; 
        10'b0000011101: data <= 9'h000; 
        10'b0000011110: data <= 9'h000; 
        10'b0000011111: data <= 9'h000; 
        10'b0000100000: data <= 9'h000; 
        10'b0000100001: data <= 9'h001; 
        10'b0000100010: data <= 9'h000; 
        10'b0000100011: data <= 9'h000; 
        10'b0000100100: data <= 9'h000; 
        10'b0000100101: data <= 9'h000; 
        10'b0000100110: data <= 9'h000; 
        10'b0000100111: data <= 9'h000; 
        10'b0000101000: data <= 9'h000; 
        10'b0000101001: data <= 9'h000; 
        10'b0000101010: data <= 9'h000; 
        10'b0000101011: data <= 9'h000; 
        10'b0000101100: data <= 9'h000; 
        10'b0000101101: data <= 9'h000; 
        10'b0000101110: data <= 9'h000; 
        10'b0000101111: data <= 9'h000; 
        10'b0000110000: data <= 9'h000; 
        10'b0000110001: data <= 9'h000; 
        10'b0000110010: data <= 9'h000; 
        10'b0000110011: data <= 9'h000; 
        10'b0000110100: data <= 9'h000; 
        10'b0000110101: data <= 9'h000; 
        10'b0000110110: data <= 9'h000; 
        10'b0000110111: data <= 9'h000; 
        10'b0000111000: data <= 9'h000; 
        10'b0000111001: data <= 9'h000; 
        10'b0000111010: data <= 9'h000; 
        10'b0000111011: data <= 9'h000; 
        10'b0000111100: data <= 9'h000; 
        10'b0000111101: data <= 9'h000; 
        10'b0000111110: data <= 9'h000; 
        10'b0000111111: data <= 9'h000; 
        10'b0001000000: data <= 9'h000; 
        10'b0001000001: data <= 9'h000; 
        10'b0001000010: data <= 9'h000; 
        10'b0001000011: data <= 9'h000; 
        10'b0001000100: data <= 9'h1ff; 
        10'b0001000101: data <= 9'h000; 
        10'b0001000110: data <= 9'h1ff; 
        10'b0001000111: data <= 9'h1ff; 
        10'b0001001000: data <= 9'h1ff; 
        10'b0001001001: data <= 9'h000; 
        10'b0001001010: data <= 9'h000; 
        10'b0001001011: data <= 9'h000; 
        10'b0001001100: data <= 9'h000; 
        10'b0001001101: data <= 9'h000; 
        10'b0001001110: data <= 9'h000; 
        10'b0001001111: data <= 9'h000; 
        10'b0001010000: data <= 9'h000; 
        10'b0001010001: data <= 9'h000; 
        10'b0001010010: data <= 9'h000; 
        10'b0001010011: data <= 9'h000; 
        10'b0001010100: data <= 9'h000; 
        10'b0001010101: data <= 9'h000; 
        10'b0001010110: data <= 9'h000; 
        10'b0001010111: data <= 9'h000; 
        10'b0001011000: data <= 9'h000; 
        10'b0001011001: data <= 9'h000; 
        10'b0001011010: data <= 9'h000; 
        10'b0001011011: data <= 9'h000; 
        10'b0001011100: data <= 9'h000; 
        10'b0001011101: data <= 9'h000; 
        10'b0001011110: data <= 9'h1ff; 
        10'b0001011111: data <= 9'h1ff; 
        10'b0001100000: data <= 9'h1fe; 
        10'b0001100001: data <= 9'h1fe; 
        10'b0001100010: data <= 9'h1fe; 
        10'b0001100011: data <= 9'h1fe; 
        10'b0001100100: data <= 9'h1ff; 
        10'b0001100101: data <= 9'h1ff; 
        10'b0001100110: data <= 9'h000; 
        10'b0001100111: data <= 9'h000; 
        10'b0001101000: data <= 9'h000; 
        10'b0001101001: data <= 9'h001; 
        10'b0001101010: data <= 9'h000; 
        10'b0001101011: data <= 9'h000; 
        10'b0001101100: data <= 9'h001; 
        10'b0001101101: data <= 9'h001; 
        10'b0001101110: data <= 9'h000; 
        10'b0001101111: data <= 9'h000; 
        10'b0001110000: data <= 9'h001; 
        10'b0001110001: data <= 9'h000; 
        10'b0001110010: data <= 9'h000; 
        10'b0001110011: data <= 9'h000; 
        10'b0001110100: data <= 9'h000; 
        10'b0001110101: data <= 9'h000; 
        10'b0001110110: data <= 9'h000; 
        10'b0001110111: data <= 9'h000; 
        10'b0001111000: data <= 9'h1ff; 
        10'b0001111001: data <= 9'h1ff; 
        10'b0001111010: data <= 9'h1fe; 
        10'b0001111011: data <= 9'h1ff; 
        10'b0001111100: data <= 9'h1fe; 
        10'b0001111101: data <= 9'h1fe; 
        10'b0001111110: data <= 9'h1fe; 
        10'b0001111111: data <= 9'h1fe; 
        10'b0010000000: data <= 9'h1ff; 
        10'b0010000001: data <= 9'h1ff; 
        10'b0010000010: data <= 9'h000; 
        10'b0010000011: data <= 9'h000; 
        10'b0010000100: data <= 9'h001; 
        10'b0010000101: data <= 9'h001; 
        10'b0010000110: data <= 9'h001; 
        10'b0010000111: data <= 9'h001; 
        10'b0010001000: data <= 9'h000; 
        10'b0010001001: data <= 9'h000; 
        10'b0010001010: data <= 9'h000; 
        10'b0010001011: data <= 9'h000; 
        10'b0010001100: data <= 9'h001; 
        10'b0010001101: data <= 9'h000; 
        10'b0010001110: data <= 9'h000; 
        10'b0010001111: data <= 9'h000; 
        10'b0010010000: data <= 9'h000; 
        10'b0010010001: data <= 9'h000; 
        10'b0010010010: data <= 9'h000; 
        10'b0010010011: data <= 9'h000; 
        10'b0010010100: data <= 9'h000; 
        10'b0010010101: data <= 9'h000; 
        10'b0010010110: data <= 9'h1ff; 
        10'b0010010111: data <= 9'h1ff; 
        10'b0010011000: data <= 9'h1ff; 
        10'b0010011001: data <= 9'h1fe; 
        10'b0010011010: data <= 9'h1ff; 
        10'b0010011011: data <= 9'h1ff; 
        10'b0010011100: data <= 9'h000; 
        10'b0010011101: data <= 9'h000; 
        10'b0010011110: data <= 9'h000; 
        10'b0010011111: data <= 9'h000; 
        10'b0010100000: data <= 9'h000; 
        10'b0010100001: data <= 9'h001; 
        10'b0010100010: data <= 9'h001; 
        10'b0010100011: data <= 9'h002; 
        10'b0010100100: data <= 9'h001; 
        10'b0010100101: data <= 9'h000; 
        10'b0010100110: data <= 9'h000; 
        10'b0010100111: data <= 9'h000; 
        10'b0010101000: data <= 9'h000; 
        10'b0010101001: data <= 9'h001; 
        10'b0010101010: data <= 9'h000; 
        10'b0010101011: data <= 9'h000; 
        10'b0010101100: data <= 9'h000; 
        10'b0010101101: data <= 9'h000; 
        10'b0010101110: data <= 9'h000; 
        10'b0010101111: data <= 9'h000; 
        10'b0010110000: data <= 9'h000; 
        10'b0010110001: data <= 9'h000; 
        10'b0010110010: data <= 9'h1ff; 
        10'b0010110011: data <= 9'h1fe; 
        10'b0010110100: data <= 9'h1fe; 
        10'b0010110101: data <= 9'h1fd; 
        10'b0010110110: data <= 9'h1fd; 
        10'b0010110111: data <= 9'h1fd; 
        10'b0010111000: data <= 9'h1fd; 
        10'b0010111001: data <= 9'h1fe; 
        10'b0010111010: data <= 9'h1fe; 
        10'b0010111011: data <= 9'h1ff; 
        10'b0010111100: data <= 9'h000; 
        10'b0010111101: data <= 9'h000; 
        10'b0010111110: data <= 9'h002; 
        10'b0010111111: data <= 9'h002; 
        10'b0011000000: data <= 9'h001; 
        10'b0011000001: data <= 9'h001; 
        10'b0011000010: data <= 9'h000; 
        10'b0011000011: data <= 9'h000; 
        10'b0011000100: data <= 9'h000; 
        10'b0011000101: data <= 9'h000; 
        10'b0011000110: data <= 9'h000; 
        10'b0011000111: data <= 9'h000; 
        10'b0011001000: data <= 9'h000; 
        10'b0011001001: data <= 9'h000; 
        10'b0011001010: data <= 9'h000; 
        10'b0011001011: data <= 9'h000; 
        10'b0011001100: data <= 9'h000; 
        10'b0011001101: data <= 9'h1ff; 
        10'b0011001110: data <= 9'h1fe; 
        10'b0011001111: data <= 9'h1fe; 
        10'b0011010000: data <= 9'h1fd; 
        10'b0011010001: data <= 9'h1fe; 
        10'b0011010010: data <= 9'h1fd; 
        10'b0011010011: data <= 9'h1fd; 
        10'b0011010100: data <= 9'h1fd; 
        10'b0011010101: data <= 9'h1fe; 
        10'b0011010110: data <= 9'h1fe; 
        10'b0011010111: data <= 9'h1ff; 
        10'b0011011000: data <= 9'h1fe; 
        10'b0011011001: data <= 9'h1ff; 
        10'b0011011010: data <= 9'h001; 
        10'b0011011011: data <= 9'h002; 
        10'b0011011100: data <= 9'h001; 
        10'b0011011101: data <= 9'h001; 
        10'b0011011110: data <= 9'h000; 
        10'b0011011111: data <= 9'h000; 
        10'b0011100000: data <= 9'h000; 
        10'b0011100001: data <= 9'h000; 
        10'b0011100010: data <= 9'h001; 
        10'b0011100011: data <= 9'h000; 
        10'b0011100100: data <= 9'h000; 
        10'b0011100101: data <= 9'h000; 
        10'b0011100110: data <= 9'h000; 
        10'b0011100111: data <= 9'h000; 
        10'b0011101000: data <= 9'h1ff; 
        10'b0011101001: data <= 9'h1ff; 
        10'b0011101010: data <= 9'h1ff; 
        10'b0011101011: data <= 9'h1fe; 
        10'b0011101100: data <= 9'h1fe; 
        10'b0011101101: data <= 9'h1ff; 
        10'b0011101110: data <= 9'h1fd; 
        10'b0011101111: data <= 9'h1fd; 
        10'b0011110000: data <= 9'h1fd; 
        10'b0011110001: data <= 9'h1fe; 
        10'b0011110010: data <= 9'h1ff; 
        10'b0011110011: data <= 9'h000; 
        10'b0011110100: data <= 9'h1ff; 
        10'b0011110101: data <= 9'h1ff; 
        10'b0011110110: data <= 9'h001; 
        10'b0011110111: data <= 9'h001; 
        10'b0011111000: data <= 9'h001; 
        10'b0011111001: data <= 9'h000; 
        10'b0011111010: data <= 9'h000; 
        10'b0011111011: data <= 9'h000; 
        10'b0011111100: data <= 9'h001; 
        10'b0011111101: data <= 9'h000; 
        10'b0011111110: data <= 9'h000; 
        10'b0011111111: data <= 9'h000; 
        10'b0100000000: data <= 9'h000; 
        10'b0100000001: data <= 9'h000; 
        10'b0100000010: data <= 9'h1ff; 
        10'b0100000011: data <= 9'h1ff; 
        10'b0100000100: data <= 9'h000; 
        10'b0100000101: data <= 9'h000; 
        10'b0100000110: data <= 9'h000; 
        10'b0100000111: data <= 9'h000; 
        10'b0100001000: data <= 9'h000; 
        10'b0100001001: data <= 9'h1ff; 
        10'b0100001010: data <= 9'h1fb; 
        10'b0100001011: data <= 9'h1fc; 
        10'b0100001100: data <= 9'h1ff; 
        10'b0100001101: data <= 9'h1ff; 
        10'b0100001110: data <= 9'h000; 
        10'b0100001111: data <= 9'h000; 
        10'b0100010000: data <= 9'h000; 
        10'b0100010001: data <= 9'h000; 
        10'b0100010010: data <= 9'h000; 
        10'b0100010011: data <= 9'h000; 
        10'b0100010100: data <= 9'h1ff; 
        10'b0100010101: data <= 9'h1ff; 
        10'b0100010110: data <= 9'h000; 
        10'b0100010111: data <= 9'h000; 
        10'b0100011000: data <= 9'h000; 
        10'b0100011001: data <= 9'h000; 
        10'b0100011010: data <= 9'h000; 
        10'b0100011011: data <= 9'h000; 
        10'b0100011100: data <= 9'h000; 
        10'b0100011101: data <= 9'h1ff; 
        10'b0100011110: data <= 9'h1ff; 
        10'b0100011111: data <= 9'h1ff; 
        10'b0100100000: data <= 9'h000; 
        10'b0100100001: data <= 9'h001; 
        10'b0100100010: data <= 9'h001; 
        10'b0100100011: data <= 9'h001; 
        10'b0100100100: data <= 9'h001; 
        10'b0100100101: data <= 9'h1fe; 
        10'b0100100110: data <= 9'h1fb; 
        10'b0100100111: data <= 9'h1fe; 
        10'b0100101000: data <= 9'h000; 
        10'b0100101001: data <= 9'h000; 
        10'b0100101010: data <= 9'h000; 
        10'b0100101011: data <= 9'h000; 
        10'b0100101100: data <= 9'h1ff; 
        10'b0100101101: data <= 9'h1ff; 
        10'b0100101110: data <= 9'h000; 
        10'b0100101111: data <= 9'h1ff; 
        10'b0100110000: data <= 9'h1ff; 
        10'b0100110001: data <= 9'h000; 
        10'b0100110010: data <= 9'h000; 
        10'b0100110011: data <= 9'h001; 
        10'b0100110100: data <= 9'h000; 
        10'b0100110101: data <= 9'h000; 
        10'b0100110110: data <= 9'h000; 
        10'b0100110111: data <= 9'h000; 
        10'b0100111000: data <= 9'h000; 
        10'b0100111001: data <= 9'h000; 
        10'b0100111010: data <= 9'h000; 
        10'b0100111011: data <= 9'h000; 
        10'b0100111100: data <= 9'h001; 
        10'b0100111101: data <= 9'h002; 
        10'b0100111110: data <= 9'h002; 
        10'b0100111111: data <= 9'h002; 
        10'b0101000000: data <= 9'h002; 
        10'b0101000001: data <= 9'h1fd; 
        10'b0101000010: data <= 9'h1fc; 
        10'b0101000011: data <= 9'h000; 
        10'b0101000100: data <= 9'h002; 
        10'b0101000101: data <= 9'h000; 
        10'b0101000110: data <= 9'h000; 
        10'b0101000111: data <= 9'h000; 
        10'b0101001000: data <= 9'h1ff; 
        10'b0101001001: data <= 9'h1ff; 
        10'b0101001010: data <= 9'h000; 
        10'b0101001011: data <= 9'h1ff; 
        10'b0101001100: data <= 9'h1ff; 
        10'b0101001101: data <= 9'h000; 
        10'b0101001110: data <= 9'h000; 
        10'b0101001111: data <= 9'h000; 
        10'b0101010000: data <= 9'h000; 
        10'b0101010001: data <= 9'h000; 
        10'b0101010010: data <= 9'h000; 
        10'b0101010011: data <= 9'h000; 
        10'b0101010100: data <= 9'h000; 
        10'b0101010101: data <= 9'h000; 
        10'b0101010110: data <= 9'h001; 
        10'b0101010111: data <= 9'h002; 
        10'b0101011000: data <= 9'h003; 
        10'b0101011001: data <= 9'h002; 
        10'b0101011010: data <= 9'h004; 
        10'b0101011011: data <= 9'h004; 
        10'b0101011100: data <= 9'h004; 
        10'b0101011101: data <= 9'h000; 
        10'b0101011110: data <= 9'h1fe; 
        10'b0101011111: data <= 9'h002; 
        10'b0101100000: data <= 9'h003; 
        10'b0101100001: data <= 9'h000; 
        10'b0101100010: data <= 9'h000; 
        10'b0101100011: data <= 9'h000; 
        10'b0101100100: data <= 9'h000; 
        10'b0101100101: data <= 9'h000; 
        10'b0101100110: data <= 9'h000; 
        10'b0101100111: data <= 9'h1ff; 
        10'b0101101000: data <= 9'h1ff; 
        10'b0101101001: data <= 9'h000; 
        10'b0101101010: data <= 9'h001; 
        10'b0101101011: data <= 9'h000; 
        10'b0101101100: data <= 9'h000; 
        10'b0101101101: data <= 9'h000; 
        10'b0101101110: data <= 9'h000; 
        10'b0101101111: data <= 9'h000; 
        10'b0101110000: data <= 9'h000; 
        10'b0101110001: data <= 9'h001; 
        10'b0101110010: data <= 9'h002; 
        10'b0101110011: data <= 9'h003; 
        10'b0101110100: data <= 9'h003; 
        10'b0101110101: data <= 9'h003; 
        10'b0101110110: data <= 9'h003; 
        10'b0101110111: data <= 9'h005; 
        10'b0101111000: data <= 9'h004; 
        10'b0101111001: data <= 9'h000; 
        10'b0101111010: data <= 9'h1ff; 
        10'b0101111011: data <= 9'h002; 
        10'b0101111100: data <= 9'h002; 
        10'b0101111101: data <= 9'h002; 
        10'b0101111110: data <= 9'h001; 
        10'b0101111111: data <= 9'h001; 
        10'b0110000000: data <= 9'h001; 
        10'b0110000001: data <= 9'h001; 
        10'b0110000010: data <= 9'h001; 
        10'b0110000011: data <= 9'h000; 
        10'b0110000100: data <= 9'h000; 
        10'b0110000101: data <= 9'h000; 
        10'b0110000110: data <= 9'h000; 
        10'b0110000111: data <= 9'h000; 
        10'b0110001000: data <= 9'h000; 
        10'b0110001001: data <= 9'h000; 
        10'b0110001010: data <= 9'h000; 
        10'b0110001011: data <= 9'h001; 
        10'b0110001100: data <= 9'h001; 
        10'b0110001101: data <= 9'h002; 
        10'b0110001110: data <= 9'h003; 
        10'b0110001111: data <= 9'h003; 
        10'b0110010000: data <= 9'h002; 
        10'b0110010001: data <= 9'h002; 
        10'b0110010010: data <= 9'h003; 
        10'b0110010011: data <= 9'h003; 
        10'b0110010100: data <= 9'h002; 
        10'b0110010101: data <= 9'h000; 
        10'b0110010110: data <= 9'h000; 
        10'b0110010111: data <= 9'h001; 
        10'b0110011000: data <= 9'h002; 
        10'b0110011001: data <= 9'h003; 
        10'b0110011010: data <= 9'h002; 
        10'b0110011011: data <= 9'h002; 
        10'b0110011100: data <= 9'h001; 
        10'b0110011101: data <= 9'h001; 
        10'b0110011110: data <= 9'h000; 
        10'b0110011111: data <= 9'h000; 
        10'b0110100000: data <= 9'h000; 
        10'b0110100001: data <= 9'h000; 
        10'b0110100010: data <= 9'h000; 
        10'b0110100011: data <= 9'h000; 
        10'b0110100100: data <= 9'h000; 
        10'b0110100101: data <= 9'h001; 
        10'b0110100110: data <= 9'h000; 
        10'b0110100111: data <= 9'h000; 
        10'b0110101000: data <= 9'h001; 
        10'b0110101001: data <= 9'h001; 
        10'b0110101010: data <= 9'h002; 
        10'b0110101011: data <= 9'h002; 
        10'b0110101100: data <= 9'h003; 
        10'b0110101101: data <= 9'h002; 
        10'b0110101110: data <= 9'h002; 
        10'b0110101111: data <= 9'h001; 
        10'b0110110000: data <= 9'h001; 
        10'b0110110001: data <= 9'h000; 
        10'b0110110010: data <= 9'h001; 
        10'b0110110011: data <= 9'h001; 
        10'b0110110100: data <= 9'h003; 
        10'b0110110101: data <= 9'h003; 
        10'b0110110110: data <= 9'h002; 
        10'b0110110111: data <= 9'h001; 
        10'b0110111000: data <= 9'h000; 
        10'b0110111001: data <= 9'h000; 
        10'b0110111010: data <= 9'h001; 
        10'b0110111011: data <= 9'h000; 
        10'b0110111100: data <= 9'h000; 
        10'b0110111101: data <= 9'h000; 
        10'b0110111110: data <= 9'h000; 
        10'b0110111111: data <= 9'h000; 
        10'b0111000000: data <= 9'h000; 
        10'b0111000001: data <= 9'h000; 
        10'b0111000010: data <= 9'h000; 
        10'b0111000011: data <= 9'h000; 
        10'b0111000100: data <= 9'h000; 
        10'b0111000101: data <= 9'h001; 
        10'b0111000110: data <= 9'h001; 
        10'b0111000111: data <= 9'h002; 
        10'b0111001000: data <= 9'h003; 
        10'b0111001001: data <= 9'h002; 
        10'b0111001010: data <= 9'h001; 
        10'b0111001011: data <= 9'h000; 
        10'b0111001100: data <= 9'h001; 
        10'b0111001101: data <= 9'h001; 
        10'b0111001110: data <= 9'h002; 
        10'b0111001111: data <= 9'h003; 
        10'b0111010000: data <= 9'h004; 
        10'b0111010001: data <= 9'h003; 
        10'b0111010010: data <= 9'h002; 
        10'b0111010011: data <= 9'h000; 
        10'b0111010100: data <= 9'h001; 
        10'b0111010101: data <= 9'h001; 
        10'b0111010110: data <= 9'h000; 
        10'b0111010111: data <= 9'h000; 
        10'b0111011000: data <= 9'h000; 
        10'b0111011001: data <= 9'h000; 
        10'b0111011010: data <= 9'h000; 
        10'b0111011011: data <= 9'h000; 
        10'b0111011100: data <= 9'h000; 
        10'b0111011101: data <= 9'h000; 
        10'b0111011110: data <= 9'h000; 
        10'b0111011111: data <= 9'h000; 
        10'b0111100000: data <= 9'h000; 
        10'b0111100001: data <= 9'h1ff; 
        10'b0111100010: data <= 9'h000; 
        10'b0111100011: data <= 9'h001; 
        10'b0111100100: data <= 9'h003; 
        10'b0111100101: data <= 9'h002; 
        10'b0111100110: data <= 9'h001; 
        10'b0111100111: data <= 9'h001; 
        10'b0111101000: data <= 9'h001; 
        10'b0111101001: data <= 9'h002; 
        10'b0111101010: data <= 9'h004; 
        10'b0111101011: data <= 9'h003; 
        10'b0111101100: data <= 9'h003; 
        10'b0111101101: data <= 9'h001; 
        10'b0111101110: data <= 9'h000; 
        10'b0111101111: data <= 9'h1ff; 
        10'b0111110000: data <= 9'h000; 
        10'b0111110001: data <= 9'h000; 
        10'b0111110010: data <= 9'h1ff; 
        10'b0111110011: data <= 9'h000; 
        10'b0111110100: data <= 9'h000; 
        10'b0111110101: data <= 9'h000; 
        10'b0111110110: data <= 9'h000; 
        10'b0111110111: data <= 9'h000; 
        10'b0111111000: data <= 9'h000; 
        10'b0111111001: data <= 9'h000; 
        10'b0111111010: data <= 9'h000; 
        10'b0111111011: data <= 9'h000; 
        10'b0111111100: data <= 9'h000; 
        10'b0111111101: data <= 9'h1ff; 
        10'b0111111110: data <= 9'h1ff; 
        10'b0111111111: data <= 9'h000; 
        10'b1000000000: data <= 9'h001; 
        10'b1000000001: data <= 9'h000; 
        10'b1000000010: data <= 9'h1ff; 
        10'b1000000011: data <= 9'h000; 
        10'b1000000100: data <= 9'h001; 
        10'b1000000101: data <= 9'h001; 
        10'b1000000110: data <= 9'h002; 
        10'b1000000111: data <= 9'h002; 
        10'b1000001000: data <= 9'h001; 
        10'b1000001001: data <= 9'h1ff; 
        10'b1000001010: data <= 9'h1ff; 
        10'b1000001011: data <= 9'h1fe; 
        10'b1000001100: data <= 9'h1ff; 
        10'b1000001101: data <= 9'h1ff; 
        10'b1000001110: data <= 9'h1ff; 
        10'b1000001111: data <= 9'h1ff; 
        10'b1000010000: data <= 9'h000; 
        10'b1000010001: data <= 9'h000; 
        10'b1000010010: data <= 9'h000; 
        10'b1000010011: data <= 9'h000; 
        10'b1000010100: data <= 9'h000; 
        10'b1000010101: data <= 9'h000; 
        10'b1000010110: data <= 9'h000; 
        10'b1000010111: data <= 9'h000; 
        10'b1000011000: data <= 9'h1ff; 
        10'b1000011001: data <= 9'h1ff; 
        10'b1000011010: data <= 9'h1ff; 
        10'b1000011011: data <= 9'h1fe; 
        10'b1000011100: data <= 9'h1fe; 
        10'b1000011101: data <= 9'h1fe; 
        10'b1000011110: data <= 9'h1fd; 
        10'b1000011111: data <= 9'h1fd; 
        10'b1000100000: data <= 9'h1fe; 
        10'b1000100001: data <= 9'h1ff; 
        10'b1000100010: data <= 9'h000; 
        10'b1000100011: data <= 9'h000; 
        10'b1000100100: data <= 9'h1ff; 
        10'b1000100101: data <= 9'h1ff; 
        10'b1000100110: data <= 9'h1ff; 
        10'b1000100111: data <= 9'h1fe; 
        10'b1000101000: data <= 9'h1fe; 
        10'b1000101001: data <= 9'h1fe; 
        10'b1000101010: data <= 9'h1fe; 
        10'b1000101011: data <= 9'h1ff; 
        10'b1000101100: data <= 9'h000; 
        10'b1000101101: data <= 9'h000; 
        10'b1000101110: data <= 9'h000; 
        10'b1000101111: data <= 9'h000; 
        10'b1000110000: data <= 9'h001; 
        10'b1000110001: data <= 9'h001; 
        10'b1000110010: data <= 9'h000; 
        10'b1000110011: data <= 9'h000; 
        10'b1000110100: data <= 9'h1ff; 
        10'b1000110101: data <= 9'h1ff; 
        10'b1000110110: data <= 9'h1fe; 
        10'b1000110111: data <= 9'h1fd; 
        10'b1000111000: data <= 9'h1fd; 
        10'b1000111001: data <= 9'h1fd; 
        10'b1000111010: data <= 9'h1fd; 
        10'b1000111011: data <= 9'h1fe; 
        10'b1000111100: data <= 9'h1fe; 
        10'b1000111101: data <= 9'h1fe; 
        10'b1000111110: data <= 9'h1ff; 
        10'b1000111111: data <= 9'h1ff; 
        10'b1001000000: data <= 9'h000; 
        10'b1001000001: data <= 9'h000; 
        10'b1001000010: data <= 9'h1ff; 
        10'b1001000011: data <= 9'h1ff; 
        10'b1001000100: data <= 9'h1ff; 
        10'b1001000101: data <= 9'h1ff; 
        10'b1001000110: data <= 9'h1ff; 
        10'b1001000111: data <= 9'h1ff; 
        10'b1001001000: data <= 9'h1ff; 
        10'b1001001001: data <= 9'h000; 
        10'b1001001010: data <= 9'h000; 
        10'b1001001011: data <= 9'h000; 
        10'b1001001100: data <= 9'h000; 
        10'b1001001101: data <= 9'h000; 
        10'b1001001110: data <= 9'h000; 
        10'b1001001111: data <= 9'h000; 
        10'b1001010000: data <= 9'h000; 
        10'b1001010001: data <= 9'h1ff; 
        10'b1001010010: data <= 9'h1fe; 
        10'b1001010011: data <= 9'h1fe; 
        10'b1001010100: data <= 9'h1fe; 
        10'b1001010101: data <= 9'h1fe; 
        10'b1001010110: data <= 9'h1fe; 
        10'b1001010111: data <= 9'h1ff; 
        10'b1001011000: data <= 9'h1ff; 
        10'b1001011001: data <= 9'h1ff; 
        10'b1001011010: data <= 9'h1ff; 
        10'b1001011011: data <= 9'h1ff; 
        10'b1001011100: data <= 9'h1ff; 
        10'b1001011101: data <= 9'h000; 
        10'b1001011110: data <= 9'h000; 
        10'b1001011111: data <= 9'h000; 
        10'b1001100000: data <= 9'h000; 
        10'b1001100001: data <= 9'h1ff; 
        10'b1001100010: data <= 9'h1ff; 
        10'b1001100011: data <= 9'h000; 
        10'b1001100100: data <= 9'h000; 
        10'b1001100101: data <= 9'h000; 
        10'b1001100110: data <= 9'h000; 
        10'b1001100111: data <= 9'h000; 
        10'b1001101000: data <= 9'h000; 
        10'b1001101001: data <= 9'h000; 
        10'b1001101010: data <= 9'h000; 
        10'b1001101011: data <= 9'h000; 
        10'b1001101100: data <= 9'h000; 
        10'b1001101101: data <= 9'h000; 
        10'b1001101110: data <= 9'h1ff; 
        10'b1001101111: data <= 9'h1ff; 
        10'b1001110000: data <= 9'h1ff; 
        10'b1001110001: data <= 9'h1ff; 
        10'b1001110010: data <= 9'h1ff; 
        10'b1001110011: data <= 9'h1ff; 
        10'b1001110100: data <= 9'h1ff; 
        10'b1001110101: data <= 9'h1ff; 
        10'b1001110110: data <= 9'h1ff; 
        10'b1001110111: data <= 9'h000; 
        10'b1001111000: data <= 9'h000; 
        10'b1001111001: data <= 9'h000; 
        10'b1001111010: data <= 9'h001; 
        10'b1001111011: data <= 9'h001; 
        10'b1001111100: data <= 9'h001; 
        10'b1001111101: data <= 9'h001; 
        10'b1001111110: data <= 9'h000; 
        10'b1001111111: data <= 9'h000; 
        10'b1010000000: data <= 9'h000; 
        10'b1010000001: data <= 9'h000; 
        10'b1010000010: data <= 9'h000; 
        10'b1010000011: data <= 9'h000; 
        10'b1010000100: data <= 9'h000; 
        10'b1010000101: data <= 9'h000; 
        10'b1010000110: data <= 9'h000; 
        10'b1010000111: data <= 9'h000; 
        10'b1010001000: data <= 9'h000; 
        10'b1010001001: data <= 9'h000; 
        10'b1010001010: data <= 9'h000; 
        10'b1010001011: data <= 9'h000; 
        10'b1010001100: data <= 9'h1ff; 
        10'b1010001101: data <= 9'h000; 
        10'b1010001110: data <= 9'h1ff; 
        10'b1010001111: data <= 9'h000; 
        10'b1010010000: data <= 9'h1ff; 
        10'b1010010001: data <= 9'h000; 
        10'b1010010010: data <= 9'h000; 
        10'b1010010011: data <= 9'h000; 
        10'b1010010100: data <= 9'h000; 
        10'b1010010101: data <= 9'h000; 
        10'b1010010110: data <= 9'h001; 
        10'b1010010111: data <= 9'h001; 
        10'b1010011000: data <= 9'h001; 
        10'b1010011001: data <= 9'h000; 
        10'b1010011010: data <= 9'h000; 
        10'b1010011011: data <= 9'h000; 
        10'b1010011100: data <= 9'h000; 
        10'b1010011101: data <= 9'h000; 
        10'b1010011110: data <= 9'h000; 
        10'b1010011111: data <= 9'h000; 
        10'b1010100000: data <= 9'h000; 
        10'b1010100001: data <= 9'h000; 
        10'b1010100010: data <= 9'h000; 
        10'b1010100011: data <= 9'h000; 
        10'b1010100100: data <= 9'h000; 
        10'b1010100101: data <= 9'h000; 
        10'b1010100110: data <= 9'h000; 
        10'b1010100111: data <= 9'h1ff; 
        10'b1010101000: data <= 9'h1ff; 
        10'b1010101001: data <= 9'h000; 
        10'b1010101010: data <= 9'h1ff; 
        10'b1010101011: data <= 9'h000; 
        10'b1010101100: data <= 9'h000; 
        10'b1010101101: data <= 9'h000; 
        10'b1010101110: data <= 9'h1ff; 
        10'b1010101111: data <= 9'h1ff; 
        10'b1010110000: data <= 9'h000; 
        10'b1010110001: data <= 9'h000; 
        10'b1010110010: data <= 9'h000; 
        10'b1010110011: data <= 9'h001; 
        10'b1010110100: data <= 9'h000; 
        10'b1010110101: data <= 9'h000; 
        10'b1010110110: data <= 9'h000; 
        10'b1010110111: data <= 9'h000; 
        10'b1010111000: data <= 9'h000; 
        10'b1010111001: data <= 9'h000; 
        10'b1010111010: data <= 9'h000; 
        10'b1010111011: data <= 9'h000; 
        10'b1010111100: data <= 9'h001; 
        10'b1010111101: data <= 9'h000; 
        10'b1010111110: data <= 9'h000; 
        10'b1010111111: data <= 9'h000; 
        10'b1011000000: data <= 9'h000; 
        10'b1011000001: data <= 9'h000; 
        10'b1011000010: data <= 9'h000; 
        10'b1011000011: data <= 9'h1ff; 
        10'b1011000100: data <= 9'h1ff; 
        10'b1011000101: data <= 9'h1ff; 
        10'b1011000110: data <= 9'h1ff; 
        10'b1011000111: data <= 9'h1fe; 
        10'b1011001000: data <= 9'h1ff; 
        10'b1011001001: data <= 9'h1ff; 
        10'b1011001010: data <= 9'h1ff; 
        10'b1011001011: data <= 9'h1ff; 
        10'b1011001100: data <= 9'h1fe; 
        10'b1011001101: data <= 9'h1fe; 
        10'b1011001110: data <= 9'h1fe; 
        10'b1011001111: data <= 9'h1ff; 
        10'b1011010000: data <= 9'h1ff; 
        10'b1011010001: data <= 9'h000; 
        10'b1011010010: data <= 9'h000; 
        10'b1011010011: data <= 9'h000; 
        10'b1011010100: data <= 9'h000; 
        10'b1011010101: data <= 9'h000; 
        10'b1011010110: data <= 9'h000; 
        10'b1011010111: data <= 9'h000; 
        10'b1011011000: data <= 9'h000; 
        10'b1011011001: data <= 9'h000; 
        10'b1011011010: data <= 9'h000; 
        10'b1011011011: data <= 9'h000; 
        10'b1011011100: data <= 9'h000; 
        10'b1011011101: data <= 9'h000; 
        10'b1011011110: data <= 9'h000; 
        10'b1011011111: data <= 9'h000; 
        10'b1011100000: data <= 9'h000; 
        10'b1011100001: data <= 9'h000; 
        10'b1011100010: data <= 9'h1ff; 
        10'b1011100011: data <= 9'h1ff; 
        10'b1011100100: data <= 9'h1ff; 
        10'b1011100101: data <= 9'h1fe; 
        10'b1011100110: data <= 9'h1fe; 
        10'b1011100111: data <= 9'h1ff; 
        10'b1011101000: data <= 9'h1ff; 
        10'b1011101001: data <= 9'h1ff; 
        10'b1011101010: data <= 9'h1ff; 
        10'b1011101011: data <= 9'h1ff; 
        10'b1011101100: data <= 9'h000; 
        10'b1011101101: data <= 9'h000; 
        10'b1011101110: data <= 9'h000; 
        10'b1011101111: data <= 9'h000; 
        10'b1011110000: data <= 9'h000; 
        10'b1011110001: data <= 9'h000; 
        10'b1011110010: data <= 9'h001; 
        10'b1011110011: data <= 9'h000; 
        10'b1011110100: data <= 9'h000; 
        10'b1011110101: data <= 9'h000; 
        10'b1011110110: data <= 9'h000; 
        10'b1011110111: data <= 9'h001; 
        10'b1011111000: data <= 9'h000; 
        10'b1011111001: data <= 9'h000; 
        10'b1011111010: data <= 9'h000; 
        10'b1011111011: data <= 9'h001; 
        10'b1011111100: data <= 9'h000; 
        10'b1011111101: data <= 9'h000; 
        10'b1011111110: data <= 9'h000; 
        10'b1011111111: data <= 9'h000; 
        10'b1100000000: data <= 9'h000; 
        10'b1100000001: data <= 9'h000; 
        10'b1100000010: data <= 9'h000; 
        10'b1100000011: data <= 9'h000; 
        10'b1100000100: data <= 9'h000; 
        10'b1100000101: data <= 9'h000; 
        10'b1100000110: data <= 9'h000; 
        10'b1100000111: data <= 9'h000; 
        10'b1100001000: data <= 9'h000; 
        10'b1100001001: data <= 9'h000; 
        10'b1100001010: data <= 9'h000; 
        10'b1100001011: data <= 9'h000; 
        10'b1100001100: data <= 9'h000; 
        10'b1100001101: data <= 9'h000; 
        10'b1100001110: data <= 9'h000; 
        10'b1100001111: data <= 9'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 4) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 10'h000; 
        10'b0000000001: data <= 10'h000; 
        10'b0000000010: data <= 10'h001; 
        10'b0000000011: data <= 10'h001; 
        10'b0000000100: data <= 10'h000; 
        10'b0000000101: data <= 10'h000; 
        10'b0000000110: data <= 10'h001; 
        10'b0000000111: data <= 10'h000; 
        10'b0000001000: data <= 10'h000; 
        10'b0000001001: data <= 10'h000; 
        10'b0000001010: data <= 10'h000; 
        10'b0000001011: data <= 10'h001; 
        10'b0000001100: data <= 10'h001; 
        10'b0000001101: data <= 10'h001; 
        10'b0000001110: data <= 10'h001; 
        10'b0000001111: data <= 10'h000; 
        10'b0000010000: data <= 10'h001; 
        10'b0000010001: data <= 10'h001; 
        10'b0000010010: data <= 10'h000; 
        10'b0000010011: data <= 10'h001; 
        10'b0000010100: data <= 10'h000; 
        10'b0000010101: data <= 10'h000; 
        10'b0000010110: data <= 10'h001; 
        10'b0000010111: data <= 10'h000; 
        10'b0000011000: data <= 10'h001; 
        10'b0000011001: data <= 10'h000; 
        10'b0000011010: data <= 10'h001; 
        10'b0000011011: data <= 10'h000; 
        10'b0000011100: data <= 10'h000; 
        10'b0000011101: data <= 10'h000; 
        10'b0000011110: data <= 10'h000; 
        10'b0000011111: data <= 10'h000; 
        10'b0000100000: data <= 10'h000; 
        10'b0000100001: data <= 10'h001; 
        10'b0000100010: data <= 10'h000; 
        10'b0000100011: data <= 10'h000; 
        10'b0000100100: data <= 10'h001; 
        10'b0000100101: data <= 10'h000; 
        10'b0000100110: data <= 10'h000; 
        10'b0000100111: data <= 10'h000; 
        10'b0000101000: data <= 10'h000; 
        10'b0000101001: data <= 10'h000; 
        10'b0000101010: data <= 10'h000; 
        10'b0000101011: data <= 10'h001; 
        10'b0000101100: data <= 10'h001; 
        10'b0000101101: data <= 10'h000; 
        10'b0000101110: data <= 10'h000; 
        10'b0000101111: data <= 10'h000; 
        10'b0000110000: data <= 10'h001; 
        10'b0000110001: data <= 10'h000; 
        10'b0000110010: data <= 10'h000; 
        10'b0000110011: data <= 10'h000; 
        10'b0000110100: data <= 10'h001; 
        10'b0000110101: data <= 10'h001; 
        10'b0000110110: data <= 10'h000; 
        10'b0000110111: data <= 10'h001; 
        10'b0000111000: data <= 10'h001; 
        10'b0000111001: data <= 10'h001; 
        10'b0000111010: data <= 10'h001; 
        10'b0000111011: data <= 10'h001; 
        10'b0000111100: data <= 10'h001; 
        10'b0000111101: data <= 10'h001; 
        10'b0000111110: data <= 10'h001; 
        10'b0000111111: data <= 10'h000; 
        10'b0001000000: data <= 10'h000; 
        10'b0001000001: data <= 10'h000; 
        10'b0001000010: data <= 10'h000; 
        10'b0001000011: data <= 10'h3ff; 
        10'b0001000100: data <= 10'h3fe; 
        10'b0001000101: data <= 10'h3ff; 
        10'b0001000110: data <= 10'h3ff; 
        10'b0001000111: data <= 10'h3ff; 
        10'b0001001000: data <= 10'h3ff; 
        10'b0001001001: data <= 10'h000; 
        10'b0001001010: data <= 10'h000; 
        10'b0001001011: data <= 10'h001; 
        10'b0001001100: data <= 10'h001; 
        10'b0001001101: data <= 10'h001; 
        10'b0001001110: data <= 10'h001; 
        10'b0001001111: data <= 10'h000; 
        10'b0001010000: data <= 10'h000; 
        10'b0001010001: data <= 10'h001; 
        10'b0001010010: data <= 10'h000; 
        10'b0001010011: data <= 10'h000; 
        10'b0001010100: data <= 10'h001; 
        10'b0001010101: data <= 10'h001; 
        10'b0001010110: data <= 10'h000; 
        10'b0001010111: data <= 10'h000; 
        10'b0001011000: data <= 10'h000; 
        10'b0001011001: data <= 10'h000; 
        10'b0001011010: data <= 10'h001; 
        10'b0001011011: data <= 10'h3ff; 
        10'b0001011100: data <= 10'h3ff; 
        10'b0001011101: data <= 10'h000; 
        10'b0001011110: data <= 10'h3fe; 
        10'b0001011111: data <= 10'h3fe; 
        10'b0001100000: data <= 10'h3fd; 
        10'b0001100001: data <= 10'h3fd; 
        10'b0001100010: data <= 10'h3fd; 
        10'b0001100011: data <= 10'h3fc; 
        10'b0001100100: data <= 10'h3fd; 
        10'b0001100101: data <= 10'h3ff; 
        10'b0001100110: data <= 10'h000; 
        10'b0001100111: data <= 10'h000; 
        10'b0001101000: data <= 10'h001; 
        10'b0001101001: data <= 10'h001; 
        10'b0001101010: data <= 10'h000; 
        10'b0001101011: data <= 10'h000; 
        10'b0001101100: data <= 10'h001; 
        10'b0001101101: data <= 10'h001; 
        10'b0001101110: data <= 10'h000; 
        10'b0001101111: data <= 10'h001; 
        10'b0001110000: data <= 10'h001; 
        10'b0001110001: data <= 10'h001; 
        10'b0001110010: data <= 10'h001; 
        10'b0001110011: data <= 10'h001; 
        10'b0001110100: data <= 10'h000; 
        10'b0001110101: data <= 10'h001; 
        10'b0001110110: data <= 10'h3ff; 
        10'b0001110111: data <= 10'h000; 
        10'b0001111000: data <= 10'h3ff; 
        10'b0001111001: data <= 10'h3ff; 
        10'b0001111010: data <= 10'h3fd; 
        10'b0001111011: data <= 10'h3fd; 
        10'b0001111100: data <= 10'h3fc; 
        10'b0001111101: data <= 10'h3fd; 
        10'b0001111110: data <= 10'h3fc; 
        10'b0001111111: data <= 10'h3fc; 
        10'b0010000000: data <= 10'h3fe; 
        10'b0010000001: data <= 10'h3fe; 
        10'b0010000010: data <= 10'h3ff; 
        10'b0010000011: data <= 10'h001; 
        10'b0010000100: data <= 10'h001; 
        10'b0010000101: data <= 10'h001; 
        10'b0010000110: data <= 10'h001; 
        10'b0010000111: data <= 10'h002; 
        10'b0010001000: data <= 10'h000; 
        10'b0010001001: data <= 10'h001; 
        10'b0010001010: data <= 10'h000; 
        10'b0010001011: data <= 10'h000; 
        10'b0010001100: data <= 10'h001; 
        10'b0010001101: data <= 10'h000; 
        10'b0010001110: data <= 10'h001; 
        10'b0010001111: data <= 10'h000; 
        10'b0010010000: data <= 10'h001; 
        10'b0010010001: data <= 10'h000; 
        10'b0010010010: data <= 10'h000; 
        10'b0010010011: data <= 10'h3ff; 
        10'b0010010100: data <= 10'h000; 
        10'b0010010101: data <= 10'h3ff; 
        10'b0010010110: data <= 10'h3fe; 
        10'b0010010111: data <= 10'h3fe; 
        10'b0010011000: data <= 10'h3fd; 
        10'b0010011001: data <= 10'h3fd; 
        10'b0010011010: data <= 10'h3fe; 
        10'b0010011011: data <= 10'h3fe; 
        10'b0010011100: data <= 10'h000; 
        10'b0010011101: data <= 10'h000; 
        10'b0010011110: data <= 10'h000; 
        10'b0010011111: data <= 10'h001; 
        10'b0010100000: data <= 10'h001; 
        10'b0010100001: data <= 10'h001; 
        10'b0010100010: data <= 10'h003; 
        10'b0010100011: data <= 10'h003; 
        10'b0010100100: data <= 10'h002; 
        10'b0010100101: data <= 10'h000; 
        10'b0010100110: data <= 10'h000; 
        10'b0010100111: data <= 10'h000; 
        10'b0010101000: data <= 10'h001; 
        10'b0010101001: data <= 10'h001; 
        10'b0010101010: data <= 10'h000; 
        10'b0010101011: data <= 10'h001; 
        10'b0010101100: data <= 10'h001; 
        10'b0010101101: data <= 10'h001; 
        10'b0010101110: data <= 10'h001; 
        10'b0010101111: data <= 10'h000; 
        10'b0010110000: data <= 10'h000; 
        10'b0010110001: data <= 10'h3ff; 
        10'b0010110010: data <= 10'h3fe; 
        10'b0010110011: data <= 10'h3fd; 
        10'b0010110100: data <= 10'h3fb; 
        10'b0010110101: data <= 10'h3fa; 
        10'b0010110110: data <= 10'h3fa; 
        10'b0010110111: data <= 10'h3fb; 
        10'b0010111000: data <= 10'h3fb; 
        10'b0010111001: data <= 10'h3fd; 
        10'b0010111010: data <= 10'h3fd; 
        10'b0010111011: data <= 10'h3ff; 
        10'b0010111100: data <= 10'h3ff; 
        10'b0010111101: data <= 10'h000; 
        10'b0010111110: data <= 10'h004; 
        10'b0010111111: data <= 10'h004; 
        10'b0011000000: data <= 10'h002; 
        10'b0011000001: data <= 10'h001; 
        10'b0011000010: data <= 10'h001; 
        10'b0011000011: data <= 10'h000; 
        10'b0011000100: data <= 10'h000; 
        10'b0011000101: data <= 10'h000; 
        10'b0011000110: data <= 10'h000; 
        10'b0011000111: data <= 10'h001; 
        10'b0011001000: data <= 10'h000; 
        10'b0011001001: data <= 10'h001; 
        10'b0011001010: data <= 10'h000; 
        10'b0011001011: data <= 10'h000; 
        10'b0011001100: data <= 10'h3ff; 
        10'b0011001101: data <= 10'h3ff; 
        10'b0011001110: data <= 10'h3fd; 
        10'b0011001111: data <= 10'h3fb; 
        10'b0011010000: data <= 10'h3fa; 
        10'b0011010001: data <= 10'h3fc; 
        10'b0011010010: data <= 10'h3fa; 
        10'b0011010011: data <= 10'h3fa; 
        10'b0011010100: data <= 10'h3fa; 
        10'b0011010101: data <= 10'h3fc; 
        10'b0011010110: data <= 10'h3fc; 
        10'b0011010111: data <= 10'h3fd; 
        10'b0011011000: data <= 10'h3fd; 
        10'b0011011001: data <= 10'h3ff; 
        10'b0011011010: data <= 10'h003; 
        10'b0011011011: data <= 10'h003; 
        10'b0011011100: data <= 10'h002; 
        10'b0011011101: data <= 10'h001; 
        10'b0011011110: data <= 10'h001; 
        10'b0011011111: data <= 10'h001; 
        10'b0011100000: data <= 10'h001; 
        10'b0011100001: data <= 10'h001; 
        10'b0011100010: data <= 10'h001; 
        10'b0011100011: data <= 10'h000; 
        10'b0011100100: data <= 10'h000; 
        10'b0011100101: data <= 10'h000; 
        10'b0011100110: data <= 10'h000; 
        10'b0011100111: data <= 10'h000; 
        10'b0011101000: data <= 10'h3fe; 
        10'b0011101001: data <= 10'h3ff; 
        10'b0011101010: data <= 10'h3fe; 
        10'b0011101011: data <= 10'h3fd; 
        10'b0011101100: data <= 10'h3fb; 
        10'b0011101101: data <= 10'h3fd; 
        10'b0011101110: data <= 10'h3f9; 
        10'b0011101111: data <= 10'h3f9; 
        10'b0011110000: data <= 10'h3fb; 
        10'b0011110001: data <= 10'h3fd; 
        10'b0011110010: data <= 10'h3fd; 
        10'b0011110011: data <= 10'h3ff; 
        10'b0011110100: data <= 10'h3fe; 
        10'b0011110101: data <= 10'h3fe; 
        10'b0011110110: data <= 10'h001; 
        10'b0011110111: data <= 10'h002; 
        10'b0011111000: data <= 10'h001; 
        10'b0011111001: data <= 10'h000; 
        10'b0011111010: data <= 10'h000; 
        10'b0011111011: data <= 10'h001; 
        10'b0011111100: data <= 10'h001; 
        10'b0011111101: data <= 10'h001; 
        10'b0011111110: data <= 10'h001; 
        10'b0011111111: data <= 10'h000; 
        10'b0100000000: data <= 10'h3ff; 
        10'b0100000001: data <= 10'h000; 
        10'b0100000010: data <= 10'h3ff; 
        10'b0100000011: data <= 10'h3ff; 
        10'b0100000100: data <= 10'h3ff; 
        10'b0100000101: data <= 10'h000; 
        10'b0100000110: data <= 10'h3ff; 
        10'b0100000111: data <= 10'h3ff; 
        10'b0100001000: data <= 10'h3ff; 
        10'b0100001001: data <= 10'h3fd; 
        10'b0100001010: data <= 10'h3f7; 
        10'b0100001011: data <= 10'h3f9; 
        10'b0100001100: data <= 10'h3fe; 
        10'b0100001101: data <= 10'h3ff; 
        10'b0100001110: data <= 10'h000; 
        10'b0100001111: data <= 10'h000; 
        10'b0100010000: data <= 10'h3ff; 
        10'b0100010001: data <= 10'h3ff; 
        10'b0100010010: data <= 10'h000; 
        10'b0100010011: data <= 10'h000; 
        10'b0100010100: data <= 10'h3ff; 
        10'b0100010101: data <= 10'h3ff; 
        10'b0100010110: data <= 10'h3ff; 
        10'b0100010111: data <= 10'h001; 
        10'b0100011000: data <= 10'h001; 
        10'b0100011001: data <= 10'h000; 
        10'b0100011010: data <= 10'h000; 
        10'b0100011011: data <= 10'h000; 
        10'b0100011100: data <= 10'h000; 
        10'b0100011101: data <= 10'h3ff; 
        10'b0100011110: data <= 10'h3fe; 
        10'b0100011111: data <= 10'h3ff; 
        10'b0100100000: data <= 10'h000; 
        10'b0100100001: data <= 10'h003; 
        10'b0100100010: data <= 10'h002; 
        10'b0100100011: data <= 10'h001; 
        10'b0100100100: data <= 10'h001; 
        10'b0100100101: data <= 10'h3fc; 
        10'b0100100110: data <= 10'h3f6; 
        10'b0100100111: data <= 10'h3fd; 
        10'b0100101000: data <= 10'h000; 
        10'b0100101001: data <= 10'h000; 
        10'b0100101010: data <= 10'h000; 
        10'b0100101011: data <= 10'h000; 
        10'b0100101100: data <= 10'h3fe; 
        10'b0100101101: data <= 10'h3ff; 
        10'b0100101110: data <= 10'h000; 
        10'b0100101111: data <= 10'h3fe; 
        10'b0100110000: data <= 10'h3ff; 
        10'b0100110001: data <= 10'h3ff; 
        10'b0100110010: data <= 10'h001; 
        10'b0100110011: data <= 10'h001; 
        10'b0100110100: data <= 10'h001; 
        10'b0100110101: data <= 10'h001; 
        10'b0100110110: data <= 10'h001; 
        10'b0100110111: data <= 10'h000; 
        10'b0100111000: data <= 10'h000; 
        10'b0100111001: data <= 10'h3ff; 
        10'b0100111010: data <= 10'h3ff; 
        10'b0100111011: data <= 10'h001; 
        10'b0100111100: data <= 10'h002; 
        10'b0100111101: data <= 10'h003; 
        10'b0100111110: data <= 10'h005; 
        10'b0100111111: data <= 10'h003; 
        10'b0101000000: data <= 10'h003; 
        10'b0101000001: data <= 10'h3fa; 
        10'b0101000010: data <= 10'h3f8; 
        10'b0101000011: data <= 10'h001; 
        10'b0101000100: data <= 10'h004; 
        10'b0101000101: data <= 10'h001; 
        10'b0101000110: data <= 10'h000; 
        10'b0101000111: data <= 10'h3ff; 
        10'b0101001000: data <= 10'h3fe; 
        10'b0101001001: data <= 10'h3fe; 
        10'b0101001010: data <= 10'h3ff; 
        10'b0101001011: data <= 10'h3fe; 
        10'b0101001100: data <= 10'h3fe; 
        10'b0101001101: data <= 10'h000; 
        10'b0101001110: data <= 10'h000; 
        10'b0101001111: data <= 10'h000; 
        10'b0101010000: data <= 10'h001; 
        10'b0101010001: data <= 10'h001; 
        10'b0101010010: data <= 10'h000; 
        10'b0101010011: data <= 10'h000; 
        10'b0101010100: data <= 10'h000; 
        10'b0101010101: data <= 10'h3ff; 
        10'b0101010110: data <= 10'h002; 
        10'b0101010111: data <= 10'h003; 
        10'b0101011000: data <= 10'h005; 
        10'b0101011001: data <= 10'h004; 
        10'b0101011010: data <= 10'h007; 
        10'b0101011011: data <= 10'h008; 
        10'b0101011100: data <= 10'h008; 
        10'b0101011101: data <= 10'h000; 
        10'b0101011110: data <= 10'h3fc; 
        10'b0101011111: data <= 10'h003; 
        10'b0101100000: data <= 10'h005; 
        10'b0101100001: data <= 10'h001; 
        10'b0101100010: data <= 10'h000; 
        10'b0101100011: data <= 10'h001; 
        10'b0101100100: data <= 10'h000; 
        10'b0101100101: data <= 10'h000; 
        10'b0101100110: data <= 10'h000; 
        10'b0101100111: data <= 10'h3ff; 
        10'b0101101000: data <= 10'h3ff; 
        10'b0101101001: data <= 10'h000; 
        10'b0101101010: data <= 10'h001; 
        10'b0101101011: data <= 10'h001; 
        10'b0101101100: data <= 10'h000; 
        10'b0101101101: data <= 10'h001; 
        10'b0101101110: data <= 10'h000; 
        10'b0101101111: data <= 10'h000; 
        10'b0101110000: data <= 10'h001; 
        10'b0101110001: data <= 10'h002; 
        10'b0101110010: data <= 10'h005; 
        10'b0101110011: data <= 10'h006; 
        10'b0101110100: data <= 10'h007; 
        10'b0101110101: data <= 10'h005; 
        10'b0101110110: data <= 10'h006; 
        10'b0101110111: data <= 10'h00a; 
        10'b0101111000: data <= 10'h008; 
        10'b0101111001: data <= 10'h000; 
        10'b0101111010: data <= 10'h3ff; 
        10'b0101111011: data <= 10'h004; 
        10'b0101111100: data <= 10'h004; 
        10'b0101111101: data <= 10'h004; 
        10'b0101111110: data <= 10'h003; 
        10'b0101111111: data <= 10'h001; 
        10'b0110000000: data <= 10'h003; 
        10'b0110000001: data <= 10'h002; 
        10'b0110000010: data <= 10'h001; 
        10'b0110000011: data <= 10'h3ff; 
        10'b0110000100: data <= 10'h3ff; 
        10'b0110000101: data <= 10'h000; 
        10'b0110000110: data <= 10'h001; 
        10'b0110000111: data <= 10'h001; 
        10'b0110001000: data <= 10'h000; 
        10'b0110001001: data <= 10'h001; 
        10'b0110001010: data <= 10'h000; 
        10'b0110001011: data <= 10'h001; 
        10'b0110001100: data <= 10'h002; 
        10'b0110001101: data <= 10'h004; 
        10'b0110001110: data <= 10'h006; 
        10'b0110001111: data <= 10'h007; 
        10'b0110010000: data <= 10'h005; 
        10'b0110010001: data <= 10'h005; 
        10'b0110010010: data <= 10'h006; 
        10'b0110010011: data <= 10'h007; 
        10'b0110010100: data <= 10'h005; 
        10'b0110010101: data <= 10'h000; 
        10'b0110010110: data <= 10'h3ff; 
        10'b0110010111: data <= 10'h001; 
        10'b0110011000: data <= 10'h004; 
        10'b0110011001: data <= 10'h007; 
        10'b0110011010: data <= 10'h005; 
        10'b0110011011: data <= 10'h004; 
        10'b0110011100: data <= 10'h002; 
        10'b0110011101: data <= 10'h002; 
        10'b0110011110: data <= 10'h001; 
        10'b0110011111: data <= 10'h000; 
        10'b0110100000: data <= 10'h000; 
        10'b0110100001: data <= 10'h000; 
        10'b0110100010: data <= 10'h001; 
        10'b0110100011: data <= 10'h000; 
        10'b0110100100: data <= 10'h001; 
        10'b0110100101: data <= 10'h001; 
        10'b0110100110: data <= 10'h001; 
        10'b0110100111: data <= 10'h001; 
        10'b0110101000: data <= 10'h002; 
        10'b0110101001: data <= 10'h002; 
        10'b0110101010: data <= 10'h003; 
        10'b0110101011: data <= 10'h003; 
        10'b0110101100: data <= 10'h005; 
        10'b0110101101: data <= 10'h004; 
        10'b0110101110: data <= 10'h003; 
        10'b0110101111: data <= 10'h002; 
        10'b0110110000: data <= 10'h003; 
        10'b0110110001: data <= 10'h001; 
        10'b0110110010: data <= 10'h002; 
        10'b0110110011: data <= 10'h003; 
        10'b0110110100: data <= 10'h006; 
        10'b0110110101: data <= 10'h005; 
        10'b0110110110: data <= 10'h004; 
        10'b0110110111: data <= 10'h002; 
        10'b0110111000: data <= 10'h3ff; 
        10'b0110111001: data <= 10'h001; 
        10'b0110111010: data <= 10'h002; 
        10'b0110111011: data <= 10'h000; 
        10'b0110111100: data <= 10'h3ff; 
        10'b0110111101: data <= 10'h000; 
        10'b0110111110: data <= 10'h000; 
        10'b0110111111: data <= 10'h000; 
        10'b0111000000: data <= 10'h000; 
        10'b0111000001: data <= 10'h000; 
        10'b0111000010: data <= 10'h000; 
        10'b0111000011: data <= 10'h000; 
        10'b0111000100: data <= 10'h001; 
        10'b0111000101: data <= 10'h001; 
        10'b0111000110: data <= 10'h002; 
        10'b0111000111: data <= 10'h004; 
        10'b0111001000: data <= 10'h005; 
        10'b0111001001: data <= 10'h004; 
        10'b0111001010: data <= 10'h001; 
        10'b0111001011: data <= 10'h000; 
        10'b0111001100: data <= 10'h001; 
        10'b0111001101: data <= 10'h001; 
        10'b0111001110: data <= 10'h005; 
        10'b0111001111: data <= 10'h007; 
        10'b0111010000: data <= 10'h007; 
        10'b0111010001: data <= 10'h006; 
        10'b0111010010: data <= 10'h004; 
        10'b0111010011: data <= 10'h000; 
        10'b0111010100: data <= 10'h002; 
        10'b0111010101: data <= 10'h002; 
        10'b0111010110: data <= 10'h001; 
        10'b0111010111: data <= 10'h000; 
        10'b0111011000: data <= 10'h000; 
        10'b0111011001: data <= 10'h000; 
        10'b0111011010: data <= 10'h000; 
        10'b0111011011: data <= 10'h000; 
        10'b0111011100: data <= 10'h000; 
        10'b0111011101: data <= 10'h000; 
        10'b0111011110: data <= 10'h001; 
        10'b0111011111: data <= 10'h000; 
        10'b0111100000: data <= 10'h3ff; 
        10'b0111100001: data <= 10'h3ff; 
        10'b0111100010: data <= 10'h001; 
        10'b0111100011: data <= 10'h003; 
        10'b0111100100: data <= 10'h006; 
        10'b0111100101: data <= 10'h005; 
        10'b0111100110: data <= 10'h002; 
        10'b0111100111: data <= 10'h001; 
        10'b0111101000: data <= 10'h002; 
        10'b0111101001: data <= 10'h005; 
        10'b0111101010: data <= 10'h008; 
        10'b0111101011: data <= 10'h006; 
        10'b0111101100: data <= 10'h005; 
        10'b0111101101: data <= 10'h002; 
        10'b0111101110: data <= 10'h000; 
        10'b0111101111: data <= 10'h3fe; 
        10'b0111110000: data <= 10'h001; 
        10'b0111110001: data <= 10'h000; 
        10'b0111110010: data <= 10'h3ff; 
        10'b0111110011: data <= 10'h000; 
        10'b0111110100: data <= 10'h3ff; 
        10'b0111110101: data <= 10'h000; 
        10'b0111110110: data <= 10'h001; 
        10'b0111110111: data <= 10'h001; 
        10'b0111111000: data <= 10'h000; 
        10'b0111111001: data <= 10'h001; 
        10'b0111111010: data <= 10'h001; 
        10'b0111111011: data <= 10'h000; 
        10'b0111111100: data <= 10'h3ff; 
        10'b0111111101: data <= 10'h3ff; 
        10'b0111111110: data <= 10'h3fe; 
        10'b0111111111: data <= 10'h000; 
        10'b1000000000: data <= 10'h001; 
        10'b1000000001: data <= 10'h000; 
        10'b1000000010: data <= 10'h3ff; 
        10'b1000000011: data <= 10'h3ff; 
        10'b1000000100: data <= 10'h002; 
        10'b1000000101: data <= 10'h002; 
        10'b1000000110: data <= 10'h004; 
        10'b1000000111: data <= 10'h003; 
        10'b1000001000: data <= 10'h002; 
        10'b1000001001: data <= 10'h3fe; 
        10'b1000001010: data <= 10'h3fe; 
        10'b1000001011: data <= 10'h3fd; 
        10'b1000001100: data <= 10'h3fe; 
        10'b1000001101: data <= 10'h3fe; 
        10'b1000001110: data <= 10'h3fd; 
        10'b1000001111: data <= 10'h3fe; 
        10'b1000010000: data <= 10'h3ff; 
        10'b1000010001: data <= 10'h000; 
        10'b1000010010: data <= 10'h000; 
        10'b1000010011: data <= 10'h000; 
        10'b1000010100: data <= 10'h000; 
        10'b1000010101: data <= 10'h001; 
        10'b1000010110: data <= 10'h000; 
        10'b1000010111: data <= 10'h000; 
        10'b1000011000: data <= 10'h3fe; 
        10'b1000011001: data <= 10'h3fe; 
        10'b1000011010: data <= 10'h3fd; 
        10'b1000011011: data <= 10'h3fc; 
        10'b1000011100: data <= 10'h3fc; 
        10'b1000011101: data <= 10'h3fb; 
        10'b1000011110: data <= 10'h3fb; 
        10'b1000011111: data <= 10'h3fb; 
        10'b1000100000: data <= 10'h3fb; 
        10'b1000100001: data <= 10'h3fd; 
        10'b1000100010: data <= 10'h3ff; 
        10'b1000100011: data <= 10'h001; 
        10'b1000100100: data <= 10'h3fe; 
        10'b1000100101: data <= 10'h3fe; 
        10'b1000100110: data <= 10'h3fe; 
        10'b1000100111: data <= 10'h3fd; 
        10'b1000101000: data <= 10'h3fd; 
        10'b1000101001: data <= 10'h3fd; 
        10'b1000101010: data <= 10'h3fd; 
        10'b1000101011: data <= 10'h3fe; 
        10'b1000101100: data <= 10'h3ff; 
        10'b1000101101: data <= 10'h000; 
        10'b1000101110: data <= 10'h001; 
        10'b1000101111: data <= 10'h001; 
        10'b1000110000: data <= 10'h001; 
        10'b1000110001: data <= 10'h001; 
        10'b1000110010: data <= 10'h000; 
        10'b1000110011: data <= 10'h000; 
        10'b1000110100: data <= 10'h3ff; 
        10'b1000110101: data <= 10'h3fe; 
        10'b1000110110: data <= 10'h3fd; 
        10'b1000110111: data <= 10'h3fb; 
        10'b1000111000: data <= 10'h3fa; 
        10'b1000111001: data <= 10'h3fa; 
        10'b1000111010: data <= 10'h3f9; 
        10'b1000111011: data <= 10'h3fb; 
        10'b1000111100: data <= 10'h3fc; 
        10'b1000111101: data <= 10'h3fc; 
        10'b1000111110: data <= 10'h3fd; 
        10'b1000111111: data <= 10'h3ff; 
        10'b1001000000: data <= 10'h000; 
        10'b1001000001: data <= 10'h000; 
        10'b1001000010: data <= 10'h3ff; 
        10'b1001000011: data <= 10'h3fe; 
        10'b1001000100: data <= 10'h3fe; 
        10'b1001000101: data <= 10'h3fe; 
        10'b1001000110: data <= 10'h3fe; 
        10'b1001000111: data <= 10'h3ff; 
        10'b1001001000: data <= 10'h3ff; 
        10'b1001001001: data <= 10'h000; 
        10'b1001001010: data <= 10'h000; 
        10'b1001001011: data <= 10'h001; 
        10'b1001001100: data <= 10'h000; 
        10'b1001001101: data <= 10'h000; 
        10'b1001001110: data <= 10'h000; 
        10'b1001001111: data <= 10'h000; 
        10'b1001010000: data <= 10'h000; 
        10'b1001010001: data <= 10'h3ff; 
        10'b1001010010: data <= 10'h3fd; 
        10'b1001010011: data <= 10'h3fc; 
        10'b1001010100: data <= 10'h3fc; 
        10'b1001010101: data <= 10'h3fc; 
        10'b1001010110: data <= 10'h3fc; 
        10'b1001010111: data <= 10'h3fd; 
        10'b1001011000: data <= 10'h3fe; 
        10'b1001011001: data <= 10'h3fe; 
        10'b1001011010: data <= 10'h3fd; 
        10'b1001011011: data <= 10'h3ff; 
        10'b1001011100: data <= 10'h3fe; 
        10'b1001011101: data <= 10'h000; 
        10'b1001011110: data <= 10'h000; 
        10'b1001011111: data <= 10'h000; 
        10'b1001100000: data <= 10'h000; 
        10'b1001100001: data <= 10'h3fe; 
        10'b1001100010: data <= 10'h3ff; 
        10'b1001100011: data <= 10'h000; 
        10'b1001100100: data <= 10'h000; 
        10'b1001100101: data <= 10'h000; 
        10'b1001100110: data <= 10'h001; 
        10'b1001100111: data <= 10'h001; 
        10'b1001101000: data <= 10'h001; 
        10'b1001101001: data <= 10'h001; 
        10'b1001101010: data <= 10'h000; 
        10'b1001101011: data <= 10'h001; 
        10'b1001101100: data <= 10'h000; 
        10'b1001101101: data <= 10'h3ff; 
        10'b1001101110: data <= 10'h3ff; 
        10'b1001101111: data <= 10'h3fe; 
        10'b1001110000: data <= 10'h3fd; 
        10'b1001110001: data <= 10'h3fe; 
        10'b1001110010: data <= 10'h3fe; 
        10'b1001110011: data <= 10'h3ff; 
        10'b1001110100: data <= 10'h3ff; 
        10'b1001110101: data <= 10'h3ff; 
        10'b1001110110: data <= 10'h3ff; 
        10'b1001110111: data <= 10'h3ff; 
        10'b1001111000: data <= 10'h3ff; 
        10'b1001111001: data <= 10'h000; 
        10'b1001111010: data <= 10'h001; 
        10'b1001111011: data <= 10'h002; 
        10'b1001111100: data <= 10'h002; 
        10'b1001111101: data <= 10'h001; 
        10'b1001111110: data <= 10'h3ff; 
        10'b1001111111: data <= 10'h3ff; 
        10'b1010000000: data <= 10'h000; 
        10'b1010000001: data <= 10'h000; 
        10'b1010000010: data <= 10'h000; 
        10'b1010000011: data <= 10'h000; 
        10'b1010000100: data <= 10'h000; 
        10'b1010000101: data <= 10'h000; 
        10'b1010000110: data <= 10'h000; 
        10'b1010000111: data <= 10'h001; 
        10'b1010001000: data <= 10'h000; 
        10'b1010001001: data <= 10'h000; 
        10'b1010001010: data <= 10'h3ff; 
        10'b1010001011: data <= 10'h3ff; 
        10'b1010001100: data <= 10'h3ff; 
        10'b1010001101: data <= 10'h000; 
        10'b1010001110: data <= 10'h3ff; 
        10'b1010001111: data <= 10'h000; 
        10'b1010010000: data <= 10'h3ff; 
        10'b1010010001: data <= 10'h3ff; 
        10'b1010010010: data <= 10'h3ff; 
        10'b1010010011: data <= 10'h000; 
        10'b1010010100: data <= 10'h000; 
        10'b1010010101: data <= 10'h001; 
        10'b1010010110: data <= 10'h002; 
        10'b1010010111: data <= 10'h002; 
        10'b1010011000: data <= 10'h002; 
        10'b1010011001: data <= 10'h001; 
        10'b1010011010: data <= 10'h000; 
        10'b1010011011: data <= 10'h000; 
        10'b1010011100: data <= 10'h001; 
        10'b1010011101: data <= 10'h001; 
        10'b1010011110: data <= 10'h000; 
        10'b1010011111: data <= 10'h001; 
        10'b1010100000: data <= 10'h001; 
        10'b1010100001: data <= 10'h001; 
        10'b1010100010: data <= 10'h000; 
        10'b1010100011: data <= 10'h001; 
        10'b1010100100: data <= 10'h000; 
        10'b1010100101: data <= 10'h001; 
        10'b1010100110: data <= 10'h000; 
        10'b1010100111: data <= 10'h3ff; 
        10'b1010101000: data <= 10'h3ff; 
        10'b1010101001: data <= 10'h000; 
        10'b1010101010: data <= 10'h3ff; 
        10'b1010101011: data <= 10'h000; 
        10'b1010101100: data <= 10'h3ff; 
        10'b1010101101: data <= 10'h3ff; 
        10'b1010101110: data <= 10'h3ff; 
        10'b1010101111: data <= 10'h3fe; 
        10'b1010110000: data <= 10'h3ff; 
        10'b1010110001: data <= 10'h000; 
        10'b1010110010: data <= 10'h000; 
        10'b1010110011: data <= 10'h001; 
        10'b1010110100: data <= 10'h001; 
        10'b1010110101: data <= 10'h000; 
        10'b1010110110: data <= 10'h000; 
        10'b1010110111: data <= 10'h000; 
        10'b1010111000: data <= 10'h001; 
        10'b1010111001: data <= 10'h000; 
        10'b1010111010: data <= 10'h000; 
        10'b1010111011: data <= 10'h001; 
        10'b1010111100: data <= 10'h001; 
        10'b1010111101: data <= 10'h001; 
        10'b1010111110: data <= 10'h001; 
        10'b1010111111: data <= 10'h000; 
        10'b1011000000: data <= 10'h001; 
        10'b1011000001: data <= 10'h000; 
        10'b1011000010: data <= 10'h3ff; 
        10'b1011000011: data <= 10'h3ff; 
        10'b1011000100: data <= 10'h3fe; 
        10'b1011000101: data <= 10'h3fe; 
        10'b1011000110: data <= 10'h3fd; 
        10'b1011000111: data <= 10'h3fd; 
        10'b1011001000: data <= 10'h3fd; 
        10'b1011001001: data <= 10'h3fd; 
        10'b1011001010: data <= 10'h3fe; 
        10'b1011001011: data <= 10'h3fd; 
        10'b1011001100: data <= 10'h3fd; 
        10'b1011001101: data <= 10'h3fc; 
        10'b1011001110: data <= 10'h3fd; 
        10'b1011001111: data <= 10'h3fe; 
        10'b1011010000: data <= 10'h3fe; 
        10'b1011010001: data <= 10'h3ff; 
        10'b1011010010: data <= 10'h000; 
        10'b1011010011: data <= 10'h001; 
        10'b1011010100: data <= 10'h000; 
        10'b1011010101: data <= 10'h001; 
        10'b1011010110: data <= 10'h000; 
        10'b1011010111: data <= 10'h000; 
        10'b1011011000: data <= 10'h000; 
        10'b1011011001: data <= 10'h001; 
        10'b1011011010: data <= 10'h000; 
        10'b1011011011: data <= 10'h000; 
        10'b1011011100: data <= 10'h000; 
        10'b1011011101: data <= 10'h000; 
        10'b1011011110: data <= 10'h000; 
        10'b1011011111: data <= 10'h000; 
        10'b1011100000: data <= 10'h000; 
        10'b1011100001: data <= 10'h3ff; 
        10'b1011100010: data <= 10'h3fe; 
        10'b1011100011: data <= 10'h3fe; 
        10'b1011100100: data <= 10'h3fe; 
        10'b1011100101: data <= 10'h3fd; 
        10'b1011100110: data <= 10'h3fd; 
        10'b1011100111: data <= 10'h3fd; 
        10'b1011101000: data <= 10'h3fd; 
        10'b1011101001: data <= 10'h3fd; 
        10'b1011101010: data <= 10'h3fe; 
        10'b1011101011: data <= 10'h3ff; 
        10'b1011101100: data <= 10'h000; 
        10'b1011101101: data <= 10'h001; 
        10'b1011101110: data <= 10'h001; 
        10'b1011101111: data <= 10'h000; 
        10'b1011110000: data <= 10'h000; 
        10'b1011110001: data <= 10'h000; 
        10'b1011110010: data <= 10'h001; 
        10'b1011110011: data <= 10'h000; 
        10'b1011110100: data <= 10'h001; 
        10'b1011110101: data <= 10'h000; 
        10'b1011110110: data <= 10'h000; 
        10'b1011110111: data <= 10'h001; 
        10'b1011111000: data <= 10'h000; 
        10'b1011111001: data <= 10'h001; 
        10'b1011111010: data <= 10'h000; 
        10'b1011111011: data <= 10'h001; 
        10'b1011111100: data <= 10'h000; 
        10'b1011111101: data <= 10'h000; 
        10'b1011111110: data <= 10'h000; 
        10'b1011111111: data <= 10'h000; 
        10'b1100000000: data <= 10'h000; 
        10'b1100000001: data <= 10'h000; 
        10'b1100000010: data <= 10'h000; 
        10'b1100000011: data <= 10'h001; 
        10'b1100000100: data <= 10'h000; 
        10'b1100000101: data <= 10'h000; 
        10'b1100000110: data <= 10'h000; 
        10'b1100000111: data <= 10'h000; 
        10'b1100001000: data <= 10'h000; 
        10'b1100001001: data <= 10'h000; 
        10'b1100001010: data <= 10'h000; 
        10'b1100001011: data <= 10'h001; 
        10'b1100001100: data <= 10'h001; 
        10'b1100001101: data <= 10'h001; 
        10'b1100001110: data <= 10'h001; 
        10'b1100001111: data <= 10'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 5) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 11'h000; 
        10'b0000000001: data <= 11'h000; 
        10'b0000000010: data <= 11'h002; 
        10'b0000000011: data <= 11'h002; 
        10'b0000000100: data <= 11'h000; 
        10'b0000000101: data <= 11'h000; 
        10'b0000000110: data <= 11'h001; 
        10'b0000000111: data <= 11'h000; 
        10'b0000001000: data <= 11'h000; 
        10'b0000001001: data <= 11'h000; 
        10'b0000001010: data <= 11'h000; 
        10'b0000001011: data <= 11'h001; 
        10'b0000001100: data <= 11'h002; 
        10'b0000001101: data <= 11'h001; 
        10'b0000001110: data <= 11'h001; 
        10'b0000001111: data <= 11'h000; 
        10'b0000010000: data <= 11'h001; 
        10'b0000010001: data <= 11'h002; 
        10'b0000010010: data <= 11'h000; 
        10'b0000010011: data <= 11'h001; 
        10'b0000010100: data <= 11'h000; 
        10'b0000010101: data <= 11'h001; 
        10'b0000010110: data <= 11'h002; 
        10'b0000010111: data <= 11'h000; 
        10'b0000011000: data <= 11'h002; 
        10'b0000011001: data <= 11'h000; 
        10'b0000011010: data <= 11'h002; 
        10'b0000011011: data <= 11'h001; 
        10'b0000011100: data <= 11'h001; 
        10'b0000011101: data <= 11'h001; 
        10'b0000011110: data <= 11'h000; 
        10'b0000011111: data <= 11'h000; 
        10'b0000100000: data <= 11'h001; 
        10'b0000100001: data <= 11'h002; 
        10'b0000100010: data <= 11'h000; 
        10'b0000100011: data <= 11'h000; 
        10'b0000100100: data <= 11'h001; 
        10'b0000100101: data <= 11'h000; 
        10'b0000100110: data <= 11'h001; 
        10'b0000100111: data <= 11'h7ff; 
        10'b0000101000: data <= 11'h001; 
        10'b0000101001: data <= 11'h7ff; 
        10'b0000101010: data <= 11'h000; 
        10'b0000101011: data <= 11'h001; 
        10'b0000101100: data <= 11'h001; 
        10'b0000101101: data <= 11'h000; 
        10'b0000101110: data <= 11'h000; 
        10'b0000101111: data <= 11'h000; 
        10'b0000110000: data <= 11'h002; 
        10'b0000110001: data <= 11'h000; 
        10'b0000110010: data <= 11'h000; 
        10'b0000110011: data <= 11'h000; 
        10'b0000110100: data <= 11'h001; 
        10'b0000110101: data <= 11'h001; 
        10'b0000110110: data <= 11'h000; 
        10'b0000110111: data <= 11'h001; 
        10'b0000111000: data <= 11'h002; 
        10'b0000111001: data <= 11'h001; 
        10'b0000111010: data <= 11'h002; 
        10'b0000111011: data <= 11'h002; 
        10'b0000111100: data <= 11'h002; 
        10'b0000111101: data <= 11'h001; 
        10'b0000111110: data <= 11'h002; 
        10'b0000111111: data <= 11'h7ff; 
        10'b0001000000: data <= 11'h7ff; 
        10'b0001000001: data <= 11'h000; 
        10'b0001000010: data <= 11'h000; 
        10'b0001000011: data <= 11'h7ff; 
        10'b0001000100: data <= 11'h7fc; 
        10'b0001000101: data <= 11'h7fe; 
        10'b0001000110: data <= 11'h7fe; 
        10'b0001000111: data <= 11'h7fd; 
        10'b0001001000: data <= 11'h7fe; 
        10'b0001001001: data <= 11'h000; 
        10'b0001001010: data <= 11'h001; 
        10'b0001001011: data <= 11'h002; 
        10'b0001001100: data <= 11'h002; 
        10'b0001001101: data <= 11'h001; 
        10'b0001001110: data <= 11'h002; 
        10'b0001001111: data <= 11'h000; 
        10'b0001010000: data <= 11'h001; 
        10'b0001010001: data <= 11'h001; 
        10'b0001010010: data <= 11'h000; 
        10'b0001010011: data <= 11'h001; 
        10'b0001010100: data <= 11'h002; 
        10'b0001010101: data <= 11'h001; 
        10'b0001010110: data <= 11'h001; 
        10'b0001010111: data <= 11'h001; 
        10'b0001011000: data <= 11'h001; 
        10'b0001011001: data <= 11'h000; 
        10'b0001011010: data <= 11'h001; 
        10'b0001011011: data <= 11'h7ff; 
        10'b0001011100: data <= 11'h7fe; 
        10'b0001011101: data <= 11'h7ff; 
        10'b0001011110: data <= 11'h7fc; 
        10'b0001011111: data <= 11'h7fc; 
        10'b0001100000: data <= 11'h7f9; 
        10'b0001100001: data <= 11'h7f9; 
        10'b0001100010: data <= 11'h7fa; 
        10'b0001100011: data <= 11'h7f8; 
        10'b0001100100: data <= 11'h7fb; 
        10'b0001100101: data <= 11'h7fd; 
        10'b0001100110: data <= 11'h000; 
        10'b0001100111: data <= 11'h001; 
        10'b0001101000: data <= 11'h001; 
        10'b0001101001: data <= 11'h002; 
        10'b0001101010: data <= 11'h001; 
        10'b0001101011: data <= 11'h001; 
        10'b0001101100: data <= 11'h002; 
        10'b0001101101: data <= 11'h002; 
        10'b0001101110: data <= 11'h001; 
        10'b0001101111: data <= 11'h001; 
        10'b0001110000: data <= 11'h002; 
        10'b0001110001: data <= 11'h001; 
        10'b0001110010: data <= 11'h002; 
        10'b0001110011: data <= 11'h001; 
        10'b0001110100: data <= 11'h001; 
        10'b0001110101: data <= 11'h002; 
        10'b0001110110: data <= 11'h7ff; 
        10'b0001110111: data <= 11'h000; 
        10'b0001111000: data <= 11'h7fd; 
        10'b0001111001: data <= 11'h7fe; 
        10'b0001111010: data <= 11'h7fa; 
        10'b0001111011: data <= 11'h7fa; 
        10'b0001111100: data <= 11'h7f8; 
        10'b0001111101: data <= 11'h7f9; 
        10'b0001111110: data <= 11'h7f8; 
        10'b0001111111: data <= 11'h7f9; 
        10'b0010000000: data <= 11'h7fd; 
        10'b0010000001: data <= 11'h7fd; 
        10'b0010000010: data <= 11'h7fe; 
        10'b0010000011: data <= 11'h002; 
        10'b0010000100: data <= 11'h002; 
        10'b0010000101: data <= 11'h003; 
        10'b0010000110: data <= 11'h003; 
        10'b0010000111: data <= 11'h003; 
        10'b0010001000: data <= 11'h001; 
        10'b0010001001: data <= 11'h002; 
        10'b0010001010: data <= 11'h000; 
        10'b0010001011: data <= 11'h000; 
        10'b0010001100: data <= 11'h002; 
        10'b0010001101: data <= 11'h001; 
        10'b0010001110: data <= 11'h001; 
        10'b0010001111: data <= 11'h000; 
        10'b0010010000: data <= 11'h001; 
        10'b0010010001: data <= 11'h000; 
        10'b0010010010: data <= 11'h001; 
        10'b0010010011: data <= 11'h7ff; 
        10'b0010010100: data <= 11'h000; 
        10'b0010010101: data <= 11'h7ff; 
        10'b0010010110: data <= 11'h7fb; 
        10'b0010010111: data <= 11'h7fd; 
        10'b0010011000: data <= 11'h7fb; 
        10'b0010011001: data <= 11'h7fa; 
        10'b0010011010: data <= 11'h7fc; 
        10'b0010011011: data <= 11'h7fc; 
        10'b0010011100: data <= 11'h7ff; 
        10'b0010011101: data <= 11'h001; 
        10'b0010011110: data <= 11'h7ff; 
        10'b0010011111: data <= 11'h001; 
        10'b0010100000: data <= 11'h002; 
        10'b0010100001: data <= 11'h002; 
        10'b0010100010: data <= 11'h006; 
        10'b0010100011: data <= 11'h007; 
        10'b0010100100: data <= 11'h004; 
        10'b0010100101: data <= 11'h000; 
        10'b0010100110: data <= 11'h001; 
        10'b0010100111: data <= 11'h000; 
        10'b0010101000: data <= 11'h002; 
        10'b0010101001: data <= 11'h002; 
        10'b0010101010: data <= 11'h001; 
        10'b0010101011: data <= 11'h002; 
        10'b0010101100: data <= 11'h002; 
        10'b0010101101: data <= 11'h002; 
        10'b0010101110: data <= 11'h001; 
        10'b0010101111: data <= 11'h000; 
        10'b0010110000: data <= 11'h000; 
        10'b0010110001: data <= 11'h7fe; 
        10'b0010110010: data <= 11'h7fc; 
        10'b0010110011: data <= 11'h7fa; 
        10'b0010110100: data <= 11'h7f6; 
        10'b0010110101: data <= 11'h7f5; 
        10'b0010110110: data <= 11'h7f4; 
        10'b0010110111: data <= 11'h7f6; 
        10'b0010111000: data <= 11'h7f5; 
        10'b0010111001: data <= 11'h7fa; 
        10'b0010111010: data <= 11'h7fa; 
        10'b0010111011: data <= 11'h7fd; 
        10'b0010111100: data <= 11'h7fe; 
        10'b0010111101: data <= 11'h000; 
        10'b0010111110: data <= 11'h008; 
        10'b0010111111: data <= 11'h009; 
        10'b0011000000: data <= 11'h003; 
        10'b0011000001: data <= 11'h003; 
        10'b0011000010: data <= 11'h002; 
        10'b0011000011: data <= 11'h000; 
        10'b0011000100: data <= 11'h001; 
        10'b0011000101: data <= 11'h000; 
        10'b0011000110: data <= 11'h001; 
        10'b0011000111: data <= 11'h001; 
        10'b0011001000: data <= 11'h001; 
        10'b0011001001: data <= 11'h002; 
        10'b0011001010: data <= 11'h7ff; 
        10'b0011001011: data <= 11'h000; 
        10'b0011001100: data <= 11'h7ff; 
        10'b0011001101: data <= 11'h7fe; 
        10'b0011001110: data <= 11'h7fa; 
        10'b0011001111: data <= 11'h7f6; 
        10'b0011010000: data <= 11'h7f4; 
        10'b0011010001: data <= 11'h7f7; 
        10'b0011010010: data <= 11'h7f5; 
        10'b0011010011: data <= 11'h7f5; 
        10'b0011010100: data <= 11'h7f5; 
        10'b0011010101: data <= 11'h7f9; 
        10'b0011010110: data <= 11'h7f9; 
        10'b0011010111: data <= 11'h7fb; 
        10'b0011011000: data <= 11'h7fa; 
        10'b0011011001: data <= 11'h7fd; 
        10'b0011011010: data <= 11'h005; 
        10'b0011011011: data <= 11'h007; 
        10'b0011011100: data <= 11'h004; 
        10'b0011011101: data <= 11'h002; 
        10'b0011011110: data <= 11'h002; 
        10'b0011011111: data <= 11'h001; 
        10'b0011100000: data <= 11'h002; 
        10'b0011100001: data <= 11'h002; 
        10'b0011100010: data <= 11'h002; 
        10'b0011100011: data <= 11'h000; 
        10'b0011100100: data <= 11'h001; 
        10'b0011100101: data <= 11'h001; 
        10'b0011100110: data <= 11'h001; 
        10'b0011100111: data <= 11'h000; 
        10'b0011101000: data <= 11'h7fb; 
        10'b0011101001: data <= 11'h7fe; 
        10'b0011101010: data <= 11'h7fd; 
        10'b0011101011: data <= 11'h7fa; 
        10'b0011101100: data <= 11'h7f7; 
        10'b0011101101: data <= 11'h7fa; 
        10'b0011101110: data <= 11'h7f3; 
        10'b0011101111: data <= 11'h7f2; 
        10'b0011110000: data <= 11'h7f5; 
        10'b0011110001: data <= 11'h7f9; 
        10'b0011110010: data <= 11'h7fa; 
        10'b0011110011: data <= 11'h7fe; 
        10'b0011110100: data <= 11'h7fc; 
        10'b0011110101: data <= 11'h7fc; 
        10'b0011110110: data <= 11'h002; 
        10'b0011110111: data <= 11'h004; 
        10'b0011111000: data <= 11'h003; 
        10'b0011111001: data <= 11'h001; 
        10'b0011111010: data <= 11'h001; 
        10'b0011111011: data <= 11'h001; 
        10'b0011111100: data <= 11'h002; 
        10'b0011111101: data <= 11'h002; 
        10'b0011111110: data <= 11'h002; 
        10'b0011111111: data <= 11'h000; 
        10'b0100000000: data <= 11'h7ff; 
        10'b0100000001: data <= 11'h000; 
        10'b0100000010: data <= 11'h7fd; 
        10'b0100000011: data <= 11'h7fe; 
        10'b0100000100: data <= 11'h7ff; 
        10'b0100000101: data <= 11'h000; 
        10'b0100000110: data <= 11'h7fe; 
        10'b0100000111: data <= 11'h7fe; 
        10'b0100001000: data <= 11'h7fe; 
        10'b0100001001: data <= 11'h7fb; 
        10'b0100001010: data <= 11'h7ed; 
        10'b0100001011: data <= 11'h7f2; 
        10'b0100001100: data <= 11'h7fd; 
        10'b0100001101: data <= 11'h7fd; 
        10'b0100001110: data <= 11'h7ff; 
        10'b0100001111: data <= 11'h000; 
        10'b0100010000: data <= 11'h7fe; 
        10'b0100010001: data <= 11'h7fe; 
        10'b0100010010: data <= 11'h001; 
        10'b0100010011: data <= 11'h000; 
        10'b0100010100: data <= 11'h7fe; 
        10'b0100010101: data <= 11'h7fe; 
        10'b0100010110: data <= 11'h7ff; 
        10'b0100010111: data <= 11'h002; 
        10'b0100011000: data <= 11'h001; 
        10'b0100011001: data <= 11'h001; 
        10'b0100011010: data <= 11'h001; 
        10'b0100011011: data <= 11'h000; 
        10'b0100011100: data <= 11'h001; 
        10'b0100011101: data <= 11'h7fd; 
        10'b0100011110: data <= 11'h7fc; 
        10'b0100011111: data <= 11'h7fe; 
        10'b0100100000: data <= 11'h001; 
        10'b0100100001: data <= 11'h005; 
        10'b0100100010: data <= 11'h003; 
        10'b0100100011: data <= 11'h002; 
        10'b0100100100: data <= 11'h003; 
        10'b0100100101: data <= 11'h7f9; 
        10'b0100100110: data <= 11'h7ec; 
        10'b0100100111: data <= 11'h7fa; 
        10'b0100101000: data <= 11'h001; 
        10'b0100101001: data <= 11'h7ff; 
        10'b0100101010: data <= 11'h7ff; 
        10'b0100101011: data <= 11'h001; 
        10'b0100101100: data <= 11'h7fc; 
        10'b0100101101: data <= 11'h7fd; 
        10'b0100101110: data <= 11'h000; 
        10'b0100101111: data <= 11'h7fc; 
        10'b0100110000: data <= 11'h7fe; 
        10'b0100110001: data <= 11'h7fe; 
        10'b0100110010: data <= 11'h001; 
        10'b0100110011: data <= 11'h002; 
        10'b0100110100: data <= 11'h001; 
        10'b0100110101: data <= 11'h001; 
        10'b0100110110: data <= 11'h001; 
        10'b0100110111: data <= 11'h7ff; 
        10'b0100111000: data <= 11'h000; 
        10'b0100111001: data <= 11'h7ff; 
        10'b0100111010: data <= 11'h7fe; 
        10'b0100111011: data <= 11'h001; 
        10'b0100111100: data <= 11'h004; 
        10'b0100111101: data <= 11'h007; 
        10'b0100111110: data <= 11'h00a; 
        10'b0100111111: data <= 11'h006; 
        10'b0101000000: data <= 11'h007; 
        10'b0101000001: data <= 11'h7f5; 
        10'b0101000010: data <= 11'h7f1; 
        10'b0101000011: data <= 11'h002; 
        10'b0101000100: data <= 11'h008; 
        10'b0101000101: data <= 11'h001; 
        10'b0101000110: data <= 11'h000; 
        10'b0101000111: data <= 11'h7ff; 
        10'b0101001000: data <= 11'h7fc; 
        10'b0101001001: data <= 11'h7fc; 
        10'b0101001010: data <= 11'h7fe; 
        10'b0101001011: data <= 11'h7fd; 
        10'b0101001100: data <= 11'h7fc; 
        10'b0101001101: data <= 11'h000; 
        10'b0101001110: data <= 11'h000; 
        10'b0101001111: data <= 11'h001; 
        10'b0101010000: data <= 11'h002; 
        10'b0101010001: data <= 11'h001; 
        10'b0101010010: data <= 11'h001; 
        10'b0101010011: data <= 11'h001; 
        10'b0101010100: data <= 11'h000; 
        10'b0101010101: data <= 11'h7ff; 
        10'b0101010110: data <= 11'h004; 
        10'b0101010111: data <= 11'h007; 
        10'b0101011000: data <= 11'h00a; 
        10'b0101011001: data <= 11'h009; 
        10'b0101011010: data <= 11'h00f; 
        10'b0101011011: data <= 11'h011; 
        10'b0101011100: data <= 11'h010; 
        10'b0101011101: data <= 11'h000; 
        10'b0101011110: data <= 11'h7f8; 
        10'b0101011111: data <= 11'h006; 
        10'b0101100000: data <= 11'h00a; 
        10'b0101100001: data <= 11'h001; 
        10'b0101100010: data <= 11'h000; 
        10'b0101100011: data <= 11'h001; 
        10'b0101100100: data <= 11'h000; 
        10'b0101100101: data <= 11'h000; 
        10'b0101100110: data <= 11'h000; 
        10'b0101100111: data <= 11'h7fe; 
        10'b0101101000: data <= 11'h7fe; 
        10'b0101101001: data <= 11'h7ff; 
        10'b0101101010: data <= 11'h002; 
        10'b0101101011: data <= 11'h001; 
        10'b0101101100: data <= 11'h000; 
        10'b0101101101: data <= 11'h001; 
        10'b0101101110: data <= 11'h000; 
        10'b0101101111: data <= 11'h001; 
        10'b0101110000: data <= 11'h002; 
        10'b0101110001: data <= 11'h005; 
        10'b0101110010: data <= 11'h00a; 
        10'b0101110011: data <= 11'h00b; 
        10'b0101110100: data <= 11'h00d; 
        10'b0101110101: data <= 11'h00b; 
        10'b0101110110: data <= 11'h00d; 
        10'b0101110111: data <= 11'h015; 
        10'b0101111000: data <= 11'h010; 
        10'b0101111001: data <= 11'h000; 
        10'b0101111010: data <= 11'h7fe; 
        10'b0101111011: data <= 11'h007; 
        10'b0101111100: data <= 11'h008; 
        10'b0101111101: data <= 11'h008; 
        10'b0101111110: data <= 11'h006; 
        10'b0101111111: data <= 11'h003; 
        10'b0110000000: data <= 11'h006; 
        10'b0110000001: data <= 11'h004; 
        10'b0110000010: data <= 11'h002; 
        10'b0110000011: data <= 11'h7ff; 
        10'b0110000100: data <= 11'h7ff; 
        10'b0110000101: data <= 11'h000; 
        10'b0110000110: data <= 11'h002; 
        10'b0110000111: data <= 11'h001; 
        10'b0110001000: data <= 11'h000; 
        10'b0110001001: data <= 11'h002; 
        10'b0110001010: data <= 11'h000; 
        10'b0110001011: data <= 11'h002; 
        10'b0110001100: data <= 11'h004; 
        10'b0110001101: data <= 11'h009; 
        10'b0110001110: data <= 11'h00c; 
        10'b0110001111: data <= 11'h00d; 
        10'b0110010000: data <= 11'h00a; 
        10'b0110010001: data <= 11'h009; 
        10'b0110010010: data <= 11'h00b; 
        10'b0110010011: data <= 11'h00e; 
        10'b0110010100: data <= 11'h00a; 
        10'b0110010101: data <= 11'h001; 
        10'b0110010110: data <= 11'h7ff; 
        10'b0110010111: data <= 11'h003; 
        10'b0110011000: data <= 11'h008; 
        10'b0110011001: data <= 11'h00e; 
        10'b0110011010: data <= 11'h009; 
        10'b0110011011: data <= 11'h009; 
        10'b0110011100: data <= 11'h005; 
        10'b0110011101: data <= 11'h003; 
        10'b0110011110: data <= 11'h001; 
        10'b0110011111: data <= 11'h001; 
        10'b0110100000: data <= 11'h000; 
        10'b0110100001: data <= 11'h001; 
        10'b0110100010: data <= 11'h001; 
        10'b0110100011: data <= 11'h001; 
        10'b0110100100: data <= 11'h001; 
        10'b0110100101: data <= 11'h002; 
        10'b0110100110: data <= 11'h001; 
        10'b0110100111: data <= 11'h002; 
        10'b0110101000: data <= 11'h004; 
        10'b0110101001: data <= 11'h004; 
        10'b0110101010: data <= 11'h007; 
        10'b0110101011: data <= 11'h006; 
        10'b0110101100: data <= 11'h00a; 
        10'b0110101101: data <= 11'h009; 
        10'b0110101110: data <= 11'h006; 
        10'b0110101111: data <= 11'h004; 
        10'b0110110000: data <= 11'h005; 
        10'b0110110001: data <= 11'h001; 
        10'b0110110010: data <= 11'h004; 
        10'b0110110011: data <= 11'h006; 
        10'b0110110100: data <= 11'h00c; 
        10'b0110110101: data <= 11'h00b; 
        10'b0110110110: data <= 11'h008; 
        10'b0110110111: data <= 11'h005; 
        10'b0110111000: data <= 11'h7ff; 
        10'b0110111001: data <= 11'h002; 
        10'b0110111010: data <= 11'h003; 
        10'b0110111011: data <= 11'h000; 
        10'b0110111100: data <= 11'h7fe; 
        10'b0110111101: data <= 11'h001; 
        10'b0110111110: data <= 11'h000; 
        10'b0110111111: data <= 11'h001; 
        10'b0111000000: data <= 11'h001; 
        10'b0111000001: data <= 11'h000; 
        10'b0111000010: data <= 11'h000; 
        10'b0111000011: data <= 11'h000; 
        10'b0111000100: data <= 11'h001; 
        10'b0111000101: data <= 11'h003; 
        10'b0111000110: data <= 11'h004; 
        10'b0111000111: data <= 11'h007; 
        10'b0111001000: data <= 11'h00b; 
        10'b0111001001: data <= 11'h008; 
        10'b0111001010: data <= 11'h002; 
        10'b0111001011: data <= 11'h000; 
        10'b0111001100: data <= 11'h002; 
        10'b0111001101: data <= 11'h003; 
        10'b0111001110: data <= 11'h00a; 
        10'b0111001111: data <= 11'h00e; 
        10'b0111010000: data <= 11'h00e; 
        10'b0111010001: data <= 11'h00c; 
        10'b0111010010: data <= 11'h008; 
        10'b0111010011: data <= 11'h001; 
        10'b0111010100: data <= 11'h003; 
        10'b0111010101: data <= 11'h005; 
        10'b0111010110: data <= 11'h001; 
        10'b0111010111: data <= 11'h7ff; 
        10'b0111011000: data <= 11'h000; 
        10'b0111011001: data <= 11'h000; 
        10'b0111011010: data <= 11'h001; 
        10'b0111011011: data <= 11'h001; 
        10'b0111011100: data <= 11'h001; 
        10'b0111011101: data <= 11'h001; 
        10'b0111011110: data <= 11'h002; 
        10'b0111011111: data <= 11'h000; 
        10'b0111100000: data <= 11'h7ff; 
        10'b0111100001: data <= 11'h7fe; 
        10'b0111100010: data <= 11'h001; 
        10'b0111100011: data <= 11'h006; 
        10'b0111100100: data <= 11'h00b; 
        10'b0111100101: data <= 11'h00a; 
        10'b0111100110: data <= 11'h004; 
        10'b0111100111: data <= 11'h003; 
        10'b0111101000: data <= 11'h004; 
        10'b0111101001: data <= 11'h00a; 
        10'b0111101010: data <= 11'h010; 
        10'b0111101011: data <= 11'h00d; 
        10'b0111101100: data <= 11'h00b; 
        10'b0111101101: data <= 11'h003; 
        10'b0111101110: data <= 11'h001; 
        10'b0111101111: data <= 11'h7fc; 
        10'b0111110000: data <= 11'h001; 
        10'b0111110001: data <= 11'h000; 
        10'b0111110010: data <= 11'h7fe; 
        10'b0111110011: data <= 11'h7ff; 
        10'b0111110100: data <= 11'h7ff; 
        10'b0111110101: data <= 11'h7ff; 
        10'b0111110110: data <= 11'h001; 
        10'b0111110111: data <= 11'h002; 
        10'b0111111000: data <= 11'h001; 
        10'b0111111001: data <= 11'h001; 
        10'b0111111010: data <= 11'h001; 
        10'b0111111011: data <= 11'h000; 
        10'b0111111100: data <= 11'h7ff; 
        10'b0111111101: data <= 11'h7fd; 
        10'b0111111110: data <= 11'h7fd; 
        10'b0111111111: data <= 11'h000; 
        10'b1000000000: data <= 11'h003; 
        10'b1000000001: data <= 11'h001; 
        10'b1000000010: data <= 11'h7fe; 
        10'b1000000011: data <= 11'h7ff; 
        10'b1000000100: data <= 11'h004; 
        10'b1000000101: data <= 11'h004; 
        10'b1000000110: data <= 11'h007; 
        10'b1000000111: data <= 11'h006; 
        10'b1000001000: data <= 11'h003; 
        10'b1000001001: data <= 11'h7fb; 
        10'b1000001010: data <= 11'h7fb; 
        10'b1000001011: data <= 11'h7f9; 
        10'b1000001100: data <= 11'h7fc; 
        10'b1000001101: data <= 11'h7fc; 
        10'b1000001110: data <= 11'h7fa; 
        10'b1000001111: data <= 11'h7fc; 
        10'b1000010000: data <= 11'h7ff; 
        10'b1000010001: data <= 11'h7ff; 
        10'b1000010010: data <= 11'h001; 
        10'b1000010011: data <= 11'h000; 
        10'b1000010100: data <= 11'h001; 
        10'b1000010101: data <= 11'h002; 
        10'b1000010110: data <= 11'h001; 
        10'b1000010111: data <= 11'h000; 
        10'b1000011000: data <= 11'h7fd; 
        10'b1000011001: data <= 11'h7fc; 
        10'b1000011010: data <= 11'h7fb; 
        10'b1000011011: data <= 11'h7f8; 
        10'b1000011100: data <= 11'h7f7; 
        10'b1000011101: data <= 11'h7f7; 
        10'b1000011110: data <= 11'h7f5; 
        10'b1000011111: data <= 11'h7f6; 
        10'b1000100000: data <= 11'h7f7; 
        10'b1000100001: data <= 11'h7fb; 
        10'b1000100010: data <= 11'h7fe; 
        10'b1000100011: data <= 11'h001; 
        10'b1000100100: data <= 11'h7fc; 
        10'b1000100101: data <= 11'h7fc; 
        10'b1000100110: data <= 11'h7fc; 
        10'b1000100111: data <= 11'h7fa; 
        10'b1000101000: data <= 11'h7f9; 
        10'b1000101001: data <= 11'h7fa; 
        10'b1000101010: data <= 11'h7fa; 
        10'b1000101011: data <= 11'h7fc; 
        10'b1000101100: data <= 11'h7ff; 
        10'b1000101101: data <= 11'h001; 
        10'b1000101110: data <= 11'h002; 
        10'b1000101111: data <= 11'h001; 
        10'b1000110000: data <= 11'h002; 
        10'b1000110001: data <= 11'h002; 
        10'b1000110010: data <= 11'h001; 
        10'b1000110011: data <= 11'h000; 
        10'b1000110100: data <= 11'h7fd; 
        10'b1000110101: data <= 11'h7fc; 
        10'b1000110110: data <= 11'h7fa; 
        10'b1000110111: data <= 11'h7f6; 
        10'b1000111000: data <= 11'h7f4; 
        10'b1000111001: data <= 11'h7f3; 
        10'b1000111010: data <= 11'h7f3; 
        10'b1000111011: data <= 11'h7f6; 
        10'b1000111100: data <= 11'h7f8; 
        10'b1000111101: data <= 11'h7f7; 
        10'b1000111110: data <= 11'h7fb; 
        10'b1000111111: data <= 11'h7fd; 
        10'b1001000000: data <= 11'h7ff; 
        10'b1001000001: data <= 11'h7ff; 
        10'b1001000010: data <= 11'h7fe; 
        10'b1001000011: data <= 11'h7fb; 
        10'b1001000100: data <= 11'h7fd; 
        10'b1001000101: data <= 11'h7fc; 
        10'b1001000110: data <= 11'h7fc; 
        10'b1001000111: data <= 11'h7fe; 
        10'b1001001000: data <= 11'h7fe; 
        10'b1001001001: data <= 11'h000; 
        10'b1001001010: data <= 11'h001; 
        10'b1001001011: data <= 11'h002; 
        10'b1001001100: data <= 11'h000; 
        10'b1001001101: data <= 11'h001; 
        10'b1001001110: data <= 11'h000; 
        10'b1001001111: data <= 11'h000; 
        10'b1001010000: data <= 11'h000; 
        10'b1001010001: data <= 11'h7fe; 
        10'b1001010010: data <= 11'h7fa; 
        10'b1001010011: data <= 11'h7f7; 
        10'b1001010100: data <= 11'h7f8; 
        10'b1001010101: data <= 11'h7f7; 
        10'b1001010110: data <= 11'h7f8; 
        10'b1001010111: data <= 11'h7fa; 
        10'b1001011000: data <= 11'h7fb; 
        10'b1001011001: data <= 11'h7fc; 
        10'b1001011010: data <= 11'h7fb; 
        10'b1001011011: data <= 11'h7fe; 
        10'b1001011100: data <= 11'h7fd; 
        10'b1001011101: data <= 11'h001; 
        10'b1001011110: data <= 11'h7ff; 
        10'b1001011111: data <= 11'h000; 
        10'b1001100000: data <= 11'h000; 
        10'b1001100001: data <= 11'h7fd; 
        10'b1001100010: data <= 11'h7fd; 
        10'b1001100011: data <= 11'h000; 
        10'b1001100100: data <= 11'h000; 
        10'b1001100101: data <= 11'h001; 
        10'b1001100110: data <= 11'h001; 
        10'b1001100111: data <= 11'h001; 
        10'b1001101000: data <= 11'h001; 
        10'b1001101001: data <= 11'h001; 
        10'b1001101010: data <= 11'h001; 
        10'b1001101011: data <= 11'h001; 
        10'b1001101100: data <= 11'h000; 
        10'b1001101101: data <= 11'h7ff; 
        10'b1001101110: data <= 11'h7fd; 
        10'b1001101111: data <= 11'h7fc; 
        10'b1001110000: data <= 11'h7fa; 
        10'b1001110001: data <= 11'h7fd; 
        10'b1001110010: data <= 11'h7fc; 
        10'b1001110011: data <= 11'h7fe; 
        10'b1001110100: data <= 11'h7fd; 
        10'b1001110101: data <= 11'h7fe; 
        10'b1001110110: data <= 11'h7fd; 
        10'b1001110111: data <= 11'h7fe; 
        10'b1001111000: data <= 11'h7fe; 
        10'b1001111001: data <= 11'h001; 
        10'b1001111010: data <= 11'h003; 
        10'b1001111011: data <= 11'h004; 
        10'b1001111100: data <= 11'h003; 
        10'b1001111101: data <= 11'h002; 
        10'b1001111110: data <= 11'h7ff; 
        10'b1001111111: data <= 11'h7ff; 
        10'b1010000000: data <= 11'h000; 
        10'b1010000001: data <= 11'h001; 
        10'b1010000010: data <= 11'h000; 
        10'b1010000011: data <= 11'h001; 
        10'b1010000100: data <= 11'h001; 
        10'b1010000101: data <= 11'h000; 
        10'b1010000110: data <= 11'h001; 
        10'b1010000111: data <= 11'h001; 
        10'b1010001000: data <= 11'h001; 
        10'b1010001001: data <= 11'h001; 
        10'b1010001010: data <= 11'h7ff; 
        10'b1010001011: data <= 11'h7fe; 
        10'b1010001100: data <= 11'h7fe; 
        10'b1010001101: data <= 11'h001; 
        10'b1010001110: data <= 11'h7fe; 
        10'b1010001111: data <= 11'h000; 
        10'b1010010000: data <= 11'h7fe; 
        10'b1010010001: data <= 11'h7fe; 
        10'b1010010010: data <= 11'h7fe; 
        10'b1010010011: data <= 11'h000; 
        10'b1010010100: data <= 11'h001; 
        10'b1010010101: data <= 11'h002; 
        10'b1010010110: data <= 11'h005; 
        10'b1010010111: data <= 11'h005; 
        10'b1010011000: data <= 11'h004; 
        10'b1010011001: data <= 11'h002; 
        10'b1010011010: data <= 11'h7ff; 
        10'b1010011011: data <= 11'h001; 
        10'b1010011100: data <= 11'h001; 
        10'b1010011101: data <= 11'h001; 
        10'b1010011110: data <= 11'h000; 
        10'b1010011111: data <= 11'h002; 
        10'b1010100000: data <= 11'h001; 
        10'b1010100001: data <= 11'h002; 
        10'b1010100010: data <= 11'h001; 
        10'b1010100011: data <= 11'h002; 
        10'b1010100100: data <= 11'h000; 
        10'b1010100101: data <= 11'h001; 
        10'b1010100110: data <= 11'h000; 
        10'b1010100111: data <= 11'h7fe; 
        10'b1010101000: data <= 11'h7fe; 
        10'b1010101001: data <= 11'h7ff; 
        10'b1010101010: data <= 11'h7fe; 
        10'b1010101011: data <= 11'h000; 
        10'b1010101100: data <= 11'h7fe; 
        10'b1010101101: data <= 11'h7fe; 
        10'b1010101110: data <= 11'h7fd; 
        10'b1010101111: data <= 11'h7fd; 
        10'b1010110000: data <= 11'h7ff; 
        10'b1010110001: data <= 11'h7ff; 
        10'b1010110010: data <= 11'h000; 
        10'b1010110011: data <= 11'h002; 
        10'b1010110100: data <= 11'h002; 
        10'b1010110101: data <= 11'h7ff; 
        10'b1010110110: data <= 11'h000; 
        10'b1010110111: data <= 11'h001; 
        10'b1010111000: data <= 11'h002; 
        10'b1010111001: data <= 11'h000; 
        10'b1010111010: data <= 11'h000; 
        10'b1010111011: data <= 11'h001; 
        10'b1010111100: data <= 11'h002; 
        10'b1010111101: data <= 11'h002; 
        10'b1010111110: data <= 11'h002; 
        10'b1010111111: data <= 11'h000; 
        10'b1011000000: data <= 11'h002; 
        10'b1011000001: data <= 11'h000; 
        10'b1011000010: data <= 11'h7ff; 
        10'b1011000011: data <= 11'h7fe; 
        10'b1011000100: data <= 11'h7fd; 
        10'b1011000101: data <= 11'h7fd; 
        10'b1011000110: data <= 11'h7fb; 
        10'b1011000111: data <= 11'h7fa; 
        10'b1011001000: data <= 11'h7fa; 
        10'b1011001001: data <= 11'h7fa; 
        10'b1011001010: data <= 11'h7fb; 
        10'b1011001011: data <= 11'h7fb; 
        10'b1011001100: data <= 11'h7f9; 
        10'b1011001101: data <= 11'h7f8; 
        10'b1011001110: data <= 11'h7f9; 
        10'b1011001111: data <= 11'h7fc; 
        10'b1011010000: data <= 11'h7fd; 
        10'b1011010001: data <= 11'h7ff; 
        10'b1011010010: data <= 11'h000; 
        10'b1011010011: data <= 11'h001; 
        10'b1011010100: data <= 11'h000; 
        10'b1011010101: data <= 11'h002; 
        10'b1011010110: data <= 11'h001; 
        10'b1011010111: data <= 11'h001; 
        10'b1011011000: data <= 11'h001; 
        10'b1011011001: data <= 11'h001; 
        10'b1011011010: data <= 11'h000; 
        10'b1011011011: data <= 11'h001; 
        10'b1011011100: data <= 11'h000; 
        10'b1011011101: data <= 11'h000; 
        10'b1011011110: data <= 11'h001; 
        10'b1011011111: data <= 11'h000; 
        10'b1011100000: data <= 11'h000; 
        10'b1011100001: data <= 11'h7fe; 
        10'b1011100010: data <= 11'h7fb; 
        10'b1011100011: data <= 11'h7fc; 
        10'b1011100100: data <= 11'h7fb; 
        10'b1011100101: data <= 11'h7fa; 
        10'b1011100110: data <= 11'h7f9; 
        10'b1011100111: data <= 11'h7fb; 
        10'b1011101000: data <= 11'h7fa; 
        10'b1011101001: data <= 11'h7fb; 
        10'b1011101010: data <= 11'h7fc; 
        10'b1011101011: data <= 11'h7fe; 
        10'b1011101100: data <= 11'h7ff; 
        10'b1011101101: data <= 11'h001; 
        10'b1011101110: data <= 11'h001; 
        10'b1011101111: data <= 11'h000; 
        10'b1011110000: data <= 11'h001; 
        10'b1011110001: data <= 11'h000; 
        10'b1011110010: data <= 11'h002; 
        10'b1011110011: data <= 11'h001; 
        10'b1011110100: data <= 11'h001; 
        10'b1011110101: data <= 11'h000; 
        10'b1011110110: data <= 11'h000; 
        10'b1011110111: data <= 11'h002; 
        10'b1011111000: data <= 11'h001; 
        10'b1011111001: data <= 11'h002; 
        10'b1011111010: data <= 11'h001; 
        10'b1011111011: data <= 11'h002; 
        10'b1011111100: data <= 11'h000; 
        10'b1011111101: data <= 11'h001; 
        10'b1011111110: data <= 11'h000; 
        10'b1011111111: data <= 11'h000; 
        10'b1100000000: data <= 11'h000; 
        10'b1100000001: data <= 11'h000; 
        10'b1100000010: data <= 11'h7ff; 
        10'b1100000011: data <= 11'h002; 
        10'b1100000100: data <= 11'h000; 
        10'b1100000101: data <= 11'h000; 
        10'b1100000110: data <= 11'h000; 
        10'b1100000111: data <= 11'h001; 
        10'b1100001000: data <= 11'h001; 
        10'b1100001001: data <= 11'h001; 
        10'b1100001010: data <= 11'h001; 
        10'b1100001011: data <= 11'h001; 
        10'b1100001100: data <= 11'h001; 
        10'b1100001101: data <= 11'h002; 
        10'b1100001110: data <= 11'h001; 
        10'b1100001111: data <= 11'h001; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 6) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 12'h000; 
        10'b0000000001: data <= 12'h001; 
        10'b0000000010: data <= 12'h004; 
        10'b0000000011: data <= 12'h004; 
        10'b0000000100: data <= 12'h000; 
        10'b0000000101: data <= 12'h000; 
        10'b0000000110: data <= 12'h003; 
        10'b0000000111: data <= 12'h001; 
        10'b0000001000: data <= 12'h000; 
        10'b0000001001: data <= 12'h001; 
        10'b0000001010: data <= 12'h000; 
        10'b0000001011: data <= 12'h003; 
        10'b0000001100: data <= 12'h004; 
        10'b0000001101: data <= 12'h002; 
        10'b0000001110: data <= 12'h003; 
        10'b0000001111: data <= 12'h000; 
        10'b0000010000: data <= 12'h002; 
        10'b0000010001: data <= 12'h003; 
        10'b0000010010: data <= 12'h001; 
        10'b0000010011: data <= 12'h003; 
        10'b0000010100: data <= 12'h000; 
        10'b0000010101: data <= 12'h002; 
        10'b0000010110: data <= 12'h004; 
        10'b0000010111: data <= 12'h000; 
        10'b0000011000: data <= 12'h004; 
        10'b0000011001: data <= 12'h001; 
        10'b0000011010: data <= 12'h004; 
        10'b0000011011: data <= 12'h002; 
        10'b0000011100: data <= 12'h001; 
        10'b0000011101: data <= 12'h002; 
        10'b0000011110: data <= 12'h000; 
        10'b0000011111: data <= 12'h000; 
        10'b0000100000: data <= 12'h002; 
        10'b0000100001: data <= 12'h004; 
        10'b0000100010: data <= 12'h001; 
        10'b0000100011: data <= 12'hfff; 
        10'b0000100100: data <= 12'h002; 
        10'b0000100101: data <= 12'h000; 
        10'b0000100110: data <= 12'h002; 
        10'b0000100111: data <= 12'hfff; 
        10'b0000101000: data <= 12'h001; 
        10'b0000101001: data <= 12'hffe; 
        10'b0000101010: data <= 12'h000; 
        10'b0000101011: data <= 12'h002; 
        10'b0000101100: data <= 12'h003; 
        10'b0000101101: data <= 12'h001; 
        10'b0000101110: data <= 12'h000; 
        10'b0000101111: data <= 12'h001; 
        10'b0000110000: data <= 12'h003; 
        10'b0000110001: data <= 12'h000; 
        10'b0000110010: data <= 12'h000; 
        10'b0000110011: data <= 12'h000; 
        10'b0000110100: data <= 12'h003; 
        10'b0000110101: data <= 12'h003; 
        10'b0000110110: data <= 12'h001; 
        10'b0000110111: data <= 12'h003; 
        10'b0000111000: data <= 12'h003; 
        10'b0000111001: data <= 12'h002; 
        10'b0000111010: data <= 12'h003; 
        10'b0000111011: data <= 12'h003; 
        10'b0000111100: data <= 12'h003; 
        10'b0000111101: data <= 12'h003; 
        10'b0000111110: data <= 12'h004; 
        10'b0000111111: data <= 12'hfff; 
        10'b0001000000: data <= 12'hfff; 
        10'b0001000001: data <= 12'h001; 
        10'b0001000010: data <= 12'h000; 
        10'b0001000011: data <= 12'hffe; 
        10'b0001000100: data <= 12'hff7; 
        10'b0001000101: data <= 12'hffd; 
        10'b0001000110: data <= 12'hffc; 
        10'b0001000111: data <= 12'hffa; 
        10'b0001001000: data <= 12'hffc; 
        10'b0001001001: data <= 12'hfff; 
        10'b0001001010: data <= 12'h001; 
        10'b0001001011: data <= 12'h003; 
        10'b0001001100: data <= 12'h004; 
        10'b0001001101: data <= 12'h002; 
        10'b0001001110: data <= 12'h004; 
        10'b0001001111: data <= 12'h001; 
        10'b0001010000: data <= 12'h001; 
        10'b0001010001: data <= 12'h002; 
        10'b0001010010: data <= 12'h000; 
        10'b0001010011: data <= 12'h002; 
        10'b0001010100: data <= 12'h003; 
        10'b0001010101: data <= 12'h003; 
        10'b0001010110: data <= 12'h001; 
        10'b0001010111: data <= 12'h002; 
        10'b0001011000: data <= 12'h002; 
        10'b0001011001: data <= 12'h000; 
        10'b0001011010: data <= 12'h002; 
        10'b0001011011: data <= 12'hffe; 
        10'b0001011100: data <= 12'hffd; 
        10'b0001011101: data <= 12'hffe; 
        10'b0001011110: data <= 12'hff9; 
        10'b0001011111: data <= 12'hff7; 
        10'b0001100000: data <= 12'hff2; 
        10'b0001100001: data <= 12'hff3; 
        10'b0001100010: data <= 12'hff3; 
        10'b0001100011: data <= 12'hff1; 
        10'b0001100100: data <= 12'hff6; 
        10'b0001100101: data <= 12'hffb; 
        10'b0001100110: data <= 12'h001; 
        10'b0001100111: data <= 12'h002; 
        10'b0001101000: data <= 12'h003; 
        10'b0001101001: data <= 12'h004; 
        10'b0001101010: data <= 12'h001; 
        10'b0001101011: data <= 12'h001; 
        10'b0001101100: data <= 12'h004; 
        10'b0001101101: data <= 12'h004; 
        10'b0001101110: data <= 12'h001; 
        10'b0001101111: data <= 12'h002; 
        10'b0001110000: data <= 12'h004; 
        10'b0001110001: data <= 12'h003; 
        10'b0001110010: data <= 12'h003; 
        10'b0001110011: data <= 12'h003; 
        10'b0001110100: data <= 12'h002; 
        10'b0001110101: data <= 12'h003; 
        10'b0001110110: data <= 12'hffd; 
        10'b0001110111: data <= 12'hfff; 
        10'b0001111000: data <= 12'hffb; 
        10'b0001111001: data <= 12'hffc; 
        10'b0001111010: data <= 12'hff4; 
        10'b0001111011: data <= 12'hff4; 
        10'b0001111100: data <= 12'hff0; 
        10'b0001111101: data <= 12'hff3; 
        10'b0001111110: data <= 12'hff0; 
        10'b0001111111: data <= 12'hff2; 
        10'b0010000000: data <= 12'hff9; 
        10'b0010000001: data <= 12'hffa; 
        10'b0010000010: data <= 12'hffc; 
        10'b0010000011: data <= 12'h004; 
        10'b0010000100: data <= 12'h005; 
        10'b0010000101: data <= 12'h006; 
        10'b0010000110: data <= 12'h005; 
        10'b0010000111: data <= 12'h007; 
        10'b0010001000: data <= 12'h002; 
        10'b0010001001: data <= 12'h004; 
        10'b0010001010: data <= 12'h001; 
        10'b0010001011: data <= 12'h001; 
        10'b0010001100: data <= 12'h004; 
        10'b0010001101: data <= 12'h001; 
        10'b0010001110: data <= 12'h003; 
        10'b0010001111: data <= 12'h001; 
        10'b0010010000: data <= 12'h003; 
        10'b0010010001: data <= 12'h001; 
        10'b0010010010: data <= 12'h002; 
        10'b0010010011: data <= 12'hffe; 
        10'b0010010100: data <= 12'h001; 
        10'b0010010101: data <= 12'hffd; 
        10'b0010010110: data <= 12'hff7; 
        10'b0010010111: data <= 12'hffa; 
        10'b0010011000: data <= 12'hff6; 
        10'b0010011001: data <= 12'hff3; 
        10'b0010011010: data <= 12'hff7; 
        10'b0010011011: data <= 12'hff9; 
        10'b0010011100: data <= 12'hfff; 
        10'b0010011101: data <= 12'h001; 
        10'b0010011110: data <= 12'hffe; 
        10'b0010011111: data <= 12'h003; 
        10'b0010100000: data <= 12'h004; 
        10'b0010100001: data <= 12'h005; 
        10'b0010100010: data <= 12'h00c; 
        10'b0010100011: data <= 12'h00d; 
        10'b0010100100: data <= 12'h007; 
        10'b0010100101: data <= 12'hfff; 
        10'b0010100110: data <= 12'h001; 
        10'b0010100111: data <= 12'h001; 
        10'b0010101000: data <= 12'h004; 
        10'b0010101001: data <= 12'h004; 
        10'b0010101010: data <= 12'h001; 
        10'b0010101011: data <= 12'h003; 
        10'b0010101100: data <= 12'h004; 
        10'b0010101101: data <= 12'h003; 
        10'b0010101110: data <= 12'h003; 
        10'b0010101111: data <= 12'h000; 
        10'b0010110000: data <= 12'hfff; 
        10'b0010110001: data <= 12'hffc; 
        10'b0010110010: data <= 12'hff9; 
        10'b0010110011: data <= 12'hff3; 
        10'b0010110100: data <= 12'hfed; 
        10'b0010110101: data <= 12'hfe9; 
        10'b0010110110: data <= 12'hfe8; 
        10'b0010110111: data <= 12'hfeb; 
        10'b0010111000: data <= 12'hfeb; 
        10'b0010111001: data <= 12'hff4; 
        10'b0010111010: data <= 12'hff3; 
        10'b0010111011: data <= 12'hffa; 
        10'b0010111100: data <= 12'hffc; 
        10'b0010111101: data <= 12'h000; 
        10'b0010111110: data <= 12'h011; 
        10'b0010111111: data <= 12'h011; 
        10'b0011000000: data <= 12'h007; 
        10'b0011000001: data <= 12'h005; 
        10'b0011000010: data <= 12'h004; 
        10'b0011000011: data <= 12'h000; 
        10'b0011000100: data <= 12'h002; 
        10'b0011000101: data <= 12'h001; 
        10'b0011000110: data <= 12'h001; 
        10'b0011000111: data <= 12'h002; 
        10'b0011001000: data <= 12'h001; 
        10'b0011001001: data <= 12'h003; 
        10'b0011001010: data <= 12'hffe; 
        10'b0011001011: data <= 12'h000; 
        10'b0011001100: data <= 12'hffe; 
        10'b0011001101: data <= 12'hffb; 
        10'b0011001110: data <= 12'hff4; 
        10'b0011001111: data <= 12'hfed; 
        10'b0011010000: data <= 12'hfe7; 
        10'b0011010001: data <= 12'hfee; 
        10'b0011010010: data <= 12'hfea; 
        10'b0011010011: data <= 12'hfea; 
        10'b0011010100: data <= 12'hfe9; 
        10'b0011010101: data <= 12'hff1; 
        10'b0011010110: data <= 12'hff1; 
        10'b0011010111: data <= 12'hff6; 
        10'b0011011000: data <= 12'hff4; 
        10'b0011011001: data <= 12'hffb; 
        10'b0011011010: data <= 12'h00a; 
        10'b0011011011: data <= 12'h00e; 
        10'b0011011100: data <= 12'h007; 
        10'b0011011101: data <= 12'h004; 
        10'b0011011110: data <= 12'h004; 
        10'b0011011111: data <= 12'h002; 
        10'b0011100000: data <= 12'h004; 
        10'b0011100001: data <= 12'h003; 
        10'b0011100010: data <= 12'h004; 
        10'b0011100011: data <= 12'h001; 
        10'b0011100100: data <= 12'h001; 
        10'b0011100101: data <= 12'h002; 
        10'b0011100110: data <= 12'h001; 
        10'b0011100111: data <= 12'hfff; 
        10'b0011101000: data <= 12'hff7; 
        10'b0011101001: data <= 12'hffb; 
        10'b0011101010: data <= 12'hffa; 
        10'b0011101011: data <= 12'hff4; 
        10'b0011101100: data <= 12'hfee; 
        10'b0011101101: data <= 12'hff4; 
        10'b0011101110: data <= 12'hfe6; 
        10'b0011101111: data <= 12'hfe5; 
        10'b0011110000: data <= 12'hfeb; 
        10'b0011110001: data <= 12'hff3; 
        10'b0011110010: data <= 12'hff4; 
        10'b0011110011: data <= 12'hffc; 
        10'b0011110100: data <= 12'hff9; 
        10'b0011110101: data <= 12'hff9; 
        10'b0011110110: data <= 12'h005; 
        10'b0011110111: data <= 12'h007; 
        10'b0011111000: data <= 12'h006; 
        10'b0011111001: data <= 12'h001; 
        10'b0011111010: data <= 12'h001; 
        10'b0011111011: data <= 12'h003; 
        10'b0011111100: data <= 12'h004; 
        10'b0011111101: data <= 12'h004; 
        10'b0011111110: data <= 12'h003; 
        10'b0011111111: data <= 12'h001; 
        10'b0100000000: data <= 12'hffe; 
        10'b0100000001: data <= 12'h000; 
        10'b0100000010: data <= 12'hffa; 
        10'b0100000011: data <= 12'hffc; 
        10'b0100000100: data <= 12'hffd; 
        10'b0100000101: data <= 12'hfff; 
        10'b0100000110: data <= 12'hffd; 
        10'b0100000111: data <= 12'hffc; 
        10'b0100001000: data <= 12'hffc; 
        10'b0100001001: data <= 12'hff6; 
        10'b0100001010: data <= 12'hfda; 
        10'b0100001011: data <= 12'hfe4; 
        10'b0100001100: data <= 12'hff9; 
        10'b0100001101: data <= 12'hffb; 
        10'b0100001110: data <= 12'hffe; 
        10'b0100001111: data <= 12'h001; 
        10'b0100010000: data <= 12'hffc; 
        10'b0100010001: data <= 12'hffc; 
        10'b0100010010: data <= 12'h002; 
        10'b0100010011: data <= 12'h000; 
        10'b0100010100: data <= 12'hffb; 
        10'b0100010101: data <= 12'hffb; 
        10'b0100010110: data <= 12'hffe; 
        10'b0100010111: data <= 12'h003; 
        10'b0100011000: data <= 12'h002; 
        10'b0100011001: data <= 12'h002; 
        10'b0100011010: data <= 12'h002; 
        10'b0100011011: data <= 12'h000; 
        10'b0100011100: data <= 12'h002; 
        10'b0100011101: data <= 12'hffb; 
        10'b0100011110: data <= 12'hff8; 
        10'b0100011111: data <= 12'hffc; 
        10'b0100100000: data <= 12'h001; 
        10'b0100100001: data <= 12'h00b; 
        10'b0100100010: data <= 12'h007; 
        10'b0100100011: data <= 12'h005; 
        10'b0100100100: data <= 12'h006; 
        10'b0100100101: data <= 12'hff1; 
        10'b0100100110: data <= 12'hfd8; 
        10'b0100100111: data <= 12'hff4; 
        10'b0100101000: data <= 12'h001; 
        10'b0100101001: data <= 12'hffe; 
        10'b0100101010: data <= 12'hfff; 
        10'b0100101011: data <= 12'h001; 
        10'b0100101100: data <= 12'hff8; 
        10'b0100101101: data <= 12'hffb; 
        10'b0100101110: data <= 12'hfff; 
        10'b0100101111: data <= 12'hff7; 
        10'b0100110000: data <= 12'hffb; 
        10'b0100110001: data <= 12'hffd; 
        10'b0100110010: data <= 12'h002; 
        10'b0100110011: data <= 12'h004; 
        10'b0100110100: data <= 12'h003; 
        10'b0100110101: data <= 12'h003; 
        10'b0100110110: data <= 12'h002; 
        10'b0100110111: data <= 12'hffe; 
        10'b0100111000: data <= 12'hfff; 
        10'b0100111001: data <= 12'hffd; 
        10'b0100111010: data <= 12'hffd; 
        10'b0100111011: data <= 12'h003; 
        10'b0100111100: data <= 12'h008; 
        10'b0100111101: data <= 12'h00e; 
        10'b0100111110: data <= 12'h013; 
        10'b0100111111: data <= 12'h00c; 
        10'b0101000000: data <= 12'h00e; 
        10'b0101000001: data <= 12'hfea; 
        10'b0101000010: data <= 12'hfe2; 
        10'b0101000011: data <= 12'h004; 
        10'b0101000100: data <= 12'h010; 
        10'b0101000101: data <= 12'h003; 
        10'b0101000110: data <= 12'hfff; 
        10'b0101000111: data <= 12'hffd; 
        10'b0101001000: data <= 12'hff7; 
        10'b0101001001: data <= 12'hff9; 
        10'b0101001010: data <= 12'hffc; 
        10'b0101001011: data <= 12'hff9; 
        10'b0101001100: data <= 12'hff8; 
        10'b0101001101: data <= 12'h000; 
        10'b0101001110: data <= 12'h000; 
        10'b0101001111: data <= 12'h001; 
        10'b0101010000: data <= 12'h003; 
        10'b0101010001: data <= 12'h003; 
        10'b0101010010: data <= 12'h001; 
        10'b0101010011: data <= 12'h002; 
        10'b0101010100: data <= 12'h000; 
        10'b0101010101: data <= 12'hffd; 
        10'b0101010110: data <= 12'h008; 
        10'b0101010111: data <= 12'h00d; 
        10'b0101011000: data <= 12'h014; 
        10'b0101011001: data <= 12'h012; 
        10'b0101011010: data <= 12'h01e; 
        10'b0101011011: data <= 12'h022; 
        10'b0101011100: data <= 12'h020; 
        10'b0101011101: data <= 12'hfff; 
        10'b0101011110: data <= 12'hff0; 
        10'b0101011111: data <= 12'h00d; 
        10'b0101100000: data <= 12'h014; 
        10'b0101100001: data <= 12'h002; 
        10'b0101100010: data <= 12'h001; 
        10'b0101100011: data <= 12'h003; 
        10'b0101100100: data <= 12'h000; 
        10'b0101100101: data <= 12'h001; 
        10'b0101100110: data <= 12'hfff; 
        10'b0101100111: data <= 12'hffc; 
        10'b0101101000: data <= 12'hffc; 
        10'b0101101001: data <= 12'hfff; 
        10'b0101101010: data <= 12'h004; 
        10'b0101101011: data <= 12'h003; 
        10'b0101101100: data <= 12'h000; 
        10'b0101101101: data <= 12'h003; 
        10'b0101101110: data <= 12'h000; 
        10'b0101101111: data <= 12'h001; 
        10'b0101110000: data <= 12'h003; 
        10'b0101110001: data <= 12'h00a; 
        10'b0101110010: data <= 12'h014; 
        10'b0101110011: data <= 12'h017; 
        10'b0101110100: data <= 12'h01a; 
        10'b0101110101: data <= 12'h016; 
        10'b0101110110: data <= 12'h01a; 
        10'b0101110111: data <= 12'h02a; 
        10'b0101111000: data <= 12'h020; 
        10'b0101111001: data <= 12'h000; 
        10'b0101111010: data <= 12'hffc; 
        10'b0101111011: data <= 12'h00f; 
        10'b0101111100: data <= 12'h00f; 
        10'b0101111101: data <= 12'h011; 
        10'b0101111110: data <= 12'h00c; 
        10'b0101111111: data <= 12'h005; 
        10'b0110000000: data <= 12'h00c; 
        10'b0110000001: data <= 12'h009; 
        10'b0110000010: data <= 12'h004; 
        10'b0110000011: data <= 12'hffe; 
        10'b0110000100: data <= 12'hffe; 
        10'b0110000101: data <= 12'h000; 
        10'b0110000110: data <= 12'h004; 
        10'b0110000111: data <= 12'h003; 
        10'b0110001000: data <= 12'h000; 
        10'b0110001001: data <= 12'h004; 
        10'b0110001010: data <= 12'h000; 
        10'b0110001011: data <= 12'h004; 
        10'b0110001100: data <= 12'h009; 
        10'b0110001101: data <= 12'h011; 
        10'b0110001110: data <= 12'h018; 
        10'b0110001111: data <= 12'h01a; 
        10'b0110010000: data <= 12'h014; 
        10'b0110010001: data <= 12'h013; 
        10'b0110010010: data <= 12'h017; 
        10'b0110010011: data <= 12'h01b; 
        10'b0110010100: data <= 12'h014; 
        10'b0110010101: data <= 12'h002; 
        10'b0110010110: data <= 12'hffd; 
        10'b0110010111: data <= 12'h005; 
        10'b0110011000: data <= 12'h011; 
        10'b0110011001: data <= 12'h01c; 
        10'b0110011010: data <= 12'h013; 
        10'b0110011011: data <= 12'h011; 
        10'b0110011100: data <= 12'h00a; 
        10'b0110011101: data <= 12'h006; 
        10'b0110011110: data <= 12'h002; 
        10'b0110011111: data <= 12'h001; 
        10'b0110100000: data <= 12'hfff; 
        10'b0110100001: data <= 12'h001; 
        10'b0110100010: data <= 12'h002; 
        10'b0110100011: data <= 12'h001; 
        10'b0110100100: data <= 12'h003; 
        10'b0110100101: data <= 12'h004; 
        10'b0110100110: data <= 12'h003; 
        10'b0110100111: data <= 12'h004; 
        10'b0110101000: data <= 12'h008; 
        10'b0110101001: data <= 12'h009; 
        10'b0110101010: data <= 12'h00e; 
        10'b0110101011: data <= 12'h00d; 
        10'b0110101100: data <= 12'h014; 
        10'b0110101101: data <= 12'h011; 
        10'b0110101110: data <= 12'h00c; 
        10'b0110101111: data <= 12'h009; 
        10'b0110110000: data <= 12'h00a; 
        10'b0110110001: data <= 12'h002; 
        10'b0110110010: data <= 12'h008; 
        10'b0110110011: data <= 12'h00c; 
        10'b0110110100: data <= 12'h018; 
        10'b0110110101: data <= 12'h015; 
        10'b0110110110: data <= 12'h00f; 
        10'b0110110111: data <= 12'h009; 
        10'b0110111000: data <= 12'hffe; 
        10'b0110111001: data <= 12'h003; 
        10'b0110111010: data <= 12'h006; 
        10'b0110111011: data <= 12'h001; 
        10'b0110111100: data <= 12'hffc; 
        10'b0110111101: data <= 12'h002; 
        10'b0110111110: data <= 12'h000; 
        10'b0110111111: data <= 12'h001; 
        10'b0111000000: data <= 12'h001; 
        10'b0111000001: data <= 12'h000; 
        10'b0111000010: data <= 12'h000; 
        10'b0111000011: data <= 12'hfff; 
        10'b0111000100: data <= 12'h002; 
        10'b0111000101: data <= 12'h005; 
        10'b0111000110: data <= 12'h008; 
        10'b0111000111: data <= 12'h00f; 
        10'b0111001000: data <= 12'h015; 
        10'b0111001001: data <= 12'h00f; 
        10'b0111001010: data <= 12'h004; 
        10'b0111001011: data <= 12'hfff; 
        10'b0111001100: data <= 12'h004; 
        10'b0111001101: data <= 12'h005; 
        10'b0111001110: data <= 12'h014; 
        10'b0111001111: data <= 12'h01b; 
        10'b0111010000: data <= 12'h01c; 
        10'b0111010001: data <= 12'h017; 
        10'b0111010010: data <= 12'h010; 
        10'b0111010011: data <= 12'h002; 
        10'b0111010100: data <= 12'h007; 
        10'b0111010101: data <= 12'h009; 
        10'b0111010110: data <= 12'h002; 
        10'b0111010111: data <= 12'hffe; 
        10'b0111011000: data <= 12'h000; 
        10'b0111011001: data <= 12'h001; 
        10'b0111011010: data <= 12'h002; 
        10'b0111011011: data <= 12'h002; 
        10'b0111011100: data <= 12'h002; 
        10'b0111011101: data <= 12'h002; 
        10'b0111011110: data <= 12'h003; 
        10'b0111011111: data <= 12'h000; 
        10'b0111100000: data <= 12'hffe; 
        10'b0111100001: data <= 12'hffb; 
        10'b0111100010: data <= 12'h003; 
        10'b0111100011: data <= 12'h00c; 
        10'b0111100100: data <= 12'h017; 
        10'b0111100101: data <= 12'h014; 
        10'b0111100110: data <= 12'h007; 
        10'b0111100111: data <= 12'h006; 
        10'b0111101000: data <= 12'h008; 
        10'b0111101001: data <= 12'h013; 
        10'b0111101010: data <= 12'h020; 
        10'b0111101011: data <= 12'h019; 
        10'b0111101100: data <= 12'h015; 
        10'b0111101101: data <= 12'h007; 
        10'b0111101110: data <= 12'h001; 
        10'b0111101111: data <= 12'hff9; 
        10'b0111110000: data <= 12'h002; 
        10'b0111110001: data <= 12'h001; 
        10'b0111110010: data <= 12'hffc; 
        10'b0111110011: data <= 12'hffe; 
        10'b0111110100: data <= 12'hffd; 
        10'b0111110101: data <= 12'hffe; 
        10'b0111110110: data <= 12'h003; 
        10'b0111110111: data <= 12'h003; 
        10'b0111111000: data <= 12'h002; 
        10'b0111111001: data <= 12'h003; 
        10'b0111111010: data <= 12'h002; 
        10'b0111111011: data <= 12'h000; 
        10'b0111111100: data <= 12'hffd; 
        10'b0111111101: data <= 12'hffa; 
        10'b0111111110: data <= 12'hff9; 
        10'b0111111111: data <= 12'h000; 
        10'b1000000000: data <= 12'h006; 
        10'b1000000001: data <= 12'h001; 
        10'b1000000010: data <= 12'hffb; 
        10'b1000000011: data <= 12'hffd; 
        10'b1000000100: data <= 12'h007; 
        10'b1000000101: data <= 12'h008; 
        10'b1000000110: data <= 12'h00e; 
        10'b1000000111: data <= 12'h00c; 
        10'b1000001000: data <= 12'h006; 
        10'b1000001001: data <= 12'hff6; 
        10'b1000001010: data <= 12'hff7; 
        10'b1000001011: data <= 12'hff2; 
        10'b1000001100: data <= 12'hff8; 
        10'b1000001101: data <= 12'hff8; 
        10'b1000001110: data <= 12'hff5; 
        10'b1000001111: data <= 12'hff7; 
        10'b1000010000: data <= 12'hffe; 
        10'b1000010001: data <= 12'hfff; 
        10'b1000010010: data <= 12'h001; 
        10'b1000010011: data <= 12'h000; 
        10'b1000010100: data <= 12'h002; 
        10'b1000010101: data <= 12'h003; 
        10'b1000010110: data <= 12'h001; 
        10'b1000010111: data <= 12'h001; 
        10'b1000011000: data <= 12'hffa; 
        10'b1000011001: data <= 12'hff8; 
        10'b1000011010: data <= 12'hff6; 
        10'b1000011011: data <= 12'hff1; 
        10'b1000011100: data <= 12'hfef; 
        10'b1000011101: data <= 12'hfee; 
        10'b1000011110: data <= 12'hfea; 
        10'b1000011111: data <= 12'hfeb; 
        10'b1000100000: data <= 12'hfee; 
        10'b1000100001: data <= 12'hff5; 
        10'b1000100010: data <= 12'hffd; 
        10'b1000100011: data <= 12'h003; 
        10'b1000100100: data <= 12'hff8; 
        10'b1000100101: data <= 12'hff9; 
        10'b1000100110: data <= 12'hff7; 
        10'b1000100111: data <= 12'hff4; 
        10'b1000101000: data <= 12'hff2; 
        10'b1000101001: data <= 12'hff3; 
        10'b1000101010: data <= 12'hff3; 
        10'b1000101011: data <= 12'hff7; 
        10'b1000101100: data <= 12'hffe; 
        10'b1000101101: data <= 12'h002; 
        10'b1000101110: data <= 12'h003; 
        10'b1000101111: data <= 12'h003; 
        10'b1000110000: data <= 12'h004; 
        10'b1000110001: data <= 12'h004; 
        10'b1000110010: data <= 12'h001; 
        10'b1000110011: data <= 12'h001; 
        10'b1000110100: data <= 12'hffb; 
        10'b1000110101: data <= 12'hff7; 
        10'b1000110110: data <= 12'hff4; 
        10'b1000110111: data <= 12'hfec; 
        10'b1000111000: data <= 12'hfe8; 
        10'b1000111001: data <= 12'hfe6; 
        10'b1000111010: data <= 12'hfe6; 
        10'b1000111011: data <= 12'hfed; 
        10'b1000111100: data <= 12'hff1; 
        10'b1000111101: data <= 12'hfef; 
        10'b1000111110: data <= 12'hff5; 
        10'b1000111111: data <= 12'hffa; 
        10'b1001000000: data <= 12'hffe; 
        10'b1001000001: data <= 12'hfff; 
        10'b1001000010: data <= 12'hffc; 
        10'b1001000011: data <= 12'hff6; 
        10'b1001000100: data <= 12'hff9; 
        10'b1001000101: data <= 12'hff9; 
        10'b1001000110: data <= 12'hff7; 
        10'b1001000111: data <= 12'hffb; 
        10'b1001001000: data <= 12'hffc; 
        10'b1001001001: data <= 12'h000; 
        10'b1001001010: data <= 12'h001; 
        10'b1001001011: data <= 12'h003; 
        10'b1001001100: data <= 12'h001; 
        10'b1001001101: data <= 12'h001; 
        10'b1001001110: data <= 12'h000; 
        10'b1001001111: data <= 12'h001; 
        10'b1001010000: data <= 12'h000; 
        10'b1001010001: data <= 12'hffb; 
        10'b1001010010: data <= 12'hff4; 
        10'b1001010011: data <= 12'hfef; 
        10'b1001010100: data <= 12'hff0; 
        10'b1001010101: data <= 12'hfee; 
        10'b1001010110: data <= 12'hff1; 
        10'b1001010111: data <= 12'hff5; 
        10'b1001011000: data <= 12'hff7; 
        10'b1001011001: data <= 12'hff7; 
        10'b1001011010: data <= 12'hff6; 
        10'b1001011011: data <= 12'hffb; 
        10'b1001011100: data <= 12'hffa; 
        10'b1001011101: data <= 12'h001; 
        10'b1001011110: data <= 12'hffe; 
        10'b1001011111: data <= 12'h000; 
        10'b1001100000: data <= 12'hfff; 
        10'b1001100001: data <= 12'hffa; 
        10'b1001100010: data <= 12'hffb; 
        10'b1001100011: data <= 12'hfff; 
        10'b1001100100: data <= 12'h000; 
        10'b1001100101: data <= 12'h002; 
        10'b1001100110: data <= 12'h002; 
        10'b1001100111: data <= 12'h002; 
        10'b1001101000: data <= 12'h002; 
        10'b1001101001: data <= 12'h003; 
        10'b1001101010: data <= 12'h001; 
        10'b1001101011: data <= 12'h003; 
        10'b1001101100: data <= 12'hfff; 
        10'b1001101101: data <= 12'hffd; 
        10'b1001101110: data <= 12'hffb; 
        10'b1001101111: data <= 12'hff8; 
        10'b1001110000: data <= 12'hff5; 
        10'b1001110001: data <= 12'hff9; 
        10'b1001110010: data <= 12'hff9; 
        10'b1001110011: data <= 12'hffb; 
        10'b1001110100: data <= 12'hffb; 
        10'b1001110101: data <= 12'hffc; 
        10'b1001110110: data <= 12'hffa; 
        10'b1001110111: data <= 12'hffd; 
        10'b1001111000: data <= 12'hffd; 
        10'b1001111001: data <= 12'h001; 
        10'b1001111010: data <= 12'h005; 
        10'b1001111011: data <= 12'h008; 
        10'b1001111100: data <= 12'h006; 
        10'b1001111101: data <= 12'h004; 
        10'b1001111110: data <= 12'hffd; 
        10'b1001111111: data <= 12'hffd; 
        10'b1010000000: data <= 12'h000; 
        10'b1010000001: data <= 12'h002; 
        10'b1010000010: data <= 12'h000; 
        10'b1010000011: data <= 12'h001; 
        10'b1010000100: data <= 12'h001; 
        10'b1010000101: data <= 12'h000; 
        10'b1010000110: data <= 12'h001; 
        10'b1010000111: data <= 12'h002; 
        10'b1010001000: data <= 12'h001; 
        10'b1010001001: data <= 12'h002; 
        10'b1010001010: data <= 12'hffd; 
        10'b1010001011: data <= 12'hffd; 
        10'b1010001100: data <= 12'hffc; 
        10'b1010001101: data <= 12'h002; 
        10'b1010001110: data <= 12'hffc; 
        10'b1010001111: data <= 12'h001; 
        10'b1010010000: data <= 12'hffb; 
        10'b1010010001: data <= 12'hffc; 
        10'b1010010010: data <= 12'hffd; 
        10'b1010010011: data <= 12'h000; 
        10'b1010010100: data <= 12'h001; 
        10'b1010010101: data <= 12'h003; 
        10'b1010010110: data <= 12'h009; 
        10'b1010010111: data <= 12'h009; 
        10'b1010011000: data <= 12'h008; 
        10'b1010011001: data <= 12'h003; 
        10'b1010011010: data <= 12'hfff; 
        10'b1010011011: data <= 12'h001; 
        10'b1010011100: data <= 12'h002; 
        10'b1010011101: data <= 12'h003; 
        10'b1010011110: data <= 12'h001; 
        10'b1010011111: data <= 12'h004; 
        10'b1010100000: data <= 12'h003; 
        10'b1010100001: data <= 12'h004; 
        10'b1010100010: data <= 12'h002; 
        10'b1010100011: data <= 12'h003; 
        10'b1010100100: data <= 12'h001; 
        10'b1010100101: data <= 12'h002; 
        10'b1010100110: data <= 12'h001; 
        10'b1010100111: data <= 12'hffc; 
        10'b1010101000: data <= 12'hffc; 
        10'b1010101001: data <= 12'hfff; 
        10'b1010101010: data <= 12'hffb; 
        10'b1010101011: data <= 12'hfff; 
        10'b1010101100: data <= 12'hffd; 
        10'b1010101101: data <= 12'hffd; 
        10'b1010101110: data <= 12'hffa; 
        10'b1010101111: data <= 12'hffa; 
        10'b1010110000: data <= 12'hffd; 
        10'b1010110001: data <= 12'hfff; 
        10'b1010110010: data <= 12'h001; 
        10'b1010110011: data <= 12'h005; 
        10'b1010110100: data <= 12'h004; 
        10'b1010110101: data <= 12'hfff; 
        10'b1010110110: data <= 12'h000; 
        10'b1010110111: data <= 12'h002; 
        10'b1010111000: data <= 12'h003; 
        10'b1010111001: data <= 12'h001; 
        10'b1010111010: data <= 12'h001; 
        10'b1010111011: data <= 12'h003; 
        10'b1010111100: data <= 12'h004; 
        10'b1010111101: data <= 12'h004; 
        10'b1010111110: data <= 12'h004; 
        10'b1010111111: data <= 12'h001; 
        10'b1011000000: data <= 12'h004; 
        10'b1011000001: data <= 12'h000; 
        10'b1011000010: data <= 12'hffd; 
        10'b1011000011: data <= 12'hffc; 
        10'b1011000100: data <= 12'hffa; 
        10'b1011000101: data <= 12'hff9; 
        10'b1011000110: data <= 12'hff5; 
        10'b1011000111: data <= 12'hff4; 
        10'b1011001000: data <= 12'hff5; 
        10'b1011001001: data <= 12'hff5; 
        10'b1011001010: data <= 12'hff6; 
        10'b1011001011: data <= 12'hff6; 
        10'b1011001100: data <= 12'hff3; 
        10'b1011001101: data <= 12'hff1; 
        10'b1011001110: data <= 12'hff2; 
        10'b1011001111: data <= 12'hff9; 
        10'b1011010000: data <= 12'hff9; 
        10'b1011010001: data <= 12'hffe; 
        10'b1011010010: data <= 12'h000; 
        10'b1011010011: data <= 12'h003; 
        10'b1011010100: data <= 12'h000; 
        10'b1011010101: data <= 12'h004; 
        10'b1011010110: data <= 12'h001; 
        10'b1011010111: data <= 12'h001; 
        10'b1011011000: data <= 12'h002; 
        10'b1011011001: data <= 12'h003; 
        10'b1011011010: data <= 12'h001; 
        10'b1011011011: data <= 12'h002; 
        10'b1011011100: data <= 12'h000; 
        10'b1011011101: data <= 12'hfff; 
        10'b1011011110: data <= 12'h001; 
        10'b1011011111: data <= 12'h001; 
        10'b1011100000: data <= 12'hfff; 
        10'b1011100001: data <= 12'hffc; 
        10'b1011100010: data <= 12'hff7; 
        10'b1011100011: data <= 12'hff8; 
        10'b1011100100: data <= 12'hff7; 
        10'b1011100101: data <= 12'hff4; 
        10'b1011100110: data <= 12'hff3; 
        10'b1011100111: data <= 12'hff5; 
        10'b1011101000: data <= 12'hff4; 
        10'b1011101001: data <= 12'hff6; 
        10'b1011101010: data <= 12'hff8; 
        10'b1011101011: data <= 12'hffb; 
        10'b1011101100: data <= 12'hffe; 
        10'b1011101101: data <= 12'h003; 
        10'b1011101110: data <= 12'h003; 
        10'b1011101111: data <= 12'h000; 
        10'b1011110000: data <= 12'h002; 
        10'b1011110001: data <= 12'h000; 
        10'b1011110010: data <= 12'h004; 
        10'b1011110011: data <= 12'h002; 
        10'b1011110100: data <= 12'h003; 
        10'b1011110101: data <= 12'h000; 
        10'b1011110110: data <= 12'h001; 
        10'b1011110111: data <= 12'h004; 
        10'b1011111000: data <= 12'h002; 
        10'b1011111001: data <= 12'h003; 
        10'b1011111010: data <= 12'h002; 
        10'b1011111011: data <= 12'h004; 
        10'b1011111100: data <= 12'h000; 
        10'b1011111101: data <= 12'h002; 
        10'b1011111110: data <= 12'h001; 
        10'b1011111111: data <= 12'hfff; 
        10'b1100000000: data <= 12'h000; 
        10'b1100000001: data <= 12'h000; 
        10'b1100000010: data <= 12'hffe; 
        10'b1100000011: data <= 12'h003; 
        10'b1100000100: data <= 12'hfff; 
        10'b1100000101: data <= 12'hfff; 
        10'b1100000110: data <= 12'h000; 
        10'b1100000111: data <= 12'h002; 
        10'b1100001000: data <= 12'h001; 
        10'b1100001001: data <= 12'h001; 
        10'b1100001010: data <= 12'h001; 
        10'b1100001011: data <= 12'h002; 
        10'b1100001100: data <= 12'h002; 
        10'b1100001101: data <= 12'h003; 
        10'b1100001110: data <= 12'h002; 
        10'b1100001111: data <= 12'h001; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 7) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 13'h0000; 
        10'b0000000001: data <= 13'h0001; 
        10'b0000000010: data <= 13'h0008; 
        10'b0000000011: data <= 13'h0008; 
        10'b0000000100: data <= 13'h0000; 
        10'b0000000101: data <= 13'h0000; 
        10'b0000000110: data <= 13'h0006; 
        10'b0000000111: data <= 13'h0002; 
        10'b0000001000: data <= 13'h0000; 
        10'b0000001001: data <= 13'h0001; 
        10'b0000001010: data <= 13'h0000; 
        10'b0000001011: data <= 13'h0005; 
        10'b0000001100: data <= 13'h0007; 
        10'b0000001101: data <= 13'h0004; 
        10'b0000001110: data <= 13'h0005; 
        10'b0000001111: data <= 13'h0001; 
        10'b0000010000: data <= 13'h0005; 
        10'b0000010001: data <= 13'h0007; 
        10'b0000010010: data <= 13'h0001; 
        10'b0000010011: data <= 13'h0005; 
        10'b0000010100: data <= 13'h0000; 
        10'b0000010101: data <= 13'h0003; 
        10'b0000010110: data <= 13'h0007; 
        10'b0000010111: data <= 13'h0001; 
        10'b0000011000: data <= 13'h0007; 
        10'b0000011001: data <= 13'h0001; 
        10'b0000011010: data <= 13'h0008; 
        10'b0000011011: data <= 13'h0003; 
        10'b0000011100: data <= 13'h0002; 
        10'b0000011101: data <= 13'h0004; 
        10'b0000011110: data <= 13'h0000; 
        10'b0000011111: data <= 13'h0001; 
        10'b0000100000: data <= 13'h0004; 
        10'b0000100001: data <= 13'h0009; 
        10'b0000100010: data <= 13'h0002; 
        10'b0000100011: data <= 13'h1fff; 
        10'b0000100100: data <= 13'h0005; 
        10'b0000100101: data <= 13'h0000; 
        10'b0000100110: data <= 13'h0003; 
        10'b0000100111: data <= 13'h1ffd; 
        10'b0000101000: data <= 13'h0002; 
        10'b0000101001: data <= 13'h1ffc; 
        10'b0000101010: data <= 13'h0000; 
        10'b0000101011: data <= 13'h0005; 
        10'b0000101100: data <= 13'h0006; 
        10'b0000101101: data <= 13'h0002; 
        10'b0000101110: data <= 13'h0000; 
        10'b0000101111: data <= 13'h0001; 
        10'b0000110000: data <= 13'h0006; 
        10'b0000110001: data <= 13'h0000; 
        10'b0000110010: data <= 13'h0000; 
        10'b0000110011: data <= 13'h0001; 
        10'b0000110100: data <= 13'h0005; 
        10'b0000110101: data <= 13'h0006; 
        10'b0000110110: data <= 13'h0001; 
        10'b0000110111: data <= 13'h0006; 
        10'b0000111000: data <= 13'h0007; 
        10'b0000111001: data <= 13'h0004; 
        10'b0000111010: data <= 13'h0006; 
        10'b0000111011: data <= 13'h0007; 
        10'b0000111100: data <= 13'h0006; 
        10'b0000111101: data <= 13'h0006; 
        10'b0000111110: data <= 13'h0007; 
        10'b0000111111: data <= 13'h1ffe; 
        10'b0001000000: data <= 13'h1ffd; 
        10'b0001000001: data <= 13'h0001; 
        10'b0001000010: data <= 13'h1fff; 
        10'b0001000011: data <= 13'h1ffc; 
        10'b0001000100: data <= 13'h1fef; 
        10'b0001000101: data <= 13'h1ff9; 
        10'b0001000110: data <= 13'h1ff8; 
        10'b0001000111: data <= 13'h1ff4; 
        10'b0001001000: data <= 13'h1ff7; 
        10'b0001001001: data <= 13'h1ffe; 
        10'b0001001010: data <= 13'h0002; 
        10'b0001001011: data <= 13'h0006; 
        10'b0001001100: data <= 13'h0008; 
        10'b0001001101: data <= 13'h0004; 
        10'b0001001110: data <= 13'h0007; 
        10'b0001001111: data <= 13'h0002; 
        10'b0001010000: data <= 13'h0003; 
        10'b0001010001: data <= 13'h0005; 
        10'b0001010010: data <= 13'h0000; 
        10'b0001010011: data <= 13'h0003; 
        10'b0001010100: data <= 13'h0007; 
        10'b0001010101: data <= 13'h0006; 
        10'b0001010110: data <= 13'h0002; 
        10'b0001010111: data <= 13'h0004; 
        10'b0001011000: data <= 13'h0004; 
        10'b0001011001: data <= 13'h0000; 
        10'b0001011010: data <= 13'h0005; 
        10'b0001011011: data <= 13'h1ffc; 
        10'b0001011100: data <= 13'h1ffa; 
        10'b0001011101: data <= 13'h1ffc; 
        10'b0001011110: data <= 13'h1ff1; 
        10'b0001011111: data <= 13'h1fef; 
        10'b0001100000: data <= 13'h1fe4; 
        10'b0001100001: data <= 13'h1fe6; 
        10'b0001100010: data <= 13'h1fe7; 
        10'b0001100011: data <= 13'h1fe1; 
        10'b0001100100: data <= 13'h1fec; 
        10'b0001100101: data <= 13'h1ff6; 
        10'b0001100110: data <= 13'h0001; 
        10'b0001100111: data <= 13'h0003; 
        10'b0001101000: data <= 13'h0006; 
        10'b0001101001: data <= 13'h0009; 
        10'b0001101010: data <= 13'h0002; 
        10'b0001101011: data <= 13'h0002; 
        10'b0001101100: data <= 13'h0008; 
        10'b0001101101: data <= 13'h0008; 
        10'b0001101110: data <= 13'h0003; 
        10'b0001101111: data <= 13'h0005; 
        10'b0001110000: data <= 13'h0008; 
        10'b0001110001: data <= 13'h0005; 
        10'b0001110010: data <= 13'h0006; 
        10'b0001110011: data <= 13'h0006; 
        10'b0001110100: data <= 13'h0004; 
        10'b0001110101: data <= 13'h0007; 
        10'b0001110110: data <= 13'h1ffb; 
        10'b0001110111: data <= 13'h1fff; 
        10'b0001111000: data <= 13'h1ff6; 
        10'b0001111001: data <= 13'h1ff7; 
        10'b0001111010: data <= 13'h1fe7; 
        10'b0001111011: data <= 13'h1fe8; 
        10'b0001111100: data <= 13'h1fe0; 
        10'b0001111101: data <= 13'h1fe5; 
        10'b0001111110: data <= 13'h1fdf; 
        10'b0001111111: data <= 13'h1fe4; 
        10'b0010000000: data <= 13'h1ff2; 
        10'b0010000001: data <= 13'h1ff4; 
        10'b0010000010: data <= 13'h1ff9; 
        10'b0010000011: data <= 13'h0007; 
        10'b0010000100: data <= 13'h000a; 
        10'b0010000101: data <= 13'h000b; 
        10'b0010000110: data <= 13'h000b; 
        10'b0010000111: data <= 13'h000e; 
        10'b0010001000: data <= 13'h0004; 
        10'b0010001001: data <= 13'h0008; 
        10'b0010001010: data <= 13'h0002; 
        10'b0010001011: data <= 13'h0001; 
        10'b0010001100: data <= 13'h0008; 
        10'b0010001101: data <= 13'h0002; 
        10'b0010001110: data <= 13'h0006; 
        10'b0010001111: data <= 13'h0002; 
        10'b0010010000: data <= 13'h0005; 
        10'b0010010001: data <= 13'h0001; 
        10'b0010010010: data <= 13'h0004; 
        10'b0010010011: data <= 13'h1ffb; 
        10'b0010010100: data <= 13'h0001; 
        10'b0010010101: data <= 13'h1ffb; 
        10'b0010010110: data <= 13'h1fee; 
        10'b0010010111: data <= 13'h1ff4; 
        10'b0010011000: data <= 13'h1feb; 
        10'b0010011001: data <= 13'h1fe6; 
        10'b0010011010: data <= 13'h1fee; 
        10'b0010011011: data <= 13'h1ff1; 
        10'b0010011100: data <= 13'h1ffe; 
        10'b0010011101: data <= 13'h0002; 
        10'b0010011110: data <= 13'h1ffc; 
        10'b0010011111: data <= 13'h0006; 
        10'b0010100000: data <= 13'h0007; 
        10'b0010100001: data <= 13'h000a; 
        10'b0010100010: data <= 13'h0017; 
        10'b0010100011: data <= 13'h001a; 
        10'b0010100100: data <= 13'h000e; 
        10'b0010100101: data <= 13'h1fff; 
        10'b0010100110: data <= 13'h0002; 
        10'b0010100111: data <= 13'h0001; 
        10'b0010101000: data <= 13'h0008; 
        10'b0010101001: data <= 13'h0009; 
        10'b0010101010: data <= 13'h0003; 
        10'b0010101011: data <= 13'h0007; 
        10'b0010101100: data <= 13'h0007; 
        10'b0010101101: data <= 13'h0006; 
        10'b0010101110: data <= 13'h0006; 
        10'b0010101111: data <= 13'h0000; 
        10'b0010110000: data <= 13'h1fff; 
        10'b0010110001: data <= 13'h1ff9; 
        10'b0010110010: data <= 13'h1ff2; 
        10'b0010110011: data <= 13'h1fe7; 
        10'b0010110100: data <= 13'h1fda; 
        10'b0010110101: data <= 13'h1fd3; 
        10'b0010110110: data <= 13'h1fd1; 
        10'b0010110111: data <= 13'h1fd7; 
        10'b0010111000: data <= 13'h1fd6; 
        10'b0010111001: data <= 13'h1fe7; 
        10'b0010111010: data <= 13'h1fe6; 
        10'b0010111011: data <= 13'h1ff4; 
        10'b0010111100: data <= 13'h1ff8; 
        10'b0010111101: data <= 13'h1fff; 
        10'b0010111110: data <= 13'h0021; 
        10'b0010111111: data <= 13'h0023; 
        10'b0011000000: data <= 13'h000d; 
        10'b0011000001: data <= 13'h000a; 
        10'b0011000010: data <= 13'h0007; 
        10'b0011000011: data <= 13'h0000; 
        10'b0011000100: data <= 13'h0004; 
        10'b0011000101: data <= 13'h0002; 
        10'b0011000110: data <= 13'h0003; 
        10'b0011000111: data <= 13'h0005; 
        10'b0011001000: data <= 13'h0003; 
        10'b0011001001: data <= 13'h0006; 
        10'b0011001010: data <= 13'h1ffc; 
        10'b0011001011: data <= 13'h1fff; 
        10'b0011001100: data <= 13'h1ffc; 
        10'b0011001101: data <= 13'h1ff6; 
        10'b0011001110: data <= 13'h1fe7; 
        10'b0011001111: data <= 13'h1fda; 
        10'b0011010000: data <= 13'h1fce; 
        10'b0011010001: data <= 13'h1fdd; 
        10'b0011010010: data <= 13'h1fd4; 
        10'b0011010011: data <= 13'h1fd4; 
        10'b0011010100: data <= 13'h1fd2; 
        10'b0011010101: data <= 13'h1fe3; 
        10'b0011010110: data <= 13'h1fe2; 
        10'b0011010111: data <= 13'h1feb; 
        10'b0011011000: data <= 13'h1fe8; 
        10'b0011011001: data <= 13'h1ff5; 
        10'b0011011010: data <= 13'h0014; 
        10'b0011011011: data <= 13'h001c; 
        10'b0011011100: data <= 13'h000f; 
        10'b0011011101: data <= 13'h0008; 
        10'b0011011110: data <= 13'h0008; 
        10'b0011011111: data <= 13'h0005; 
        10'b0011100000: data <= 13'h0007; 
        10'b0011100001: data <= 13'h0006; 
        10'b0011100010: data <= 13'h0008; 
        10'b0011100011: data <= 13'h0002; 
        10'b0011100100: data <= 13'h0002; 
        10'b0011100101: data <= 13'h0003; 
        10'b0011100110: data <= 13'h0002; 
        10'b0011100111: data <= 13'h1ffe; 
        10'b0011101000: data <= 13'h1fed; 
        10'b0011101001: data <= 13'h1ff7; 
        10'b0011101010: data <= 13'h1ff4; 
        10'b0011101011: data <= 13'h1fe7; 
        10'b0011101100: data <= 13'h1fdc; 
        10'b0011101101: data <= 13'h1fe9; 
        10'b0011101110: data <= 13'h1fcb; 
        10'b0011101111: data <= 13'h1fca; 
        10'b0011110000: data <= 13'h1fd6; 
        10'b0011110001: data <= 13'h1fe6; 
        10'b0011110010: data <= 13'h1fe8; 
        10'b0011110011: data <= 13'h1ff9; 
        10'b0011110100: data <= 13'h1ff2; 
        10'b0011110101: data <= 13'h1ff2; 
        10'b0011110110: data <= 13'h0009; 
        10'b0011110111: data <= 13'h000e; 
        10'b0011111000: data <= 13'h000b; 
        10'b0011111001: data <= 13'h0002; 
        10'b0011111010: data <= 13'h0003; 
        10'b0011111011: data <= 13'h0005; 
        10'b0011111100: data <= 13'h0009; 
        10'b0011111101: data <= 13'h0007; 
        10'b0011111110: data <= 13'h0007; 
        10'b0011111111: data <= 13'h0001; 
        10'b0100000000: data <= 13'h1ffb; 
        10'b0100000001: data <= 13'h0000; 
        10'b0100000010: data <= 13'h1ff5; 
        10'b0100000011: data <= 13'h1ff8; 
        10'b0100000100: data <= 13'h1ffb; 
        10'b0100000101: data <= 13'h1ffe; 
        10'b0100000110: data <= 13'h1ffa; 
        10'b0100000111: data <= 13'h1ff8; 
        10'b0100001000: data <= 13'h1ff8; 
        10'b0100001001: data <= 13'h1feb; 
        10'b0100001010: data <= 13'h1fb4; 
        10'b0100001011: data <= 13'h1fc7; 
        10'b0100001100: data <= 13'h1ff2; 
        10'b0100001101: data <= 13'h1ff6; 
        10'b0100001110: data <= 13'h1ffd; 
        10'b0100001111: data <= 13'h0002; 
        10'b0100010000: data <= 13'h1ff8; 
        10'b0100010001: data <= 13'h1ff8; 
        10'b0100010010: data <= 13'h0004; 
        10'b0100010011: data <= 13'h0001; 
        10'b0100010100: data <= 13'h1ff7; 
        10'b0100010101: data <= 13'h1ff7; 
        10'b0100010110: data <= 13'h1ffc; 
        10'b0100010111: data <= 13'h0006; 
        10'b0100011000: data <= 13'h0005; 
        10'b0100011001: data <= 13'h0003; 
        10'b0100011010: data <= 13'h0003; 
        10'b0100011011: data <= 13'h0001; 
        10'b0100011100: data <= 13'h0004; 
        10'b0100011101: data <= 13'h1ff6; 
        10'b0100011110: data <= 13'h1fef; 
        10'b0100011111: data <= 13'h1ff8; 
        10'b0100100000: data <= 13'h0002; 
        10'b0100100001: data <= 13'h0016; 
        10'b0100100010: data <= 13'h000d; 
        10'b0100100011: data <= 13'h000a; 
        10'b0100100100: data <= 13'h000c; 
        10'b0100100101: data <= 13'h1fe3; 
        10'b0100100110: data <= 13'h1fb0; 
        10'b0100100111: data <= 13'h1fe8; 
        10'b0100101000: data <= 13'h0003; 
        10'b0100101001: data <= 13'h1ffc; 
        10'b0100101010: data <= 13'h1ffd; 
        10'b0100101011: data <= 13'h0003; 
        10'b0100101100: data <= 13'h1ff0; 
        10'b0100101101: data <= 13'h1ff5; 
        10'b0100101110: data <= 13'h1ffe; 
        10'b0100101111: data <= 13'h1fef; 
        10'b0100110000: data <= 13'h1ff6; 
        10'b0100110001: data <= 13'h1ffa; 
        10'b0100110010: data <= 13'h0005; 
        10'b0100110011: data <= 13'h0008; 
        10'b0100110100: data <= 13'h0006; 
        10'b0100110101: data <= 13'h0006; 
        10'b0100110110: data <= 13'h0005; 
        10'b0100110111: data <= 13'h1ffd; 
        10'b0100111000: data <= 13'h1fff; 
        10'b0100111001: data <= 13'h1ffa; 
        10'b0100111010: data <= 13'h1ffa; 
        10'b0100111011: data <= 13'h0005; 
        10'b0100111100: data <= 13'h0010; 
        10'b0100111101: data <= 13'h001c; 
        10'b0100111110: data <= 13'h0026; 
        10'b0100111111: data <= 13'h0018; 
        10'b0101000000: data <= 13'h001b; 
        10'b0101000001: data <= 13'h1fd4; 
        10'b0101000010: data <= 13'h1fc4; 
        10'b0101000011: data <= 13'h0008; 
        10'b0101000100: data <= 13'h001f; 
        10'b0101000101: data <= 13'h0005; 
        10'b0101000110: data <= 13'h1ffe; 
        10'b0101000111: data <= 13'h1ffb; 
        10'b0101001000: data <= 13'h1fef; 
        10'b0101001001: data <= 13'h1ff1; 
        10'b0101001010: data <= 13'h1ff9; 
        10'b0101001011: data <= 13'h1ff2; 
        10'b0101001100: data <= 13'h1ff1; 
        10'b0101001101: data <= 13'h1fff; 
        10'b0101001110: data <= 13'h1fff; 
        10'b0101001111: data <= 13'h0002; 
        10'b0101010000: data <= 13'h0006; 
        10'b0101010001: data <= 13'h0005; 
        10'b0101010010: data <= 13'h0003; 
        10'b0101010011: data <= 13'h0004; 
        10'b0101010100: data <= 13'h0000; 
        10'b0101010101: data <= 13'h1ffa; 
        10'b0101010110: data <= 13'h0010; 
        10'b0101010111: data <= 13'h001a; 
        10'b0101011000: data <= 13'h0029; 
        10'b0101011001: data <= 13'h0024; 
        10'b0101011010: data <= 13'h003c; 
        10'b0101011011: data <= 13'h0044; 
        10'b0101011100: data <= 13'h0040; 
        10'b0101011101: data <= 13'h1fff; 
        10'b0101011110: data <= 13'h1fe0; 
        10'b0101011111: data <= 13'h0019; 
        10'b0101100000: data <= 13'h0029; 
        10'b0101100001: data <= 13'h0005; 
        10'b0101100010: data <= 13'h0002; 
        10'b0101100011: data <= 13'h0006; 
        10'b0101100100: data <= 13'h1fff; 
        10'b0101100101: data <= 13'h0001; 
        10'b0101100110: data <= 13'h1ffe; 
        10'b0101100111: data <= 13'h1ff7; 
        10'b0101101000: data <= 13'h1ff8; 
        10'b0101101001: data <= 13'h1ffe; 
        10'b0101101010: data <= 13'h0009; 
        10'b0101101011: data <= 13'h0005; 
        10'b0101101100: data <= 13'h0001; 
        10'b0101101101: data <= 13'h0006; 
        10'b0101101110: data <= 13'h0001; 
        10'b0101101111: data <= 13'h0002; 
        10'b0101110000: data <= 13'h0007; 
        10'b0101110001: data <= 13'h0013; 
        10'b0101110010: data <= 13'h0027; 
        10'b0101110011: data <= 13'h002e; 
        10'b0101110100: data <= 13'h0035; 
        10'b0101110101: data <= 13'h002c; 
        10'b0101110110: data <= 13'h0033; 
        10'b0101110111: data <= 13'h0054; 
        10'b0101111000: data <= 13'h003f; 
        10'b0101111001: data <= 13'h0001; 
        10'b0101111010: data <= 13'h1ff7; 
        10'b0101111011: data <= 13'h001d; 
        10'b0101111100: data <= 13'h001e; 
        10'b0101111101: data <= 13'h0021; 
        10'b0101111110: data <= 13'h0017; 
        10'b0101111111: data <= 13'h000a; 
        10'b0110000000: data <= 13'h0017; 
        10'b0110000001: data <= 13'h0011; 
        10'b0110000010: data <= 13'h0008; 
        10'b0110000011: data <= 13'h1ffb; 
        10'b0110000100: data <= 13'h1ffc; 
        10'b0110000101: data <= 13'h0000; 
        10'b0110000110: data <= 13'h0007; 
        10'b0110000111: data <= 13'h0005; 
        10'b0110001000: data <= 13'h0001; 
        10'b0110001001: data <= 13'h0007; 
        10'b0110001010: data <= 13'h0001; 
        10'b0110001011: data <= 13'h0009; 
        10'b0110001100: data <= 13'h0011; 
        10'b0110001101: data <= 13'h0023; 
        10'b0110001110: data <= 13'h0030; 
        10'b0110001111: data <= 13'h0035; 
        10'b0110010000: data <= 13'h0027; 
        10'b0110010001: data <= 13'h0025; 
        10'b0110010010: data <= 13'h002d; 
        10'b0110010011: data <= 13'h0037; 
        10'b0110010100: data <= 13'h0028; 
        10'b0110010101: data <= 13'h0003; 
        10'b0110010110: data <= 13'h1ffa; 
        10'b0110010111: data <= 13'h000b; 
        10'b0110011000: data <= 13'h0022; 
        10'b0110011001: data <= 13'h0037; 
        10'b0110011010: data <= 13'h0025; 
        10'b0110011011: data <= 13'h0022; 
        10'b0110011100: data <= 13'h0013; 
        10'b0110011101: data <= 13'h000d; 
        10'b0110011110: data <= 13'h0004; 
        10'b0110011111: data <= 13'h0002; 
        10'b0110100000: data <= 13'h1fff; 
        10'b0110100001: data <= 13'h0002; 
        10'b0110100010: data <= 13'h0004; 
        10'b0110100011: data <= 13'h0002; 
        10'b0110100100: data <= 13'h0006; 
        10'b0110100101: data <= 13'h0009; 
        10'b0110100110: data <= 13'h0006; 
        10'b0110100111: data <= 13'h0007; 
        10'b0110101000: data <= 13'h000f; 
        10'b0110101001: data <= 13'h0012; 
        10'b0110101010: data <= 13'h001b; 
        10'b0110101011: data <= 13'h0019; 
        10'b0110101100: data <= 13'h0028; 
        10'b0110101101: data <= 13'h0023; 
        10'b0110101110: data <= 13'h0018; 
        10'b0110101111: data <= 13'h0012; 
        10'b0110110000: data <= 13'h0015; 
        10'b0110110001: data <= 13'h0004; 
        10'b0110110010: data <= 13'h0011; 
        10'b0110110011: data <= 13'h0017; 
        10'b0110110100: data <= 13'h0030; 
        10'b0110110101: data <= 13'h002b; 
        10'b0110110110: data <= 13'h001f; 
        10'b0110110111: data <= 13'h0012; 
        10'b0110111000: data <= 13'h1ffb; 
        10'b0110111001: data <= 13'h0007; 
        10'b0110111010: data <= 13'h000c; 
        10'b0110111011: data <= 13'h0001; 
        10'b0110111100: data <= 13'h1ff9; 
        10'b0110111101: data <= 13'h0004; 
        10'b0110111110: data <= 13'h0001; 
        10'b0110111111: data <= 13'h0002; 
        10'b0111000000: data <= 13'h0003; 
        10'b0111000001: data <= 13'h0000; 
        10'b0111000010: data <= 13'h0000; 
        10'b0111000011: data <= 13'h1fff; 
        10'b0111000100: data <= 13'h0004; 
        10'b0111000101: data <= 13'h000a; 
        10'b0111000110: data <= 13'h0011; 
        10'b0111000111: data <= 13'h001e; 
        10'b0111001000: data <= 13'h002b; 
        10'b0111001001: data <= 13'h001f; 
        10'b0111001010: data <= 13'h0008; 
        10'b0111001011: data <= 13'h1fff; 
        10'b0111001100: data <= 13'h0008; 
        10'b0111001101: data <= 13'h000a; 
        10'b0111001110: data <= 13'h0027; 
        10'b0111001111: data <= 13'h0037; 
        10'b0111010000: data <= 13'h0038; 
        10'b0111010001: data <= 13'h002f; 
        10'b0111010010: data <= 13'h0020; 
        10'b0111010011: data <= 13'h0004; 
        10'b0111010100: data <= 13'h000d; 
        10'b0111010101: data <= 13'h0013; 
        10'b0111010110: data <= 13'h0004; 
        10'b0111010111: data <= 13'h1ffd; 
        10'b0111011000: data <= 13'h1fff; 
        10'b0111011001: data <= 13'h0002; 
        10'b0111011010: data <= 13'h0003; 
        10'b0111011011: data <= 13'h0004; 
        10'b0111011100: data <= 13'h0003; 
        10'b0111011101: data <= 13'h0003; 
        10'b0111011110: data <= 13'h0006; 
        10'b0111011111: data <= 13'h0000; 
        10'b0111100000: data <= 13'h1ffb; 
        10'b0111100001: data <= 13'h1ff7; 
        10'b0111100010: data <= 13'h0005; 
        10'b0111100011: data <= 13'h0017; 
        10'b0111100100: data <= 13'h002d; 
        10'b0111100101: data <= 13'h0027; 
        10'b0111100110: data <= 13'h000e; 
        10'b0111100111: data <= 13'h000b; 
        10'b0111101000: data <= 13'h0010; 
        10'b0111101001: data <= 13'h0027; 
        10'b0111101010: data <= 13'h0040; 
        10'b0111101011: data <= 13'h0033; 
        10'b0111101100: data <= 13'h002a; 
        10'b0111101101: data <= 13'h000d; 
        10'b0111101110: data <= 13'h0002; 
        10'b0111101111: data <= 13'h1ff2; 
        10'b0111110000: data <= 13'h0004; 
        10'b0111110001: data <= 13'h0002; 
        10'b0111110010: data <= 13'h1ff7; 
        10'b0111110011: data <= 13'h1ffc; 
        10'b0111110100: data <= 13'h1ffa; 
        10'b0111110101: data <= 13'h1ffd; 
        10'b0111110110: data <= 13'h0006; 
        10'b0111110111: data <= 13'h0007; 
        10'b0111111000: data <= 13'h0003; 
        10'b0111111001: data <= 13'h0005; 
        10'b0111111010: data <= 13'h0005; 
        10'b0111111011: data <= 13'h0001; 
        10'b0111111100: data <= 13'h1ffb; 
        10'b0111111101: data <= 13'h1ff5; 
        10'b0111111110: data <= 13'h1ff3; 
        10'b0111111111: data <= 13'h0000; 
        10'b1000000000: data <= 13'h000c; 
        10'b1000000001: data <= 13'h0003; 
        10'b1000000010: data <= 13'h1ff7; 
        10'b1000000011: data <= 13'h1ffa; 
        10'b1000000100: data <= 13'h000f; 
        10'b1000000101: data <= 13'h0011; 
        10'b1000000110: data <= 13'h001c; 
        10'b1000000111: data <= 13'h0018; 
        10'b1000001000: data <= 13'h000d; 
        10'b1000001001: data <= 13'h1fed; 
        10'b1000001010: data <= 13'h1fee; 
        10'b1000001011: data <= 13'h1fe5; 
        10'b1000001100: data <= 13'h1ff0; 
        10'b1000001101: data <= 13'h1fef; 
        10'b1000001110: data <= 13'h1fea; 
        10'b1000001111: data <= 13'h1fef; 
        10'b1000010000: data <= 13'h1ffc; 
        10'b1000010001: data <= 13'h1ffe; 
        10'b1000010010: data <= 13'h0002; 
        10'b1000010011: data <= 13'h0000; 
        10'b1000010100: data <= 13'h0003; 
        10'b1000010101: data <= 13'h0006; 
        10'b1000010110: data <= 13'h0002; 
        10'b1000010111: data <= 13'h0001; 
        10'b1000011000: data <= 13'h1ff4; 
        10'b1000011001: data <= 13'h1ff1; 
        10'b1000011010: data <= 13'h1fec; 
        10'b1000011011: data <= 13'h1fe1; 
        10'b1000011100: data <= 13'h1fde; 
        10'b1000011101: data <= 13'h1fdb; 
        10'b1000011110: data <= 13'h1fd5; 
        10'b1000011111: data <= 13'h1fd7; 
        10'b1000100000: data <= 13'h1fdb; 
        10'b1000100001: data <= 13'h1feb; 
        10'b1000100010: data <= 13'h1ffa; 
        10'b1000100011: data <= 13'h0006; 
        10'b1000100100: data <= 13'h1fef; 
        10'b1000100101: data <= 13'h1ff2; 
        10'b1000100110: data <= 13'h1fee; 
        10'b1000100111: data <= 13'h1fe8; 
        10'b1000101000: data <= 13'h1fe5; 
        10'b1000101001: data <= 13'h1fe7; 
        10'b1000101010: data <= 13'h1fe6; 
        10'b1000101011: data <= 13'h1fef; 
        10'b1000101100: data <= 13'h1ffb; 
        10'b1000101101: data <= 13'h0003; 
        10'b1000101110: data <= 13'h0006; 
        10'b1000101111: data <= 13'h0006; 
        10'b1000110000: data <= 13'h0009; 
        10'b1000110001: data <= 13'h0008; 
        10'b1000110010: data <= 13'h0002; 
        10'b1000110011: data <= 13'h0001; 
        10'b1000110100: data <= 13'h1ff6; 
        10'b1000110101: data <= 13'h1fef; 
        10'b1000110110: data <= 13'h1fe7; 
        10'b1000110111: data <= 13'h1fd7; 
        10'b1000111000: data <= 13'h1fd0; 
        10'b1000111001: data <= 13'h1fcd; 
        10'b1000111010: data <= 13'h1fcc; 
        10'b1000111011: data <= 13'h1fda; 
        10'b1000111100: data <= 13'h1fe1; 
        10'b1000111101: data <= 13'h1fde; 
        10'b1000111110: data <= 13'h1fea; 
        10'b1000111111: data <= 13'h1ff5; 
        10'b1001000000: data <= 13'h1ffc; 
        10'b1001000001: data <= 13'h1ffe; 
        10'b1001000010: data <= 13'h1ff7; 
        10'b1001000011: data <= 13'h1fed; 
        10'b1001000100: data <= 13'h1ff3; 
        10'b1001000101: data <= 13'h1ff1; 
        10'b1001000110: data <= 13'h1fee; 
        10'b1001000111: data <= 13'h1ff7; 
        10'b1001001000: data <= 13'h1ff7; 
        10'b1001001001: data <= 13'h0001; 
        10'b1001001010: data <= 13'h0002; 
        10'b1001001011: data <= 13'h0006; 
        10'b1001001100: data <= 13'h0002; 
        10'b1001001101: data <= 13'h0003; 
        10'b1001001110: data <= 13'h0001; 
        10'b1001001111: data <= 13'h0001; 
        10'b1001010000: data <= 13'h0000; 
        10'b1001010001: data <= 13'h1ff6; 
        10'b1001010010: data <= 13'h1fe7; 
        10'b1001010011: data <= 13'h1fde; 
        10'b1001010100: data <= 13'h1fe1; 
        10'b1001010101: data <= 13'h1fdd; 
        10'b1001010110: data <= 13'h1fe1; 
        10'b1001010111: data <= 13'h1fe9; 
        10'b1001011000: data <= 13'h1fed; 
        10'b1001011001: data <= 13'h1fee; 
        10'b1001011010: data <= 13'h1fec; 
        10'b1001011011: data <= 13'h1ff7; 
        10'b1001011100: data <= 13'h1ff4; 
        10'b1001011101: data <= 13'h0002; 
        10'b1001011110: data <= 13'h1ffc; 
        10'b1001011111: data <= 13'h0001; 
        10'b1001100000: data <= 13'h1ffe; 
        10'b1001100001: data <= 13'h1ff4; 
        10'b1001100010: data <= 13'h1ff6; 
        10'b1001100011: data <= 13'h1ffe; 
        10'b1001100100: data <= 13'h0000; 
        10'b1001100101: data <= 13'h0004; 
        10'b1001100110: data <= 13'h0005; 
        10'b1001100111: data <= 13'h0005; 
        10'b1001101000: data <= 13'h0004; 
        10'b1001101001: data <= 13'h0005; 
        10'b1001101010: data <= 13'h0002; 
        10'b1001101011: data <= 13'h0006; 
        10'b1001101100: data <= 13'h1fff; 
        10'b1001101101: data <= 13'h1ffb; 
        10'b1001101110: data <= 13'h1ff6; 
        10'b1001101111: data <= 13'h1fef; 
        10'b1001110000: data <= 13'h1fe9; 
        10'b1001110001: data <= 13'h1ff2; 
        10'b1001110010: data <= 13'h1ff2; 
        10'b1001110011: data <= 13'h1ff6; 
        10'b1001110100: data <= 13'h1ff6; 
        10'b1001110101: data <= 13'h1ff7; 
        10'b1001110110: data <= 13'h1ff5; 
        10'b1001110111: data <= 13'h1ff9; 
        10'b1001111000: data <= 13'h1ff9; 
        10'b1001111001: data <= 13'h0002; 
        10'b1001111010: data <= 13'h000a; 
        10'b1001111011: data <= 13'h0010; 
        10'b1001111100: data <= 13'h000d; 
        10'b1001111101: data <= 13'h0008; 
        10'b1001111110: data <= 13'h1ffb; 
        10'b1001111111: data <= 13'h1ffb; 
        10'b1010000000: data <= 13'h0000; 
        10'b1010000001: data <= 13'h0004; 
        10'b1010000010: data <= 13'h0001; 
        10'b1010000011: data <= 13'h0003; 
        10'b1010000100: data <= 13'h0003; 
        10'b1010000101: data <= 13'h0000; 
        10'b1010000110: data <= 13'h0002; 
        10'b1010000111: data <= 13'h0005; 
        10'b1010001000: data <= 13'h0003; 
        10'b1010001001: data <= 13'h0003; 
        10'b1010001010: data <= 13'h1ffb; 
        10'b1010001011: data <= 13'h1ffa; 
        10'b1010001100: data <= 13'h1ff8; 
        10'b1010001101: data <= 13'h0004; 
        10'b1010001110: data <= 13'h1ff7; 
        10'b1010001111: data <= 13'h0001; 
        10'b1010010000: data <= 13'h1ff7; 
        10'b1010010001: data <= 13'h1ff9; 
        10'b1010010010: data <= 13'h1ff9; 
        10'b1010010011: data <= 13'h1fff; 
        10'b1010010100: data <= 13'h0002; 
        10'b1010010101: data <= 13'h0006; 
        10'b1010010110: data <= 13'h0013; 
        10'b1010010111: data <= 13'h0012; 
        10'b1010011000: data <= 13'h0010; 
        10'b1010011001: data <= 13'h0007; 
        10'b1010011010: data <= 13'h1ffd; 
        10'b1010011011: data <= 13'h0002; 
        10'b1010011100: data <= 13'h0004; 
        10'b1010011101: data <= 13'h0006; 
        10'b1010011110: data <= 13'h0002; 
        10'b1010011111: data <= 13'h0007; 
        10'b1010100000: data <= 13'h0005; 
        10'b1010100001: data <= 13'h0008; 
        10'b1010100010: data <= 13'h0004; 
        10'b1010100011: data <= 13'h0006; 
        10'b1010100100: data <= 13'h0001; 
        10'b1010100101: data <= 13'h0005; 
        10'b1010100110: data <= 13'h0002; 
        10'b1010100111: data <= 13'h1ff7; 
        10'b1010101000: data <= 13'h1ff7; 
        10'b1010101001: data <= 13'h1ffd; 
        10'b1010101010: data <= 13'h1ff7; 
        10'b1010101011: data <= 13'h1ffe; 
        10'b1010101100: data <= 13'h1ff9; 
        10'b1010101101: data <= 13'h1ffa; 
        10'b1010101110: data <= 13'h1ff5; 
        10'b1010101111: data <= 13'h1ff3; 
        10'b1010110000: data <= 13'h1ffa; 
        10'b1010110001: data <= 13'h1ffd; 
        10'b1010110010: data <= 13'h0001; 
        10'b1010110011: data <= 13'h000a; 
        10'b1010110100: data <= 13'h0007; 
        10'b1010110101: data <= 13'h1ffd; 
        10'b1010110110: data <= 13'h1fff; 
        10'b1010110111: data <= 13'h0004; 
        10'b1010111000: data <= 13'h0006; 
        10'b1010111001: data <= 13'h0001; 
        10'b1010111010: data <= 13'h0002; 
        10'b1010111011: data <= 13'h0005; 
        10'b1010111100: data <= 13'h0008; 
        10'b1010111101: data <= 13'h0008; 
        10'b1010111110: data <= 13'h0007; 
        10'b1010111111: data <= 13'h0002; 
        10'b1011000000: data <= 13'h0007; 
        10'b1011000001: data <= 13'h0000; 
        10'b1011000010: data <= 13'h1ffb; 
        10'b1011000011: data <= 13'h1ff8; 
        10'b1011000100: data <= 13'h1ff4; 
        10'b1011000101: data <= 13'h1ff3; 
        10'b1011000110: data <= 13'h1fea; 
        10'b1011000111: data <= 13'h1fe8; 
        10'b1011001000: data <= 13'h1fe9; 
        10'b1011001001: data <= 13'h1fe9; 
        10'b1011001010: data <= 13'h1fed; 
        10'b1011001011: data <= 13'h1feb; 
        10'b1011001100: data <= 13'h1fe5; 
        10'b1011001101: data <= 13'h1fe2; 
        10'b1011001110: data <= 13'h1fe5; 
        10'b1011001111: data <= 13'h1ff1; 
        10'b1011010000: data <= 13'h1ff2; 
        10'b1011010001: data <= 13'h1ffb; 
        10'b1011010010: data <= 13'h0000; 
        10'b1011010011: data <= 13'h0005; 
        10'b1011010100: data <= 13'h0000; 
        10'b1011010101: data <= 13'h0007; 
        10'b1011010110: data <= 13'h0003; 
        10'b1011010111: data <= 13'h0003; 
        10'b1011011000: data <= 13'h0004; 
        10'b1011011001: data <= 13'h0005; 
        10'b1011011010: data <= 13'h0001; 
        10'b1011011011: data <= 13'h0004; 
        10'b1011011100: data <= 13'h0000; 
        10'b1011011101: data <= 13'h1fff; 
        10'b1011011110: data <= 13'h0002; 
        10'b1011011111: data <= 13'h0002; 
        10'b1011100000: data <= 13'h1ffe; 
        10'b1011100001: data <= 13'h1ff8; 
        10'b1011100010: data <= 13'h1fee; 
        10'b1011100011: data <= 13'h1ff0; 
        10'b1011100100: data <= 13'h1fee; 
        10'b1011100101: data <= 13'h1fe7; 
        10'b1011100110: data <= 13'h1fe5; 
        10'b1011100111: data <= 13'h1feb; 
        10'b1011101000: data <= 13'h1fe8; 
        10'b1011101001: data <= 13'h1fec; 
        10'b1011101010: data <= 13'h1fef; 
        10'b1011101011: data <= 13'h1ff6; 
        10'b1011101100: data <= 13'h1ffc; 
        10'b1011101101: data <= 13'h0005; 
        10'b1011101110: data <= 13'h0005; 
        10'b1011101111: data <= 13'h0001; 
        10'b1011110000: data <= 13'h0003; 
        10'b1011110001: data <= 13'h0001; 
        10'b1011110010: data <= 13'h0009; 
        10'b1011110011: data <= 13'h0004; 
        10'b1011110100: data <= 13'h0005; 
        10'b1011110101: data <= 13'h0001; 
        10'b1011110110: data <= 13'h0001; 
        10'b1011110111: data <= 13'h0008; 
        10'b1011111000: data <= 13'h0003; 
        10'b1011111001: data <= 13'h0007; 
        10'b1011111010: data <= 13'h0003; 
        10'b1011111011: data <= 13'h0008; 
        10'b1011111100: data <= 13'h0000; 
        10'b1011111101: data <= 13'h0004; 
        10'b1011111110: data <= 13'h0002; 
        10'b1011111111: data <= 13'h1fff; 
        10'b1100000000: data <= 13'h1fff; 
        10'b1100000001: data <= 13'h0000; 
        10'b1100000010: data <= 13'h1ffd; 
        10'b1100000011: data <= 13'h0007; 
        10'b1100000100: data <= 13'h1ffe; 
        10'b1100000101: data <= 13'h1ffe; 
        10'b1100000110: data <= 13'h1fff; 
        10'b1100000111: data <= 13'h0004; 
        10'b1100001000: data <= 13'h0003; 
        10'b1100001001: data <= 13'h0003; 
        10'b1100001010: data <= 13'h0003; 
        10'b1100001011: data <= 13'h0005; 
        10'b1100001100: data <= 13'h0005; 
        10'b1100001101: data <= 13'h0006; 
        10'b1100001110: data <= 13'h0004; 
        10'b1100001111: data <= 13'h0003; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 8) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 14'h0000; 
        10'b0000000001: data <= 14'h0002; 
        10'b0000000010: data <= 14'h000f; 
        10'b0000000011: data <= 14'h000f; 
        10'b0000000100: data <= 14'h0000; 
        10'b0000000101: data <= 14'h0000; 
        10'b0000000110: data <= 14'h000c; 
        10'b0000000111: data <= 14'h0003; 
        10'b0000001000: data <= 14'h0001; 
        10'b0000001001: data <= 14'h0002; 
        10'b0000001010: data <= 14'h0000; 
        10'b0000001011: data <= 14'h000b; 
        10'b0000001100: data <= 14'h000e; 
        10'b0000001101: data <= 14'h0008; 
        10'b0000001110: data <= 14'h000b; 
        10'b0000001111: data <= 14'h0001; 
        10'b0000010000: data <= 14'h000a; 
        10'b0000010001: data <= 14'h000e; 
        10'b0000010010: data <= 14'h0003; 
        10'b0000010011: data <= 14'h000b; 
        10'b0000010100: data <= 14'h0001; 
        10'b0000010101: data <= 14'h0006; 
        10'b0000010110: data <= 14'h000f; 
        10'b0000010111: data <= 14'h0001; 
        10'b0000011000: data <= 14'h000f; 
        10'b0000011001: data <= 14'h0002; 
        10'b0000011010: data <= 14'h0010; 
        10'b0000011011: data <= 14'h0007; 
        10'b0000011100: data <= 14'h0004; 
        10'b0000011101: data <= 14'h0007; 
        10'b0000011110: data <= 14'h0000; 
        10'b0000011111: data <= 14'h0001; 
        10'b0000100000: data <= 14'h0007; 
        10'b0000100001: data <= 14'h0012; 
        10'b0000100010: data <= 14'h0004; 
        10'b0000100011: data <= 14'h3ffd; 
        10'b0000100100: data <= 14'h000a; 
        10'b0000100101: data <= 14'h0000; 
        10'b0000100110: data <= 14'h0007; 
        10'b0000100111: data <= 14'h3ffb; 
        10'b0000101000: data <= 14'h0005; 
        10'b0000101001: data <= 14'h3ff9; 
        10'b0000101010: data <= 14'h0000; 
        10'b0000101011: data <= 14'h000a; 
        10'b0000101100: data <= 14'h000b; 
        10'b0000101101: data <= 14'h0003; 
        10'b0000101110: data <= 14'h0000; 
        10'b0000101111: data <= 14'h0003; 
        10'b0000110000: data <= 14'h000c; 
        10'b0000110001: data <= 14'h0000; 
        10'b0000110010: data <= 14'h0000; 
        10'b0000110011: data <= 14'h0001; 
        10'b0000110100: data <= 14'h000b; 
        10'b0000110101: data <= 14'h000b; 
        10'b0000110110: data <= 14'h0003; 
        10'b0000110111: data <= 14'h000b; 
        10'b0000111000: data <= 14'h000d; 
        10'b0000111001: data <= 14'h0009; 
        10'b0000111010: data <= 14'h000d; 
        10'b0000111011: data <= 14'h000d; 
        10'b0000111100: data <= 14'h000d; 
        10'b0000111101: data <= 14'h000b; 
        10'b0000111110: data <= 14'h000f; 
        10'b0000111111: data <= 14'h3ffb; 
        10'b0001000000: data <= 14'h3ffb; 
        10'b0001000001: data <= 14'h0003; 
        10'b0001000010: data <= 14'h3ffe; 
        10'b0001000011: data <= 14'h3ff7; 
        10'b0001000100: data <= 14'h3fde; 
        10'b0001000101: data <= 14'h3ff2; 
        10'b0001000110: data <= 14'h3fef; 
        10'b0001000111: data <= 14'h3fe9; 
        10'b0001001000: data <= 14'h3fef; 
        10'b0001001001: data <= 14'h3ffd; 
        10'b0001001010: data <= 14'h0004; 
        10'b0001001011: data <= 14'h000c; 
        10'b0001001100: data <= 14'h0010; 
        10'b0001001101: data <= 14'h0009; 
        10'b0001001110: data <= 14'h000f; 
        10'b0001001111: data <= 14'h0004; 
        10'b0001010000: data <= 14'h0006; 
        10'b0001010001: data <= 14'h000a; 
        10'b0001010010: data <= 14'h0001; 
        10'b0001010011: data <= 14'h0007; 
        10'b0001010100: data <= 14'h000d; 
        10'b0001010101: data <= 14'h000c; 
        10'b0001010110: data <= 14'h0005; 
        10'b0001010111: data <= 14'h0007; 
        10'b0001011000: data <= 14'h0008; 
        10'b0001011001: data <= 14'h0000; 
        10'b0001011010: data <= 14'h000a; 
        10'b0001011011: data <= 14'h3ff7; 
        10'b0001011100: data <= 14'h3ff3; 
        10'b0001011101: data <= 14'h3ff9; 
        10'b0001011110: data <= 14'h3fe3; 
        10'b0001011111: data <= 14'h3fdd; 
        10'b0001100000: data <= 14'h3fc9; 
        10'b0001100001: data <= 14'h3fcb; 
        10'b0001100010: data <= 14'h3fce; 
        10'b0001100011: data <= 14'h3fc3; 
        10'b0001100100: data <= 14'h3fd7; 
        10'b0001100101: data <= 14'h3fec; 
        10'b0001100110: data <= 14'h0003; 
        10'b0001100111: data <= 14'h0007; 
        10'b0001101000: data <= 14'h000c; 
        10'b0001101001: data <= 14'h0011; 
        10'b0001101010: data <= 14'h0005; 
        10'b0001101011: data <= 14'h0005; 
        10'b0001101100: data <= 14'h0011; 
        10'b0001101101: data <= 14'h0010; 
        10'b0001101110: data <= 14'h0005; 
        10'b0001101111: data <= 14'h000a; 
        10'b0001110000: data <= 14'h0010; 
        10'b0001110001: data <= 14'h000b; 
        10'b0001110010: data <= 14'h000c; 
        10'b0001110011: data <= 14'h000c; 
        10'b0001110100: data <= 14'h0007; 
        10'b0001110101: data <= 14'h000e; 
        10'b0001110110: data <= 14'h3ff6; 
        10'b0001110111: data <= 14'h3ffe; 
        10'b0001111000: data <= 14'h3feb; 
        10'b0001111001: data <= 14'h3fef; 
        10'b0001111010: data <= 14'h3fce; 
        10'b0001111011: data <= 14'h3fd1; 
        10'b0001111100: data <= 14'h3fbf; 
        10'b0001111101: data <= 14'h3fca; 
        10'b0001111110: data <= 14'h3fbe; 
        10'b0001111111: data <= 14'h3fc8; 
        10'b0010000000: data <= 14'h3fe5; 
        10'b0010000001: data <= 14'h3fe8; 
        10'b0010000010: data <= 14'h3ff1; 
        10'b0010000011: data <= 14'h000e; 
        10'b0010000100: data <= 14'h0013; 
        10'b0010000101: data <= 14'h0016; 
        10'b0010000110: data <= 14'h0015; 
        10'b0010000111: data <= 14'h001c; 
        10'b0010001000: data <= 14'h0008; 
        10'b0010001001: data <= 14'h0010; 
        10'b0010001010: data <= 14'h0004; 
        10'b0010001011: data <= 14'h0003; 
        10'b0010001100: data <= 14'h0011; 
        10'b0010001101: data <= 14'h0005; 
        10'b0010001110: data <= 14'h000c; 
        10'b0010001111: data <= 14'h0004; 
        10'b0010010000: data <= 14'h000b; 
        10'b0010010001: data <= 14'h0002; 
        10'b0010010010: data <= 14'h0008; 
        10'b0010010011: data <= 14'h3ff7; 
        10'b0010010100: data <= 14'h0003; 
        10'b0010010101: data <= 14'h3ff5; 
        10'b0010010110: data <= 14'h3fdc; 
        10'b0010010111: data <= 14'h3fe8; 
        10'b0010011000: data <= 14'h3fd7; 
        10'b0010011001: data <= 14'h3fcd; 
        10'b0010011010: data <= 14'h3fdc; 
        10'b0010011011: data <= 14'h3fe2; 
        10'b0010011100: data <= 14'h3ffb; 
        10'b0010011101: data <= 14'h0005; 
        10'b0010011110: data <= 14'h3ff9; 
        10'b0010011111: data <= 14'h000c; 
        10'b0010100000: data <= 14'h000f; 
        10'b0010100001: data <= 14'h0014; 
        10'b0010100010: data <= 14'h002e; 
        10'b0010100011: data <= 14'h0034; 
        10'b0010100100: data <= 14'h001c; 
        10'b0010100101: data <= 14'h3ffd; 
        10'b0010100110: data <= 14'h0005; 
        10'b0010100111: data <= 14'h0003; 
        10'b0010101000: data <= 14'h0010; 
        10'b0010101001: data <= 14'h0011; 
        10'b0010101010: data <= 14'h0005; 
        10'b0010101011: data <= 14'h000e; 
        10'b0010101100: data <= 14'h000f; 
        10'b0010101101: data <= 14'h000c; 
        10'b0010101110: data <= 14'h000c; 
        10'b0010101111: data <= 14'h3fff; 
        10'b0010110000: data <= 14'h3ffd; 
        10'b0010110001: data <= 14'h3ff2; 
        10'b0010110010: data <= 14'h3fe3; 
        10'b0010110011: data <= 14'h3fcd; 
        10'b0010110100: data <= 14'h3fb3; 
        10'b0010110101: data <= 14'h3fa5; 
        10'b0010110110: data <= 14'h3fa1; 
        10'b0010110111: data <= 14'h3fae; 
        10'b0010111000: data <= 14'h3fac; 
        10'b0010111001: data <= 14'h3fcf; 
        10'b0010111010: data <= 14'h3fcd; 
        10'b0010111011: data <= 14'h3fe9; 
        10'b0010111100: data <= 14'h3ff1; 
        10'b0010111101: data <= 14'h3fff; 
        10'b0010111110: data <= 14'h0042; 
        10'b0010111111: data <= 14'h0045; 
        10'b0011000000: data <= 14'h001b; 
        10'b0011000001: data <= 14'h0015; 
        10'b0011000010: data <= 14'h000f; 
        10'b0011000011: data <= 14'h0001; 
        10'b0011000100: data <= 14'h0007; 
        10'b0011000101: data <= 14'h0004; 
        10'b0011000110: data <= 14'h0005; 
        10'b0011000111: data <= 14'h0009; 
        10'b0011001000: data <= 14'h0005; 
        10'b0011001001: data <= 14'h000d; 
        10'b0011001010: data <= 14'h3ff8; 
        10'b0011001011: data <= 14'h3fff; 
        10'b0011001100: data <= 14'h3ff7; 
        10'b0011001101: data <= 14'h3fed; 
        10'b0011001110: data <= 14'h3fcf; 
        10'b0011001111: data <= 14'h3fb3; 
        10'b0011010000: data <= 14'h3f9c; 
        10'b0011010001: data <= 14'h3fb9; 
        10'b0011010010: data <= 14'h3fa8; 
        10'b0011010011: data <= 14'h3fa7; 
        10'b0011010100: data <= 14'h3fa5; 
        10'b0011010101: data <= 14'h3fc6; 
        10'b0011010110: data <= 14'h3fc4; 
        10'b0011010111: data <= 14'h3fd6; 
        10'b0011011000: data <= 14'h3fd0; 
        10'b0011011001: data <= 14'h3fea; 
        10'b0011011010: data <= 14'h0029; 
        10'b0011011011: data <= 14'h0037; 
        10'b0011011100: data <= 14'h001d; 
        10'b0011011101: data <= 14'h0011; 
        10'b0011011110: data <= 14'h0010; 
        10'b0011011111: data <= 14'h0009; 
        10'b0011100000: data <= 14'h000f; 
        10'b0011100001: data <= 14'h000d; 
        10'b0011100010: data <= 14'h0011; 
        10'b0011100011: data <= 14'h0003; 
        10'b0011100100: data <= 14'h0005; 
        10'b0011100101: data <= 14'h0007; 
        10'b0011100110: data <= 14'h0005; 
        10'b0011100111: data <= 14'h3ffc; 
        10'b0011101000: data <= 14'h3fdb; 
        10'b0011101001: data <= 14'h3fed; 
        10'b0011101010: data <= 14'h3fe7; 
        10'b0011101011: data <= 14'h3fce; 
        10'b0011101100: data <= 14'h3fb7; 
        10'b0011101101: data <= 14'h3fd2; 
        10'b0011101110: data <= 14'h3f97; 
        10'b0011101111: data <= 14'h3f94; 
        10'b0011110000: data <= 14'h3fac; 
        10'b0011110001: data <= 14'h3fcb; 
        10'b0011110010: data <= 14'h3fd1; 
        10'b0011110011: data <= 14'h3ff1; 
        10'b0011110100: data <= 14'h3fe3; 
        10'b0011110101: data <= 14'h3fe4; 
        10'b0011110110: data <= 14'h0013; 
        10'b0011110111: data <= 14'h001d; 
        10'b0011111000: data <= 14'h0016; 
        10'b0011111001: data <= 14'h0004; 
        10'b0011111010: data <= 14'h0006; 
        10'b0011111011: data <= 14'h000b; 
        10'b0011111100: data <= 14'h0012; 
        10'b0011111101: data <= 14'h000f; 
        10'b0011111110: data <= 14'h000e; 
        10'b0011111111: data <= 14'h0003; 
        10'b0100000000: data <= 14'h3ff7; 
        10'b0100000001: data <= 14'h0000; 
        10'b0100000010: data <= 14'h3fe9; 
        10'b0100000011: data <= 14'h3ff0; 
        10'b0100000100: data <= 14'h3ff5; 
        10'b0100000101: data <= 14'h3ffc; 
        10'b0100000110: data <= 14'h3ff3; 
        10'b0100000111: data <= 14'h3ff1; 
        10'b0100001000: data <= 14'h3ff0; 
        10'b0100001001: data <= 14'h3fd6; 
        10'b0100001010: data <= 14'h3f68; 
        10'b0100001011: data <= 14'h3f8e; 
        10'b0100001100: data <= 14'h3fe4; 
        10'b0100001101: data <= 14'h3fec; 
        10'b0100001110: data <= 14'h3ffa; 
        10'b0100001111: data <= 14'h0003; 
        10'b0100010000: data <= 14'h3ff0; 
        10'b0100010001: data <= 14'h3ff0; 
        10'b0100010010: data <= 14'h0008; 
        10'b0100010011: data <= 14'h0002; 
        10'b0100010100: data <= 14'h3fee; 
        10'b0100010101: data <= 14'h3fed; 
        10'b0100010110: data <= 14'h3ff8; 
        10'b0100010111: data <= 14'h000c; 
        10'b0100011000: data <= 14'h000a; 
        10'b0100011001: data <= 14'h0007; 
        10'b0100011010: data <= 14'h0007; 
        10'b0100011011: data <= 14'h0002; 
        10'b0100011100: data <= 14'h0007; 
        10'b0100011101: data <= 14'h3fec; 
        10'b0100011110: data <= 14'h3fde; 
        10'b0100011111: data <= 14'h3ff0; 
        10'b0100100000: data <= 14'h0005; 
        10'b0100100001: data <= 14'h002b; 
        10'b0100100010: data <= 14'h001a; 
        10'b0100100011: data <= 14'h0014; 
        10'b0100100100: data <= 14'h0017; 
        10'b0100100101: data <= 14'h3fc6; 
        10'b0100100110: data <= 14'h3f60; 
        10'b0100100111: data <= 14'h3fcf; 
        10'b0100101000: data <= 14'h0006; 
        10'b0100101001: data <= 14'h3ff9; 
        10'b0100101010: data <= 14'h3ffb; 
        10'b0100101011: data <= 14'h0006; 
        10'b0100101100: data <= 14'h3fe0; 
        10'b0100101101: data <= 14'h3feb; 
        10'b0100101110: data <= 14'h3ffc; 
        10'b0100101111: data <= 14'h3fdd; 
        10'b0100110000: data <= 14'h3fec; 
        10'b0100110001: data <= 14'h3ff3; 
        10'b0100110010: data <= 14'h000a; 
        10'b0100110011: data <= 14'h0010; 
        10'b0100110100: data <= 14'h000b; 
        10'b0100110101: data <= 14'h000c; 
        10'b0100110110: data <= 14'h000a; 
        10'b0100110111: data <= 14'h3ffa; 
        10'b0100111000: data <= 14'h3ffe; 
        10'b0100111001: data <= 14'h3ff5; 
        10'b0100111010: data <= 14'h3ff4; 
        10'b0100111011: data <= 14'h000a; 
        10'b0100111100: data <= 14'h0021; 
        10'b0100111101: data <= 14'h0037; 
        10'b0100111110: data <= 14'h004c; 
        10'b0100111111: data <= 14'h0030; 
        10'b0101000000: data <= 14'h0037; 
        10'b0101000001: data <= 14'h3fa7; 
        10'b0101000010: data <= 14'h3f87; 
        10'b0101000011: data <= 14'h0010; 
        10'b0101000100: data <= 14'h003e; 
        10'b0101000101: data <= 14'h000b; 
        10'b0101000110: data <= 14'h3ffc; 
        10'b0101000111: data <= 14'h3ff6; 
        10'b0101001000: data <= 14'h3fde; 
        10'b0101001001: data <= 14'h3fe3; 
        10'b0101001010: data <= 14'h3ff1; 
        10'b0101001011: data <= 14'h3fe5; 
        10'b0101001100: data <= 14'h3fe2; 
        10'b0101001101: data <= 14'h3ffe; 
        10'b0101001110: data <= 14'h3fff; 
        10'b0101001111: data <= 14'h0004; 
        10'b0101010000: data <= 14'h000c; 
        10'b0101010001: data <= 14'h000b; 
        10'b0101010010: data <= 14'h0005; 
        10'b0101010011: data <= 14'h0007; 
        10'b0101010100: data <= 14'h3fff; 
        10'b0101010101: data <= 14'h3ff5; 
        10'b0101010110: data <= 14'h0020; 
        10'b0101010111: data <= 14'h0035; 
        10'b0101011000: data <= 14'h0052; 
        10'b0101011001: data <= 14'h0048; 
        10'b0101011010: data <= 14'h0077; 
        10'b0101011011: data <= 14'h0087; 
        10'b0101011100: data <= 14'h0080; 
        10'b0101011101: data <= 14'h3ffe; 
        10'b0101011110: data <= 14'h3fc0; 
        10'b0101011111: data <= 14'h0032; 
        10'b0101100000: data <= 14'h0051; 
        10'b0101100001: data <= 14'h0009; 
        10'b0101100010: data <= 14'h0003; 
        10'b0101100011: data <= 14'h000b; 
        10'b0101100100: data <= 14'h3ffe; 
        10'b0101100101: data <= 14'h0002; 
        10'b0101100110: data <= 14'h3ffc; 
        10'b0101100111: data <= 14'h3fee; 
        10'b0101101000: data <= 14'h3ff0; 
        10'b0101101001: data <= 14'h3ffb; 
        10'b0101101010: data <= 14'h0012; 
        10'b0101101011: data <= 14'h000a; 
        10'b0101101100: data <= 14'h0002; 
        10'b0101101101: data <= 14'h000c; 
        10'b0101101110: data <= 14'h0002; 
        10'b0101101111: data <= 14'h0005; 
        10'b0101110000: data <= 14'h000e; 
        10'b0101110001: data <= 14'h0027; 
        10'b0101110010: data <= 14'h004f; 
        10'b0101110011: data <= 14'h005b; 
        10'b0101110100: data <= 14'h0069; 
        10'b0101110101: data <= 14'h0058; 
        10'b0101110110: data <= 14'h0067; 
        10'b0101110111: data <= 14'h00a7; 
        10'b0101111000: data <= 14'h007f; 
        10'b0101111001: data <= 14'h0002; 
        10'b0101111010: data <= 14'h3fee; 
        10'b0101111011: data <= 14'h003b; 
        10'b0101111100: data <= 14'h003c; 
        10'b0101111101: data <= 14'h0043; 
        10'b0101111110: data <= 14'h002e; 
        10'b0101111111: data <= 14'h0015; 
        10'b0110000000: data <= 14'h002e; 
        10'b0110000001: data <= 14'h0022; 
        10'b0110000010: data <= 14'h0010; 
        10'b0110000011: data <= 14'h3ff7; 
        10'b0110000100: data <= 14'h3ff8; 
        10'b0110000101: data <= 14'h0001; 
        10'b0110000110: data <= 14'h000e; 
        10'b0110000111: data <= 14'h000a; 
        10'b0110001000: data <= 14'h0002; 
        10'b0110001001: data <= 14'h000f; 
        10'b0110001010: data <= 14'h0001; 
        10'b0110001011: data <= 14'h0011; 
        10'b0110001100: data <= 14'h0022; 
        10'b0110001101: data <= 14'h0045; 
        10'b0110001110: data <= 14'h0060; 
        10'b0110001111: data <= 14'h0069; 
        10'b0110010000: data <= 14'h004e; 
        10'b0110010001: data <= 14'h004b; 
        10'b0110010010: data <= 14'h005a; 
        10'b0110010011: data <= 14'h006e; 
        10'b0110010100: data <= 14'h0050; 
        10'b0110010101: data <= 14'h0007; 
        10'b0110010110: data <= 14'h3ff4; 
        10'b0110010111: data <= 14'h0015; 
        10'b0110011000: data <= 14'h0043; 
        10'b0110011001: data <= 14'h006e; 
        10'b0110011010: data <= 14'h004b; 
        10'b0110011011: data <= 14'h0045; 
        10'b0110011100: data <= 14'h0026; 
        10'b0110011101: data <= 14'h001a; 
        10'b0110011110: data <= 14'h0008; 
        10'b0110011111: data <= 14'h0005; 
        10'b0110100000: data <= 14'h3ffd; 
        10'b0110100001: data <= 14'h0005; 
        10'b0110100010: data <= 14'h0009; 
        10'b0110100011: data <= 14'h0004; 
        10'b0110100100: data <= 14'h000c; 
        10'b0110100101: data <= 14'h0011; 
        10'b0110100110: data <= 14'h000b; 
        10'b0110100111: data <= 14'h000e; 
        10'b0110101000: data <= 14'h001f; 
        10'b0110101001: data <= 14'h0023; 
        10'b0110101010: data <= 14'h0037; 
        10'b0110101011: data <= 14'h0032; 
        10'b0110101100: data <= 14'h0051; 
        10'b0110101101: data <= 14'h0046; 
        10'b0110101110: data <= 14'h0030; 
        10'b0110101111: data <= 14'h0023; 
        10'b0110110000: data <= 14'h002a; 
        10'b0110110001: data <= 14'h0008; 
        10'b0110110010: data <= 14'h0021; 
        10'b0110110011: data <= 14'h002f; 
        10'b0110110100: data <= 14'h0061; 
        10'b0110110101: data <= 14'h0056; 
        10'b0110110110: data <= 14'h003d; 
        10'b0110110111: data <= 14'h0024; 
        10'b0110111000: data <= 14'h3ff6; 
        10'b0110111001: data <= 14'h000e; 
        10'b0110111010: data <= 14'h0018; 
        10'b0110111011: data <= 14'h0003; 
        10'b0110111100: data <= 14'h3ff1; 
        10'b0110111101: data <= 14'h0008; 
        10'b0110111110: data <= 14'h0002; 
        10'b0110111111: data <= 14'h0005; 
        10'b0111000000: data <= 14'h0005; 
        10'b0111000001: data <= 14'h0000; 
        10'b0111000010: data <= 14'h0001; 
        10'b0111000011: data <= 14'h3ffe; 
        10'b0111000100: data <= 14'h0008; 
        10'b0111000101: data <= 14'h0015; 
        10'b0111000110: data <= 14'h0022; 
        10'b0111000111: data <= 14'h003b; 
        10'b0111001000: data <= 14'h0056; 
        10'b0111001001: data <= 14'h003d; 
        10'b0111001010: data <= 14'h0010; 
        10'b0111001011: data <= 14'h3ffe; 
        10'b0111001100: data <= 14'h0011; 
        10'b0111001101: data <= 14'h0015; 
        10'b0111001110: data <= 14'h004f; 
        10'b0111001111: data <= 14'h006d; 
        10'b0111010000: data <= 14'h0070; 
        10'b0111010001: data <= 14'h005d; 
        10'b0111010010: data <= 14'h003f; 
        10'b0111010011: data <= 14'h0008; 
        10'b0111010100: data <= 14'h001a; 
        10'b0111010101: data <= 14'h0026; 
        10'b0111010110: data <= 14'h0009; 
        10'b0111010111: data <= 14'h3ffa; 
        10'b0111011000: data <= 14'h3ffe; 
        10'b0111011001: data <= 14'h0004; 
        10'b0111011010: data <= 14'h0007; 
        10'b0111011011: data <= 14'h0007; 
        10'b0111011100: data <= 14'h0006; 
        10'b0111011101: data <= 14'h0006; 
        10'b0111011110: data <= 14'h000d; 
        10'b0111011111: data <= 14'h0000; 
        10'b0111100000: data <= 14'h3ff7; 
        10'b0111100001: data <= 14'h3fed; 
        10'b0111100010: data <= 14'h000b; 
        10'b0111100011: data <= 14'h002f; 
        10'b0111100100: data <= 14'h005a; 
        10'b0111100101: data <= 14'h004e; 
        10'b0111100110: data <= 14'h001c; 
        10'b0111100111: data <= 14'h0016; 
        10'b0111101000: data <= 14'h0020; 
        10'b0111101001: data <= 14'h004d; 
        10'b0111101010: data <= 14'h0080; 
        10'b0111101011: data <= 14'h0065; 
        10'b0111101100: data <= 14'h0055; 
        10'b0111101101: data <= 14'h001a; 
        10'b0111101110: data <= 14'h0004; 
        10'b0111101111: data <= 14'h3fe4; 
        10'b0111110000: data <= 14'h0008; 
        10'b0111110001: data <= 14'h0003; 
        10'b0111110010: data <= 14'h3fef; 
        10'b0111110011: data <= 14'h3ff9; 
        10'b0111110100: data <= 14'h3ff5; 
        10'b0111110101: data <= 14'h3ffa; 
        10'b0111110110: data <= 14'h000b; 
        10'b0111110111: data <= 14'h000e; 
        10'b0111111000: data <= 14'h0007; 
        10'b0111111001: data <= 14'h000b; 
        10'b0111111010: data <= 14'h0009; 
        10'b0111111011: data <= 14'h0001; 
        10'b0111111100: data <= 14'h3ff5; 
        10'b0111111101: data <= 14'h3fe9; 
        10'b0111111110: data <= 14'h3fe5; 
        10'b0111111111: data <= 14'h3fff; 
        10'b1000000000: data <= 14'h0017; 
        10'b1000000001: data <= 14'h0005; 
        10'b1000000010: data <= 14'h3fed; 
        10'b1000000011: data <= 14'h3ff5; 
        10'b1000000100: data <= 14'h001e; 
        10'b1000000101: data <= 14'h0021; 
        10'b1000000110: data <= 14'h0038; 
        10'b1000000111: data <= 14'h0030; 
        10'b1000001000: data <= 14'h0019; 
        10'b1000001001: data <= 14'h3fd9; 
        10'b1000001010: data <= 14'h3fdb; 
        10'b1000001011: data <= 14'h3fca; 
        10'b1000001100: data <= 14'h3fe0; 
        10'b1000001101: data <= 14'h3fdf; 
        10'b1000001110: data <= 14'h3fd4; 
        10'b1000001111: data <= 14'h3fde; 
        10'b1000010000: data <= 14'h3ff7; 
        10'b1000010001: data <= 14'h3ffb; 
        10'b1000010010: data <= 14'h0004; 
        10'b1000010011: data <= 14'h0001; 
        10'b1000010100: data <= 14'h0007; 
        10'b1000010101: data <= 14'h000d; 
        10'b1000010110: data <= 14'h0005; 
        10'b1000010111: data <= 14'h0003; 
        10'b1000011000: data <= 14'h3fe7; 
        10'b1000011001: data <= 14'h3fe1; 
        10'b1000011010: data <= 14'h3fd7; 
        10'b1000011011: data <= 14'h3fc3; 
        10'b1000011100: data <= 14'h3fbb; 
        10'b1000011101: data <= 14'h3fb7; 
        10'b1000011110: data <= 14'h3fa9; 
        10'b1000011111: data <= 14'h3fad; 
        10'b1000100000: data <= 14'h3fb7; 
        10'b1000100001: data <= 14'h3fd5; 
        10'b1000100010: data <= 14'h3ff3; 
        10'b1000100011: data <= 14'h000b; 
        10'b1000100100: data <= 14'h3fdf; 
        10'b1000100101: data <= 14'h3fe3; 
        10'b1000100110: data <= 14'h3fdd; 
        10'b1000100111: data <= 14'h3fcf; 
        10'b1000101000: data <= 14'h3fc9; 
        10'b1000101001: data <= 14'h3fce; 
        10'b1000101010: data <= 14'h3fcd; 
        10'b1000101011: data <= 14'h3fdd; 
        10'b1000101100: data <= 14'h3ff7; 
        10'b1000101101: data <= 14'h0007; 
        10'b1000101110: data <= 14'h000c; 
        10'b1000101111: data <= 14'h000b; 
        10'b1000110000: data <= 14'h0012; 
        10'b1000110001: data <= 14'h0011; 
        10'b1000110010: data <= 14'h0005; 
        10'b1000110011: data <= 14'h0003; 
        10'b1000110100: data <= 14'h3fec; 
        10'b1000110101: data <= 14'h3fde; 
        10'b1000110110: data <= 14'h3fce; 
        10'b1000110111: data <= 14'h3faf; 
        10'b1000111000: data <= 14'h3f9f; 
        10'b1000111001: data <= 14'h3f9a; 
        10'b1000111010: data <= 14'h3f98; 
        10'b1000111011: data <= 14'h3fb4; 
        10'b1000111100: data <= 14'h3fc2; 
        10'b1000111101: data <= 14'h3fbb; 
        10'b1000111110: data <= 14'h3fd5; 
        10'b1000111111: data <= 14'h3fe9; 
        10'b1001000000: data <= 14'h3ff8; 
        10'b1001000001: data <= 14'h3ffc; 
        10'b1001000010: data <= 14'h3fee; 
        10'b1001000011: data <= 14'h3fd9; 
        10'b1001000100: data <= 14'h3fe6; 
        10'b1001000101: data <= 14'h3fe2; 
        10'b1001000110: data <= 14'h3fdc; 
        10'b1001000111: data <= 14'h3fee; 
        10'b1001001000: data <= 14'h3fee; 
        10'b1001001001: data <= 14'h0001; 
        10'b1001001010: data <= 14'h0004; 
        10'b1001001011: data <= 14'h000c; 
        10'b1001001100: data <= 14'h0003; 
        10'b1001001101: data <= 14'h0005; 
        10'b1001001110: data <= 14'h0001; 
        10'b1001001111: data <= 14'h0002; 
        10'b1001010000: data <= 14'h0000; 
        10'b1001010001: data <= 14'h3fec; 
        10'b1001010010: data <= 14'h3fcf; 
        10'b1001010011: data <= 14'h3fbb; 
        10'b1001010100: data <= 14'h3fc2; 
        10'b1001010101: data <= 14'h3fb9; 
        10'b1001010110: data <= 14'h3fc3; 
        10'b1001010111: data <= 14'h3fd2; 
        10'b1001011000: data <= 14'h3fda; 
        10'b1001011001: data <= 14'h3fdd; 
        10'b1001011010: data <= 14'h3fd8; 
        10'b1001011011: data <= 14'h3fed; 
        10'b1001011100: data <= 14'h3fe7; 
        10'b1001011101: data <= 14'h0004; 
        10'b1001011110: data <= 14'h3ff9; 
        10'b1001011111: data <= 14'h0001; 
        10'b1001100000: data <= 14'h3ffd; 
        10'b1001100001: data <= 14'h3fe8; 
        10'b1001100010: data <= 14'h3fec; 
        10'b1001100011: data <= 14'h3ffc; 
        10'b1001100100: data <= 14'h3fff; 
        10'b1001100101: data <= 14'h0007; 
        10'b1001100110: data <= 14'h000a; 
        10'b1001100111: data <= 14'h000a; 
        10'b1001101000: data <= 14'h0009; 
        10'b1001101001: data <= 14'h000a; 
        10'b1001101010: data <= 14'h0004; 
        10'b1001101011: data <= 14'h000b; 
        10'b1001101100: data <= 14'h3ffd; 
        10'b1001101101: data <= 14'h3ff6; 
        10'b1001101110: data <= 14'h3fec; 
        10'b1001101111: data <= 14'h3fde; 
        10'b1001110000: data <= 14'h3fd3; 
        10'b1001110001: data <= 14'h3fe5; 
        10'b1001110010: data <= 14'h3fe4; 
        10'b1001110011: data <= 14'h3fec; 
        10'b1001110100: data <= 14'h3feb; 
        10'b1001110101: data <= 14'h3fee; 
        10'b1001110110: data <= 14'h3fea; 
        10'b1001110111: data <= 14'h3ff2; 
        10'b1001111000: data <= 14'h3ff3; 
        10'b1001111001: data <= 14'h0005; 
        10'b1001111010: data <= 14'h0014; 
        10'b1001111011: data <= 14'h0021; 
        10'b1001111100: data <= 14'h0019; 
        10'b1001111101: data <= 14'h0010; 
        10'b1001111110: data <= 14'h3ff5; 
        10'b1001111111: data <= 14'h3ff5; 
        10'b1010000000: data <= 14'h0000; 
        10'b1010000001: data <= 14'h0007; 
        10'b1010000010: data <= 14'h0001; 
        10'b1010000011: data <= 14'h0006; 
        10'b1010000100: data <= 14'h0006; 
        10'b1010000101: data <= 14'h0000; 
        10'b1010000110: data <= 14'h0005; 
        10'b1010000111: data <= 14'h000a; 
        10'b1010001000: data <= 14'h0006; 
        10'b1010001001: data <= 14'h0007; 
        10'b1010001010: data <= 14'h3ff5; 
        10'b1010001011: data <= 14'h3ff4; 
        10'b1010001100: data <= 14'h3ff0; 
        10'b1010001101: data <= 14'h0008; 
        10'b1010001110: data <= 14'h3fef; 
        10'b1010001111: data <= 14'h0003; 
        10'b1010010000: data <= 14'h3fee; 
        10'b1010010001: data <= 14'h3ff2; 
        10'b1010010010: data <= 14'h3ff2; 
        10'b1010010011: data <= 14'h3fff; 
        10'b1010010100: data <= 14'h0005; 
        10'b1010010101: data <= 14'h000c; 
        10'b1010010110: data <= 14'h0026; 
        10'b1010010111: data <= 14'h0025; 
        10'b1010011000: data <= 14'h001f; 
        10'b1010011001: data <= 14'h000e; 
        10'b1010011010: data <= 14'h3ffb; 
        10'b1010011011: data <= 14'h0004; 
        10'b1010011100: data <= 14'h0008; 
        10'b1010011101: data <= 14'h000b; 
        10'b1010011110: data <= 14'h0004; 
        10'b1010011111: data <= 14'h000e; 
        10'b1010100000: data <= 14'h000b; 
        10'b1010100001: data <= 14'h000f; 
        10'b1010100010: data <= 14'h0007; 
        10'b1010100011: data <= 14'h000c; 
        10'b1010100100: data <= 14'h0003; 
        10'b1010100101: data <= 14'h0009; 
        10'b1010100110: data <= 14'h0004; 
        10'b1010100111: data <= 14'h3fef; 
        10'b1010101000: data <= 14'h3fee; 
        10'b1010101001: data <= 14'h3ffa; 
        10'b1010101010: data <= 14'h3fed; 
        10'b1010101011: data <= 14'h3ffd; 
        10'b1010101100: data <= 14'h3ff3; 
        10'b1010101101: data <= 14'h3ff4; 
        10'b1010101110: data <= 14'h3fe9; 
        10'b1010101111: data <= 14'h3fe6; 
        10'b1010110000: data <= 14'h3ff5; 
        10'b1010110001: data <= 14'h3ffa; 
        10'b1010110010: data <= 14'h0002; 
        10'b1010110011: data <= 14'h0014; 
        10'b1010110100: data <= 14'h000e; 
        10'b1010110101: data <= 14'h3ffa; 
        10'b1010110110: data <= 14'h3ffe; 
        10'b1010110111: data <= 14'h0008; 
        10'b1010111000: data <= 14'h000d; 
        10'b1010111001: data <= 14'h0002; 
        10'b1010111010: data <= 14'h0003; 
        10'b1010111011: data <= 14'h000b; 
        10'b1010111100: data <= 14'h0010; 
        10'b1010111101: data <= 14'h0010; 
        10'b1010111110: data <= 14'h000e; 
        10'b1010111111: data <= 14'h0003; 
        10'b1011000000: data <= 14'h000e; 
        10'b1011000001: data <= 14'h0001; 
        10'b1011000010: data <= 14'h3ff6; 
        10'b1011000011: data <= 14'h3fef; 
        10'b1011000100: data <= 14'h3fe7; 
        10'b1011000101: data <= 14'h3fe6; 
        10'b1011000110: data <= 14'h3fd5; 
        10'b1011000111: data <= 14'h3fcf; 
        10'b1011001000: data <= 14'h3fd2; 
        10'b1011001001: data <= 14'h3fd2; 
        10'b1011001010: data <= 14'h3fd9; 
        10'b1011001011: data <= 14'h3fd7; 
        10'b1011001100: data <= 14'h3fcb; 
        10'b1011001101: data <= 14'h3fc3; 
        10'b1011001110: data <= 14'h3fca; 
        10'b1011001111: data <= 14'h3fe2; 
        10'b1011010000: data <= 14'h3fe5; 
        10'b1011010001: data <= 14'h3ff6; 
        10'b1011010010: data <= 14'h0001; 
        10'b1011010011: data <= 14'h000a; 
        10'b1011010100: data <= 14'h0001; 
        10'b1011010101: data <= 14'h000f; 
        10'b1011010110: data <= 14'h0006; 
        10'b1011010111: data <= 14'h0005; 
        10'b1011011000: data <= 14'h0007; 
        10'b1011011001: data <= 14'h000b; 
        10'b1011011010: data <= 14'h0002; 
        10'b1011011011: data <= 14'h0007; 
        10'b1011011100: data <= 14'h3fff; 
        10'b1011011101: data <= 14'h3ffe; 
        10'b1011011110: data <= 14'h0004; 
        10'b1011011111: data <= 14'h0003; 
        10'b1011100000: data <= 14'h3ffd; 
        10'b1011100001: data <= 14'h3ff1; 
        10'b1011100010: data <= 14'h3fdc; 
        10'b1011100011: data <= 14'h3fe0; 
        10'b1011100100: data <= 14'h3fdc; 
        10'b1011100101: data <= 14'h3fcf; 
        10'b1011100110: data <= 14'h3fca; 
        10'b1011100111: data <= 14'h3fd6; 
        10'b1011101000: data <= 14'h3fd0; 
        10'b1011101001: data <= 14'h3fd7; 
        10'b1011101010: data <= 14'h3fdf; 
        10'b1011101011: data <= 14'h3fec; 
        10'b1011101100: data <= 14'h3ff9; 
        10'b1011101101: data <= 14'h000b; 
        10'b1011101110: data <= 14'h000b; 
        10'b1011101111: data <= 14'h0001; 
        10'b1011110000: data <= 14'h0007; 
        10'b1011110001: data <= 14'h0001; 
        10'b1011110010: data <= 14'h0011; 
        10'b1011110011: data <= 14'h0008; 
        10'b1011110100: data <= 14'h000a; 
        10'b1011110101: data <= 14'h0002; 
        10'b1011110110: data <= 14'h0002; 
        10'b1011110111: data <= 14'h0011; 
        10'b1011111000: data <= 14'h0006; 
        10'b1011111001: data <= 14'h000e; 
        10'b1011111010: data <= 14'h0006; 
        10'b1011111011: data <= 14'h0011; 
        10'b1011111100: data <= 14'h0000; 
        10'b1011111101: data <= 14'h0007; 
        10'b1011111110: data <= 14'h0004; 
        10'b1011111111: data <= 14'h3ffe; 
        10'b1100000000: data <= 14'h3ffe; 
        10'b1100000001: data <= 14'h0001; 
        10'b1100000010: data <= 14'h3ff9; 
        10'b1100000011: data <= 14'h000d; 
        10'b1100000100: data <= 14'h3ffd; 
        10'b1100000101: data <= 14'h3ffc; 
        10'b1100000110: data <= 14'h3fff; 
        10'b1100000111: data <= 14'h0007; 
        10'b1100001000: data <= 14'h0005; 
        10'b1100001001: data <= 14'h0005; 
        10'b1100001010: data <= 14'h0006; 
        10'b1100001011: data <= 14'h000a; 
        10'b1100001100: data <= 14'h0009; 
        10'b1100001101: data <= 14'h000c; 
        10'b1100001110: data <= 14'h0009; 
        10'b1100001111: data <= 14'h0006; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 9) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 15'h0000; 
        10'b0000000001: data <= 15'h0005; 
        10'b0000000010: data <= 15'h001e; 
        10'b0000000011: data <= 15'h001e; 
        10'b0000000100: data <= 15'h0001; 
        10'b0000000101: data <= 15'h0001; 
        10'b0000000110: data <= 15'h0018; 
        10'b0000000111: data <= 15'h0006; 
        10'b0000001000: data <= 15'h0002; 
        10'b0000001001: data <= 15'h0004; 
        10'b0000001010: data <= 15'h0001; 
        10'b0000001011: data <= 15'h0016; 
        10'b0000001100: data <= 15'h001d; 
        10'b0000001101: data <= 15'h0010; 
        10'b0000001110: data <= 15'h0015; 
        10'b0000001111: data <= 15'h0002; 
        10'b0000010000: data <= 15'h0014; 
        10'b0000010001: data <= 15'h001b; 
        10'b0000010010: data <= 15'h0006; 
        10'b0000010011: data <= 15'h0016; 
        10'b0000010100: data <= 15'h0002; 
        10'b0000010101: data <= 15'h000d; 
        10'b0000010110: data <= 15'h001d; 
        10'b0000010111: data <= 15'h0003; 
        10'b0000011000: data <= 15'h001d; 
        10'b0000011001: data <= 15'h0005; 
        10'b0000011010: data <= 15'h0020; 
        10'b0000011011: data <= 15'h000d; 
        10'b0000011100: data <= 15'h0008; 
        10'b0000011101: data <= 15'h000f; 
        10'b0000011110: data <= 15'h0000; 
        10'b0000011111: data <= 15'h0003; 
        10'b0000100000: data <= 15'h000f; 
        10'b0000100001: data <= 15'h0023; 
        10'b0000100010: data <= 15'h0007; 
        10'b0000100011: data <= 15'h7ffa; 
        10'b0000100100: data <= 15'h0014; 
        10'b0000100101: data <= 15'h0001; 
        10'b0000100110: data <= 15'h000d; 
        10'b0000100111: data <= 15'h7ff6; 
        10'b0000101000: data <= 15'h0009; 
        10'b0000101001: data <= 15'h7ff2; 
        10'b0000101010: data <= 15'h0001; 
        10'b0000101011: data <= 15'h0013; 
        10'b0000101100: data <= 15'h0017; 
        10'b0000101101: data <= 15'h0007; 
        10'b0000101110: data <= 15'h0000; 
        10'b0000101111: data <= 15'h0006; 
        10'b0000110000: data <= 15'h0018; 
        10'b0000110001: data <= 15'h7fff; 
        10'b0000110010: data <= 15'h7fff; 
        10'b0000110011: data <= 15'h0002; 
        10'b0000110100: data <= 15'h0016; 
        10'b0000110101: data <= 15'h0017; 
        10'b0000110110: data <= 15'h0005; 
        10'b0000110111: data <= 15'h0017; 
        10'b0000111000: data <= 15'h001a; 
        10'b0000111001: data <= 15'h0011; 
        10'b0000111010: data <= 15'h001a; 
        10'b0000111011: data <= 15'h001b; 
        10'b0000111100: data <= 15'h0019; 
        10'b0000111101: data <= 15'h0016; 
        10'b0000111110: data <= 15'h001e; 
        10'b0000111111: data <= 15'h7ff6; 
        10'b0001000000: data <= 15'h7ff6; 
        10'b0001000001: data <= 15'h0005; 
        10'b0001000010: data <= 15'h7ffd; 
        10'b0001000011: data <= 15'h7fee; 
        10'b0001000100: data <= 15'h7fbc; 
        10'b0001000101: data <= 15'h7fe4; 
        10'b0001000110: data <= 15'h7fdf; 
        10'b0001000111: data <= 15'h7fd1; 
        10'b0001001000: data <= 15'h7fde; 
        10'b0001001001: data <= 15'h7ff9; 
        10'b0001001010: data <= 15'h0009; 
        10'b0001001011: data <= 15'h0018; 
        10'b0001001100: data <= 15'h001f; 
        10'b0001001101: data <= 15'h0012; 
        10'b0001001110: data <= 15'h001d; 
        10'b0001001111: data <= 15'h0008; 
        10'b0001010000: data <= 15'h000b; 
        10'b0001010001: data <= 15'h0014; 
        10'b0001010010: data <= 15'h0001; 
        10'b0001010011: data <= 15'h000e; 
        10'b0001010100: data <= 15'h001a; 
        10'b0001010101: data <= 15'h0018; 
        10'b0001010110: data <= 15'h0009; 
        10'b0001010111: data <= 15'h000f; 
        10'b0001011000: data <= 15'h0010; 
        10'b0001011001: data <= 15'h0000; 
        10'b0001011010: data <= 15'h0014; 
        10'b0001011011: data <= 15'h7fee; 
        10'b0001011100: data <= 15'h7fe6; 
        10'b0001011101: data <= 15'h7ff2; 
        10'b0001011110: data <= 15'h7fc5; 
        10'b0001011111: data <= 15'h7fbb; 
        10'b0001100000: data <= 15'h7f91; 
        10'b0001100001: data <= 15'h7f96; 
        10'b0001100010: data <= 15'h7f9b; 
        10'b0001100011: data <= 15'h7f86; 
        10'b0001100100: data <= 15'h7fae; 
        10'b0001100101: data <= 15'h7fd7; 
        10'b0001100110: data <= 15'h0006; 
        10'b0001100111: data <= 15'h000d; 
        10'b0001101000: data <= 15'h0018; 
        10'b0001101001: data <= 15'h0023; 
        10'b0001101010: data <= 15'h0009; 
        10'b0001101011: data <= 15'h0009; 
        10'b0001101100: data <= 15'h0022; 
        10'b0001101101: data <= 15'h0021; 
        10'b0001101110: data <= 15'h000a; 
        10'b0001101111: data <= 15'h0013; 
        10'b0001110000: data <= 15'h0021; 
        10'b0001110001: data <= 15'h0016; 
        10'b0001110010: data <= 15'h0019; 
        10'b0001110011: data <= 15'h0018; 
        10'b0001110100: data <= 15'h000e; 
        10'b0001110101: data <= 15'h001b; 
        10'b0001110110: data <= 15'h7fec; 
        10'b0001110111: data <= 15'h7ffb; 
        10'b0001111000: data <= 15'h7fd7; 
        10'b0001111001: data <= 15'h7fdd; 
        10'b0001111010: data <= 15'h7f9d; 
        10'b0001111011: data <= 15'h7fa1; 
        10'b0001111100: data <= 15'h7f7f; 
        10'b0001111101: data <= 15'h7f95; 
        10'b0001111110: data <= 15'h7f7c; 
        10'b0001111111: data <= 15'h7f8f; 
        10'b0010000000: data <= 15'h7fc9; 
        10'b0010000001: data <= 15'h7fcf; 
        10'b0010000010: data <= 15'h7fe3; 
        10'b0010000011: data <= 15'h001c; 
        10'b0010000100: data <= 15'h0027; 
        10'b0010000101: data <= 15'h002c; 
        10'b0010000110: data <= 15'h002a; 
        10'b0010000111: data <= 15'h0038; 
        10'b0010001000: data <= 15'h000f; 
        10'b0010001001: data <= 15'h001f; 
        10'b0010001010: data <= 15'h0008; 
        10'b0010001011: data <= 15'h0005; 
        10'b0010001100: data <= 15'h0022; 
        10'b0010001101: data <= 15'h0009; 
        10'b0010001110: data <= 15'h0018; 
        10'b0010001111: data <= 15'h0008; 
        10'b0010010000: data <= 15'h0016; 
        10'b0010010001: data <= 15'h0004; 
        10'b0010010010: data <= 15'h000f; 
        10'b0010010011: data <= 15'h7fed; 
        10'b0010010100: data <= 15'h0005; 
        10'b0010010101: data <= 15'h7fea; 
        10'b0010010110: data <= 15'h7fb7; 
        10'b0010010111: data <= 15'h7fd0; 
        10'b0010011000: data <= 15'h7fad; 
        10'b0010011001: data <= 15'h7f99; 
        10'b0010011010: data <= 15'h7fb8; 
        10'b0010011011: data <= 15'h7fc5; 
        10'b0010011100: data <= 15'h7ff6; 
        10'b0010011101: data <= 15'h0009; 
        10'b0010011110: data <= 15'h7ff2; 
        10'b0010011111: data <= 15'h0018; 
        10'b0010100000: data <= 15'h001d; 
        10'b0010100001: data <= 15'h0028; 
        10'b0010100010: data <= 15'h005c; 
        10'b0010100011: data <= 15'h0068; 
        10'b0010100100: data <= 15'h0039; 
        10'b0010100101: data <= 15'h7ffa; 
        10'b0010100110: data <= 15'h0009; 
        10'b0010100111: data <= 15'h0006; 
        10'b0010101000: data <= 15'h001f; 
        10'b0010101001: data <= 15'h0022; 
        10'b0010101010: data <= 15'h000a; 
        10'b0010101011: data <= 15'h001b; 
        10'b0010101100: data <= 15'h001d; 
        10'b0010101101: data <= 15'h0018; 
        10'b0010101110: data <= 15'h0018; 
        10'b0010101111: data <= 15'h7ffe; 
        10'b0010110000: data <= 15'h7ffb; 
        10'b0010110001: data <= 15'h7fe3; 
        10'b0010110010: data <= 15'h7fc6; 
        10'b0010110011: data <= 15'h7f9b; 
        10'b0010110100: data <= 15'h7f66; 
        10'b0010110101: data <= 15'h7f4a; 
        10'b0010110110: data <= 15'h7f42; 
        10'b0010110111: data <= 15'h7f5b; 
        10'b0010111000: data <= 15'h7f57; 
        10'b0010111001: data <= 15'h7f9d; 
        10'b0010111010: data <= 15'h7f9a; 
        10'b0010111011: data <= 15'h7fd2; 
        10'b0010111100: data <= 15'h7fe2; 
        10'b0010111101: data <= 15'h7ffe; 
        10'b0010111110: data <= 15'h0084; 
        10'b0010111111: data <= 15'h008b; 
        10'b0011000000: data <= 15'h0035; 
        10'b0011000001: data <= 15'h002a; 
        10'b0011000010: data <= 15'h001e; 
        10'b0011000011: data <= 15'h0001; 
        10'b0011000100: data <= 15'h000f; 
        10'b0011000101: data <= 15'h0008; 
        10'b0011000110: data <= 15'h000b; 
        10'b0011000111: data <= 15'h0013; 
        10'b0011001000: data <= 15'h000b; 
        10'b0011001001: data <= 15'h0019; 
        10'b0011001010: data <= 15'h7ff0; 
        10'b0011001011: data <= 15'h7ffd; 
        10'b0011001100: data <= 15'h7fef; 
        10'b0011001101: data <= 15'h7fd9; 
        10'b0011001110: data <= 15'h7f9d; 
        10'b0011001111: data <= 15'h7f66; 
        10'b0011010000: data <= 15'h7f38; 
        10'b0011010001: data <= 15'h7f73; 
        10'b0011010010: data <= 15'h7f50; 
        10'b0011010011: data <= 15'h7f4e; 
        10'b0011010100: data <= 15'h7f49; 
        10'b0011010101: data <= 15'h7f8c; 
        10'b0011010110: data <= 15'h7f89; 
        10'b0011010111: data <= 15'h7fad; 
        10'b0011011000: data <= 15'h7fa0; 
        10'b0011011001: data <= 15'h7fd4; 
        10'b0011011010: data <= 15'h0052; 
        10'b0011011011: data <= 15'h006e; 
        10'b0011011100: data <= 15'h003b; 
        10'b0011011101: data <= 15'h0021; 
        10'b0011011110: data <= 15'h001f; 
        10'b0011011111: data <= 15'h0012; 
        10'b0011100000: data <= 15'h001e; 
        10'b0011100001: data <= 15'h0019; 
        10'b0011100010: data <= 15'h0021; 
        10'b0011100011: data <= 15'h0006; 
        10'b0011100100: data <= 15'h000a; 
        10'b0011100101: data <= 15'h000e; 
        10'b0011100110: data <= 15'h0009; 
        10'b0011100111: data <= 15'h7ff8; 
        10'b0011101000: data <= 15'h7fb6; 
        10'b0011101001: data <= 15'h7fda; 
        10'b0011101010: data <= 15'h7fcf; 
        10'b0011101011: data <= 15'h7f9d; 
        10'b0011101100: data <= 15'h7f6f; 
        10'b0011101101: data <= 15'h7fa3; 
        10'b0011101110: data <= 15'h7f2d; 
        10'b0011101111: data <= 15'h7f28; 
        10'b0011110000: data <= 15'h7f58; 
        10'b0011110001: data <= 15'h7f97; 
        10'b0011110010: data <= 15'h7fa1; 
        10'b0011110011: data <= 15'h7fe2; 
        10'b0011110100: data <= 15'h7fc6; 
        10'b0011110101: data <= 15'h7fc7; 
        10'b0011110110: data <= 15'h0026; 
        10'b0011110111: data <= 15'h003a; 
        10'b0011111000: data <= 15'h002c; 
        10'b0011111001: data <= 15'h0009; 
        10'b0011111010: data <= 15'h000c; 
        10'b0011111011: data <= 15'h0016; 
        10'b0011111100: data <= 15'h0024; 
        10'b0011111101: data <= 15'h001e; 
        10'b0011111110: data <= 15'h001c; 
        10'b0011111111: data <= 15'h0006; 
        10'b0100000000: data <= 15'h7fed; 
        10'b0100000001: data <= 15'h0001; 
        10'b0100000010: data <= 15'h7fd2; 
        10'b0100000011: data <= 15'h7fdf; 
        10'b0100000100: data <= 15'h7feb; 
        10'b0100000101: data <= 15'h7ff9; 
        10'b0100000110: data <= 15'h7fe7; 
        10'b0100000111: data <= 15'h7fe1; 
        10'b0100001000: data <= 15'h7fe0; 
        10'b0100001001: data <= 15'h7fac; 
        10'b0100001010: data <= 15'h7ed0; 
        10'b0100001011: data <= 15'h7f1d; 
        10'b0100001100: data <= 15'h7fc9; 
        10'b0100001101: data <= 15'h7fd7; 
        10'b0100001110: data <= 15'h7ff3; 
        10'b0100001111: data <= 15'h0007; 
        10'b0100010000: data <= 15'h7fe0; 
        10'b0100010001: data <= 15'h7fe1; 
        10'b0100010010: data <= 15'h0010; 
        10'b0100010011: data <= 15'h0004; 
        10'b0100010100: data <= 15'h7fdc; 
        10'b0100010101: data <= 15'h7fda; 
        10'b0100010110: data <= 15'h7ff0; 
        10'b0100010111: data <= 15'h0018; 
        10'b0100011000: data <= 15'h0013; 
        10'b0100011001: data <= 15'h000d; 
        10'b0100011010: data <= 15'h000e; 
        10'b0100011011: data <= 15'h0004; 
        10'b0100011100: data <= 15'h000e; 
        10'b0100011101: data <= 15'h7fd7; 
        10'b0100011110: data <= 15'h7fbc; 
        10'b0100011111: data <= 15'h7fdf; 
        10'b0100100000: data <= 15'h000a; 
        10'b0100100001: data <= 15'h0057; 
        10'b0100100010: data <= 15'h0034; 
        10'b0100100011: data <= 15'h0027; 
        10'b0100100100: data <= 15'h002f; 
        10'b0100100101: data <= 15'h7f8c; 
        10'b0100100110: data <= 15'h7ebf; 
        10'b0100100111: data <= 15'h7f9e; 
        10'b0100101000: data <= 15'h000b; 
        10'b0100101001: data <= 15'h7ff2; 
        10'b0100101010: data <= 15'h7ff5; 
        10'b0100101011: data <= 15'h000b; 
        10'b0100101100: data <= 15'h7fc0; 
        10'b0100101101: data <= 15'h7fd6; 
        10'b0100101110: data <= 15'h7ff8; 
        10'b0100101111: data <= 15'h7fba; 
        10'b0100110000: data <= 15'h7fd9; 
        10'b0100110001: data <= 15'h7fe7; 
        10'b0100110010: data <= 15'h0014; 
        10'b0100110011: data <= 15'h0021; 
        10'b0100110100: data <= 15'h0016; 
        10'b0100110101: data <= 15'h0017; 
        10'b0100110110: data <= 15'h0014; 
        10'b0100110111: data <= 15'h7ff4; 
        10'b0100111000: data <= 15'h7ffb; 
        10'b0100111001: data <= 15'h7fe9; 
        10'b0100111010: data <= 15'h7fe8; 
        10'b0100111011: data <= 15'h0014; 
        10'b0100111100: data <= 15'h0041; 
        10'b0100111101: data <= 15'h006e; 
        10'b0100111110: data <= 15'h0098; 
        10'b0100111111: data <= 15'h0061; 
        10'b0101000000: data <= 15'h006d; 
        10'b0101000001: data <= 15'h7f4e; 
        10'b0101000010: data <= 15'h7f0f; 
        10'b0101000011: data <= 15'h001f; 
        10'b0101000100: data <= 15'h007d; 
        10'b0101000101: data <= 15'h0015; 
        10'b0101000110: data <= 15'h7ff9; 
        10'b0101000111: data <= 15'h7fec; 
        10'b0101001000: data <= 15'h7fbc; 
        10'b0101001001: data <= 15'h7fc6; 
        10'b0101001010: data <= 15'h7fe2; 
        10'b0101001011: data <= 15'h7fca; 
        10'b0101001100: data <= 15'h7fc4; 
        10'b0101001101: data <= 15'h7ffd; 
        10'b0101001110: data <= 15'h7ffe; 
        10'b0101001111: data <= 15'h0008; 
        10'b0101010000: data <= 15'h0019; 
        10'b0101010001: data <= 15'h0016; 
        10'b0101010010: data <= 15'h000a; 
        10'b0101010011: data <= 15'h000f; 
        10'b0101010100: data <= 15'h7ffe; 
        10'b0101010101: data <= 15'h7fea; 
        10'b0101010110: data <= 15'h0040; 
        10'b0101010111: data <= 15'h006a; 
        10'b0101011000: data <= 15'h00a4; 
        10'b0101011001: data <= 15'h0090; 
        10'b0101011010: data <= 15'h00ef; 
        10'b0101011011: data <= 15'h010f; 
        10'b0101011100: data <= 15'h0100; 
        10'b0101011101: data <= 15'h7ffc; 
        10'b0101011110: data <= 15'h7f81; 
        10'b0101011111: data <= 15'h0064; 
        10'b0101100000: data <= 15'h00a3; 
        10'b0101100001: data <= 15'h0012; 
        10'b0101100010: data <= 15'h0007; 
        10'b0101100011: data <= 15'h0016; 
        10'b0101100100: data <= 15'h7ffc; 
        10'b0101100101: data <= 15'h0005; 
        10'b0101100110: data <= 15'h7ff9; 
        10'b0101100111: data <= 15'h7fdc; 
        10'b0101101000: data <= 15'h7fe0; 
        10'b0101101001: data <= 15'h7ff7; 
        10'b0101101010: data <= 15'h0023; 
        10'b0101101011: data <= 15'h0014; 
        10'b0101101100: data <= 15'h0004; 
        10'b0101101101: data <= 15'h0017; 
        10'b0101101110: data <= 15'h0003; 
        10'b0101101111: data <= 15'h000a; 
        10'b0101110000: data <= 15'h001b; 
        10'b0101110001: data <= 15'h004d; 
        10'b0101110010: data <= 15'h009e; 
        10'b0101110011: data <= 15'h00b7; 
        10'b0101110100: data <= 15'h00d2; 
        10'b0101110101: data <= 15'h00b0; 
        10'b0101110110: data <= 15'h00cd; 
        10'b0101110111: data <= 15'h014e; 
        10'b0101111000: data <= 15'h00fd; 
        10'b0101111001: data <= 15'h0004; 
        10'b0101111010: data <= 15'h7fdc; 
        10'b0101111011: data <= 15'h0075; 
        10'b0101111100: data <= 15'h0079; 
        10'b0101111101: data <= 15'h0086; 
        10'b0101111110: data <= 15'h005c; 
        10'b0101111111: data <= 15'h002a; 
        10'b0110000000: data <= 15'h005c; 
        10'b0110000001: data <= 15'h0044; 
        10'b0110000010: data <= 15'h0020; 
        10'b0110000011: data <= 15'h7fed; 
        10'b0110000100: data <= 15'h7fef; 
        10'b0110000101: data <= 15'h0002; 
        10'b0110000110: data <= 15'h001c; 
        10'b0110000111: data <= 15'h0014; 
        10'b0110001000: data <= 15'h0004; 
        10'b0110001001: data <= 15'h001d; 
        10'b0110001010: data <= 15'h0002; 
        10'b0110001011: data <= 15'h0022; 
        10'b0110001100: data <= 15'h0045; 
        10'b0110001101: data <= 15'h008a; 
        10'b0110001110: data <= 15'h00c0; 
        10'b0110001111: data <= 15'h00d2; 
        10'b0110010000: data <= 15'h009d; 
        10'b0110010001: data <= 15'h0096; 
        10'b0110010010: data <= 15'h00b5; 
        10'b0110010011: data <= 15'h00db; 
        10'b0110010100: data <= 15'h009f; 
        10'b0110010101: data <= 15'h000d; 
        10'b0110010110: data <= 15'h7fe9; 
        10'b0110010111: data <= 15'h002a; 
        10'b0110011000: data <= 15'h0086; 
        10'b0110011001: data <= 15'h00dd; 
        10'b0110011010: data <= 15'h0096; 
        10'b0110011011: data <= 15'h008a; 
        10'b0110011100: data <= 15'h004d; 
        10'b0110011101: data <= 15'h0034; 
        10'b0110011110: data <= 15'h0011; 
        10'b0110011111: data <= 15'h0009; 
        10'b0110100000: data <= 15'h7ffb; 
        10'b0110100001: data <= 15'h0009; 
        10'b0110100010: data <= 15'h0011; 
        10'b0110100011: data <= 15'h0008; 
        10'b0110100100: data <= 15'h0018; 
        10'b0110100101: data <= 15'h0022; 
        10'b0110100110: data <= 15'h0016; 
        10'b0110100111: data <= 15'h001c; 
        10'b0110101000: data <= 15'h003e; 
        10'b0110101001: data <= 15'h0046; 
        10'b0110101010: data <= 15'h006d; 
        10'b0110101011: data <= 15'h0065; 
        10'b0110101100: data <= 15'h00a2; 
        10'b0110101101: data <= 15'h008b; 
        10'b0110101110: data <= 15'h0061; 
        10'b0110101111: data <= 15'h0046; 
        10'b0110110000: data <= 15'h0053; 
        10'b0110110001: data <= 15'h0010; 
        10'b0110110010: data <= 15'h0043; 
        10'b0110110011: data <= 15'h005d; 
        10'b0110110100: data <= 15'h00c1; 
        10'b0110110101: data <= 15'h00ac; 
        10'b0110110110: data <= 15'h007b; 
        10'b0110110111: data <= 15'h0049; 
        10'b0110111000: data <= 15'h7fec; 
        10'b0110111001: data <= 15'h001b; 
        10'b0110111010: data <= 15'h0031; 
        10'b0110111011: data <= 15'h0005; 
        10'b0110111100: data <= 15'h7fe3; 
        10'b0110111101: data <= 15'h000f; 
        10'b0110111110: data <= 15'h0004; 
        10'b0110111111: data <= 15'h000a; 
        10'b0111000000: data <= 15'h000b; 
        10'b0111000001: data <= 15'h0000; 
        10'b0111000010: data <= 15'h0001; 
        10'b0111000011: data <= 15'h7ffc; 
        10'b0111000100: data <= 15'h0011; 
        10'b0111000101: data <= 15'h0029; 
        10'b0111000110: data <= 15'h0044; 
        10'b0111000111: data <= 15'h0076; 
        10'b0111001000: data <= 15'h00ac; 
        10'b0111001001: data <= 15'h007a; 
        10'b0111001010: data <= 15'h0021; 
        10'b0111001011: data <= 15'h7ffc; 
        10'b0111001100: data <= 15'h0022; 
        10'b0111001101: data <= 15'h002a; 
        10'b0111001110: data <= 15'h009e; 
        10'b0111001111: data <= 15'h00da; 
        10'b0111010000: data <= 15'h00e1; 
        10'b0111010001: data <= 15'h00bb; 
        10'b0111010010: data <= 15'h007e; 
        10'b0111010011: data <= 15'h0010; 
        10'b0111010100: data <= 15'h0035; 
        10'b0111010101: data <= 15'h004b; 
        10'b0111010110: data <= 15'h0012; 
        10'b0111010111: data <= 15'h7ff4; 
        10'b0111011000: data <= 15'h7ffd; 
        10'b0111011001: data <= 15'h0007; 
        10'b0111011010: data <= 15'h000e; 
        10'b0111011011: data <= 15'h000e; 
        10'b0111011100: data <= 15'h000d; 
        10'b0111011101: data <= 15'h000d; 
        10'b0111011110: data <= 15'h001a; 
        10'b0111011111: data <= 15'h0000; 
        10'b0111100000: data <= 15'h7fee; 
        10'b0111100001: data <= 15'h7fdb; 
        10'b0111100010: data <= 15'h0016; 
        10'b0111100011: data <= 15'h005e; 
        10'b0111100100: data <= 15'h00b5; 
        10'b0111100101: data <= 15'h009d; 
        10'b0111100110: data <= 15'h0039; 
        10'b0111100111: data <= 15'h002d; 
        10'b0111101000: data <= 15'h0041; 
        10'b0111101001: data <= 15'h009b; 
        10'b0111101010: data <= 15'h0100; 
        10'b0111101011: data <= 15'h00cb; 
        10'b0111101100: data <= 15'h00a9; 
        10'b0111101101: data <= 15'h0034; 
        10'b0111101110: data <= 15'h0008; 
        10'b0111101111: data <= 15'h7fc7; 
        10'b0111110000: data <= 15'h0011; 
        10'b0111110001: data <= 15'h0006; 
        10'b0111110010: data <= 15'h7fdd; 
        10'b0111110011: data <= 15'h7ff1; 
        10'b0111110100: data <= 15'h7fe9; 
        10'b0111110101: data <= 15'h7ff3; 
        10'b0111110110: data <= 15'h0017; 
        10'b0111110111: data <= 15'h001c; 
        10'b0111111000: data <= 15'h000e; 
        10'b0111111001: data <= 15'h0015; 
        10'b0111111010: data <= 15'h0013; 
        10'b0111111011: data <= 15'h0003; 
        10'b0111111100: data <= 15'h7fea; 
        10'b0111111101: data <= 15'h7fd2; 
        10'b0111111110: data <= 15'h7fcb; 
        10'b0111111111: data <= 15'h7fff; 
        10'b1000000000: data <= 15'h002e; 
        10'b1000000001: data <= 15'h000b; 
        10'b1000000010: data <= 15'h7fda; 
        10'b1000000011: data <= 15'h7fea; 
        10'b1000000100: data <= 15'h003b; 
        10'b1000000101: data <= 15'h0043; 
        10'b1000000110: data <= 15'h0070; 
        10'b1000000111: data <= 15'h0060; 
        10'b1000001000: data <= 15'h0032; 
        10'b1000001001: data <= 15'h7fb2; 
        10'b1000001010: data <= 15'h7fb6; 
        10'b1000001011: data <= 15'h7f94; 
        10'b1000001100: data <= 15'h7fc0; 
        10'b1000001101: data <= 15'h7fbd; 
        10'b1000001110: data <= 15'h7fa7; 
        10'b1000001111: data <= 15'h7fbb; 
        10'b1000010000: data <= 15'h7fee; 
        10'b1000010001: data <= 15'h7ff7; 
        10'b1000010010: data <= 15'h0008; 
        10'b1000010011: data <= 15'h0001; 
        10'b1000010100: data <= 15'h000e; 
        10'b1000010101: data <= 15'h0019; 
        10'b1000010110: data <= 15'h000a; 
        10'b1000010111: data <= 15'h0006; 
        10'b1000011000: data <= 15'h7fcf; 
        10'b1000011001: data <= 15'h7fc3; 
        10'b1000011010: data <= 15'h7faf; 
        10'b1000011011: data <= 15'h7f86; 
        10'b1000011100: data <= 15'h7f76; 
        10'b1000011101: data <= 15'h7f6d; 
        10'b1000011110: data <= 15'h7f53; 
        10'b1000011111: data <= 15'h7f5a; 
        10'b1000100000: data <= 15'h7f6d; 
        10'b1000100001: data <= 15'h7faa; 
        10'b1000100010: data <= 15'h7fe6; 
        10'b1000100011: data <= 15'h0016; 
        10'b1000100100: data <= 15'h7fbd; 
        10'b1000100101: data <= 15'h7fc7; 
        10'b1000100110: data <= 15'h7fb9; 
        10'b1000100111: data <= 15'h7f9e; 
        10'b1000101000: data <= 15'h7f93; 
        10'b1000101001: data <= 15'h7f9c; 
        10'b1000101010: data <= 15'h7f9a; 
        10'b1000101011: data <= 15'h7fbb; 
        10'b1000101100: data <= 15'h7fee; 
        10'b1000101101: data <= 15'h000e; 
        10'b1000101110: data <= 15'h0018; 
        10'b1000101111: data <= 15'h0016; 
        10'b1000110000: data <= 15'h0024; 
        10'b1000110001: data <= 15'h0021; 
        10'b1000110010: data <= 15'h000a; 
        10'b1000110011: data <= 15'h0006; 
        10'b1000110100: data <= 15'h7fd8; 
        10'b1000110101: data <= 15'h7fbb; 
        10'b1000110110: data <= 15'h7f9c; 
        10'b1000110111: data <= 15'h7f5e; 
        10'b1000111000: data <= 15'h7f3f; 
        10'b1000111001: data <= 15'h7f33; 
        10'b1000111010: data <= 15'h7f30; 
        10'b1000111011: data <= 15'h7f67; 
        10'b1000111100: data <= 15'h7f85; 
        10'b1000111101: data <= 15'h7f76; 
        10'b1000111110: data <= 15'h7fa9; 
        10'b1000111111: data <= 15'h7fd3; 
        10'b1001000000: data <= 15'h7ff0; 
        10'b1001000001: data <= 15'h7ff7; 
        10'b1001000010: data <= 15'h7fdc; 
        10'b1001000011: data <= 15'h7fb2; 
        10'b1001000100: data <= 15'h7fcc; 
        10'b1001000101: data <= 15'h7fc5; 
        10'b1001000110: data <= 15'h7fb9; 
        10'b1001000111: data <= 15'h7fdb; 
        10'b1001001000: data <= 15'h7fdd; 
        10'b1001001001: data <= 15'h0003; 
        10'b1001001010: data <= 15'h0008; 
        10'b1001001011: data <= 15'h0018; 
        10'b1001001100: data <= 15'h0007; 
        10'b1001001101: data <= 15'h000a; 
        10'b1001001110: data <= 15'h0003; 
        10'b1001001111: data <= 15'h0005; 
        10'b1001010000: data <= 15'h0000; 
        10'b1001010001: data <= 15'h7fd9; 
        10'b1001010010: data <= 15'h7f9e; 
        10'b1001010011: data <= 15'h7f76; 
        10'b1001010100: data <= 15'h7f84; 
        10'b1001010101: data <= 15'h7f73; 
        10'b1001010110: data <= 15'h7f85; 
        10'b1001010111: data <= 15'h7fa5; 
        10'b1001011000: data <= 15'h7fb4; 
        10'b1001011001: data <= 15'h7fba; 
        10'b1001011010: data <= 15'h7fb0; 
        10'b1001011011: data <= 15'h7fdb; 
        10'b1001011100: data <= 15'h7fce; 
        10'b1001011101: data <= 15'h0009; 
        10'b1001011110: data <= 15'h7ff1; 
        10'b1001011111: data <= 15'h0003; 
        10'b1001100000: data <= 15'h7ffa; 
        10'b1001100001: data <= 15'h7fd0; 
        10'b1001100010: data <= 15'h7fd7; 
        10'b1001100011: data <= 15'h7ff8; 
        10'b1001100100: data <= 15'h7fff; 
        10'b1001100101: data <= 15'h000f; 
        10'b1001100110: data <= 15'h0014; 
        10'b1001100111: data <= 15'h0013; 
        10'b1001101000: data <= 15'h0011; 
        10'b1001101001: data <= 15'h0014; 
        10'b1001101010: data <= 15'h0008; 
        10'b1001101011: data <= 15'h0016; 
        10'b1001101100: data <= 15'h7ffb; 
        10'b1001101101: data <= 15'h7feb; 
        10'b1001101110: data <= 15'h7fd7; 
        10'b1001101111: data <= 15'h7fbd; 
        10'b1001110000: data <= 15'h7fa5; 
        10'b1001110001: data <= 15'h7fc9; 
        10'b1001110010: data <= 15'h7fc7; 
        10'b1001110011: data <= 15'h7fd9; 
        10'b1001110100: data <= 15'h7fd7; 
        10'b1001110101: data <= 15'h7fdc; 
        10'b1001110110: data <= 15'h7fd4; 
        10'b1001110111: data <= 15'h7fe5; 
        10'b1001111000: data <= 15'h7fe6; 
        10'b1001111001: data <= 15'h0009; 
        10'b1001111010: data <= 15'h0028; 
        10'b1001111011: data <= 15'h0042; 
        10'b1001111100: data <= 15'h0032; 
        10'b1001111101: data <= 15'h0021; 
        10'b1001111110: data <= 15'h7fea; 
        10'b1001111111: data <= 15'h7feb; 
        10'b1010000000: data <= 15'h7fff; 
        10'b1010000001: data <= 15'h000e; 
        10'b1010000010: data <= 15'h0002; 
        10'b1010000011: data <= 15'h000b; 
        10'b1010000100: data <= 15'h000b; 
        10'b1010000101: data <= 15'h0001; 
        10'b1010000110: data <= 15'h000a; 
        10'b1010000111: data <= 15'h0014; 
        10'b1010001000: data <= 15'h000b; 
        10'b1010001001: data <= 15'h000e; 
        10'b1010001010: data <= 15'h7fea; 
        10'b1010001011: data <= 15'h7fe8; 
        10'b1010001100: data <= 15'h7fdf; 
        10'b1010001101: data <= 15'h000f; 
        10'b1010001110: data <= 15'h7fdd; 
        10'b1010001111: data <= 15'h0006; 
        10'b1010010000: data <= 15'h7fdc; 
        10'b1010010001: data <= 15'h7fe4; 
        10'b1010010010: data <= 15'h7fe4; 
        10'b1010010011: data <= 15'h7ffe; 
        10'b1010010100: data <= 15'h0009; 
        10'b1010010101: data <= 15'h0018; 
        10'b1010010110: data <= 15'h004b; 
        10'b1010010111: data <= 15'h004a; 
        10'b1010011000: data <= 15'h003f; 
        10'b1010011001: data <= 15'h001c; 
        10'b1010011010: data <= 15'h7ff6; 
        10'b1010011011: data <= 15'h0008; 
        10'b1010011100: data <= 15'h0011; 
        10'b1010011101: data <= 15'h0017; 
        10'b1010011110: data <= 15'h0007; 
        10'b1010011111: data <= 15'h001c; 
        10'b1010100000: data <= 15'h0015; 
        10'b1010100001: data <= 15'h001f; 
        10'b1010100010: data <= 15'h000e; 
        10'b1010100011: data <= 15'h0018; 
        10'b1010100100: data <= 15'h0006; 
        10'b1010100101: data <= 15'h0013; 
        10'b1010100110: data <= 15'h0007; 
        10'b1010100111: data <= 15'h7fde; 
        10'b1010101000: data <= 15'h7fdd; 
        10'b1010101001: data <= 15'h7ff5; 
        10'b1010101010: data <= 15'h7fdb; 
        10'b1010101011: data <= 15'h7ffa; 
        10'b1010101100: data <= 15'h7fe5; 
        10'b1010101101: data <= 15'h7fe7; 
        10'b1010101110: data <= 15'h7fd2; 
        10'b1010101111: data <= 15'h7fcd; 
        10'b1010110000: data <= 15'h7fea; 
        10'b1010110001: data <= 15'h7ff5; 
        10'b1010110010: data <= 15'h0004; 
        10'b1010110011: data <= 15'h0028; 
        10'b1010110100: data <= 15'h001d; 
        10'b1010110101: data <= 15'h7ff4; 
        10'b1010110110: data <= 15'h7ffd; 
        10'b1010110111: data <= 15'h000f; 
        10'b1010111000: data <= 15'h0019; 
        10'b1010111001: data <= 15'h0004; 
        10'b1010111010: data <= 15'h0007; 
        10'b1010111011: data <= 15'h0016; 
        10'b1010111100: data <= 15'h0020; 
        10'b1010111101: data <= 15'h001f; 
        10'b1010111110: data <= 15'h001c; 
        10'b1010111111: data <= 15'h0006; 
        10'b1011000000: data <= 15'h001d; 
        10'b1011000001: data <= 15'h0001; 
        10'b1011000010: data <= 15'h7fec; 
        10'b1011000011: data <= 15'h7fdf; 
        10'b1011000100: data <= 15'h7fce; 
        10'b1011000101: data <= 15'h7fcb; 
        10'b1011000110: data <= 15'h7faa; 
        10'b1011000111: data <= 15'h7f9f; 
        10'b1011001000: data <= 15'h7fa4; 
        10'b1011001001: data <= 15'h7fa5; 
        10'b1011001010: data <= 15'h7fb2; 
        10'b1011001011: data <= 15'h7fae; 
        10'b1011001100: data <= 15'h7f96; 
        10'b1011001101: data <= 15'h7f87; 
        10'b1011001110: data <= 15'h7f93; 
        10'b1011001111: data <= 15'h7fc4; 
        10'b1011010000: data <= 15'h7fc9; 
        10'b1011010001: data <= 15'h7fec; 
        10'b1011010010: data <= 15'h0001; 
        10'b1011010011: data <= 15'h0015; 
        10'b1011010100: data <= 15'h0002; 
        10'b1011010101: data <= 15'h001d; 
        10'b1011010110: data <= 15'h000c; 
        10'b1011010111: data <= 15'h000b; 
        10'b1011011000: data <= 15'h000f; 
        10'b1011011001: data <= 15'h0016; 
        10'b1011011010: data <= 15'h0005; 
        10'b1011011011: data <= 15'h000e; 
        10'b1011011100: data <= 15'h7fff; 
        10'b1011011101: data <= 15'h7ffb; 
        10'b1011011110: data <= 15'h0009; 
        10'b1011011111: data <= 15'h0006; 
        10'b1011100000: data <= 15'h7ff9; 
        10'b1011100001: data <= 15'h7fe2; 
        10'b1011100010: data <= 15'h7fb7; 
        10'b1011100011: data <= 15'h7fc0; 
        10'b1011100100: data <= 15'h7fb7; 
        10'b1011100101: data <= 15'h7f9d; 
        10'b1011100110: data <= 15'h7f94; 
        10'b1011100111: data <= 15'h7fac; 
        10'b1011101000: data <= 15'h7fa0; 
        10'b1011101001: data <= 15'h7faf; 
        10'b1011101010: data <= 15'h7fbd; 
        10'b1011101011: data <= 15'h7fd8; 
        10'b1011101100: data <= 15'h7ff1; 
        10'b1011101101: data <= 15'h0016; 
        10'b1011101110: data <= 15'h0015; 
        10'b1011101111: data <= 15'h0003; 
        10'b1011110000: data <= 15'h000e; 
        10'b1011110001: data <= 15'h0002; 
        10'b1011110010: data <= 15'h0022; 
        10'b1011110011: data <= 15'h000f; 
        10'b1011110100: data <= 15'h0015; 
        10'b1011110101: data <= 15'h0003; 
        10'b1011110110: data <= 15'h0005; 
        10'b1011110111: data <= 15'h0021; 
        10'b1011111000: data <= 15'h000c; 
        10'b1011111001: data <= 15'h001b; 
        10'b1011111010: data <= 15'h000d; 
        10'b1011111011: data <= 15'h0022; 
        10'b1011111100: data <= 15'h0000; 
        10'b1011111101: data <= 15'h000f; 
        10'b1011111110: data <= 15'h0007; 
        10'b1011111111: data <= 15'h7ffb; 
        10'b1100000000: data <= 15'h7ffd; 
        10'b1100000001: data <= 15'h0001; 
        10'b1100000010: data <= 15'h7ff2; 
        10'b1100000011: data <= 15'h001b; 
        10'b1100000100: data <= 15'h7ff9; 
        10'b1100000101: data <= 15'h7ff8; 
        10'b1100000110: data <= 15'h7ffd; 
        10'b1100000111: data <= 15'h000e; 
        10'b1100001000: data <= 15'h000b; 
        10'b1100001001: data <= 15'h000b; 
        10'b1100001010: data <= 15'h000b; 
        10'b1100001011: data <= 15'h0013; 
        10'b1100001100: data <= 15'h0013; 
        10'b1100001101: data <= 15'h0019; 
        10'b1100001110: data <= 15'h0012; 
        10'b1100001111: data <= 15'h000c; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 10) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 16'h0000; 
        10'b0000000001: data <= 16'h0009; 
        10'b0000000010: data <= 16'h003c; 
        10'b0000000011: data <= 16'h003c; 
        10'b0000000100: data <= 16'h0001; 
        10'b0000000101: data <= 16'h0001; 
        10'b0000000110: data <= 16'h002f; 
        10'b0000000111: data <= 16'h000d; 
        10'b0000001000: data <= 16'h0004; 
        10'b0000001001: data <= 16'h0009; 
        10'b0000001010: data <= 16'h0002; 
        10'b0000001011: data <= 16'h002b; 
        10'b0000001100: data <= 16'h0039; 
        10'b0000001101: data <= 16'h0021; 
        10'b0000001110: data <= 16'h002a; 
        10'b0000001111: data <= 16'h0005; 
        10'b0000010000: data <= 16'h0027; 
        10'b0000010001: data <= 16'h0036; 
        10'b0000010010: data <= 16'h000b; 
        10'b0000010011: data <= 16'h002c; 
        10'b0000010100: data <= 16'h0003; 
        10'b0000010101: data <= 16'h001a; 
        10'b0000010110: data <= 16'h003a; 
        10'b0000010111: data <= 16'h0006; 
        10'b0000011000: data <= 16'h003a; 
        10'b0000011001: data <= 16'h0009; 
        10'b0000011010: data <= 16'h0040; 
        10'b0000011011: data <= 16'h001a; 
        10'b0000011100: data <= 16'h0011; 
        10'b0000011101: data <= 16'h001e; 
        10'b0000011110: data <= 16'h0000; 
        10'b0000011111: data <= 16'h0005; 
        10'b0000100000: data <= 16'h001d; 
        10'b0000100001: data <= 16'h0046; 
        10'b0000100010: data <= 16'h000f; 
        10'b0000100011: data <= 16'hfff5; 
        10'b0000100100: data <= 16'h0027; 
        10'b0000100101: data <= 16'h0001; 
        10'b0000100110: data <= 16'h001a; 
        10'b0000100111: data <= 16'hffec; 
        10'b0000101000: data <= 16'h0012; 
        10'b0000101001: data <= 16'hffe4; 
        10'b0000101010: data <= 16'h0001; 
        10'b0000101011: data <= 16'h0027; 
        10'b0000101100: data <= 16'h002d; 
        10'b0000101101: data <= 16'h000d; 
        10'b0000101110: data <= 16'h0001; 
        10'b0000101111: data <= 16'h000b; 
        10'b0000110000: data <= 16'h0031; 
        10'b0000110001: data <= 16'hffff; 
        10'b0000110010: data <= 16'hfffe; 
        10'b0000110011: data <= 16'h0004; 
        10'b0000110100: data <= 16'h002b; 
        10'b0000110101: data <= 16'h002e; 
        10'b0000110110: data <= 16'h000b; 
        10'b0000110111: data <= 16'h002e; 
        10'b0000111000: data <= 16'h0034; 
        10'b0000111001: data <= 16'h0022; 
        10'b0000111010: data <= 16'h0034; 
        10'b0000111011: data <= 16'h0035; 
        10'b0000111100: data <= 16'h0032; 
        10'b0000111101: data <= 16'h002d; 
        10'b0000111110: data <= 16'h003c; 
        10'b0000111111: data <= 16'hffed; 
        10'b0001000000: data <= 16'hffeb; 
        10'b0001000001: data <= 16'h000b; 
        10'b0001000010: data <= 16'hfff9; 
        10'b0001000011: data <= 16'hffdd; 
        10'b0001000100: data <= 16'hff77; 
        10'b0001000101: data <= 16'hffc9; 
        10'b0001000110: data <= 16'hffbe; 
        10'b0001000111: data <= 16'hffa2; 
        10'b0001001000: data <= 16'hffbc; 
        10'b0001001001: data <= 16'hfff3; 
        10'b0001001010: data <= 16'h0011; 
        10'b0001001011: data <= 16'h0030; 
        10'b0001001100: data <= 16'h003e; 
        10'b0001001101: data <= 16'h0024; 
        10'b0001001110: data <= 16'h003b; 
        10'b0001001111: data <= 16'h0010; 
        10'b0001010000: data <= 16'h0016; 
        10'b0001010001: data <= 16'h0028; 
        10'b0001010010: data <= 16'h0002; 
        10'b0001010011: data <= 16'h001c; 
        10'b0001010100: data <= 16'h0035; 
        10'b0001010101: data <= 16'h0030; 
        10'b0001010110: data <= 16'h0012; 
        10'b0001010111: data <= 16'h001e; 
        10'b0001011000: data <= 16'h001f; 
        10'b0001011001: data <= 16'h0000; 
        10'b0001011010: data <= 16'h0028; 
        10'b0001011011: data <= 16'hffdd; 
        10'b0001011100: data <= 16'hffcd; 
        10'b0001011101: data <= 16'hffe4; 
        10'b0001011110: data <= 16'hff8b; 
        10'b0001011111: data <= 16'hff75; 
        10'b0001100000: data <= 16'hff22; 
        10'b0001100001: data <= 16'hff2c; 
        10'b0001100010: data <= 16'hff37; 
        10'b0001100011: data <= 16'hff0b; 
        10'b0001100100: data <= 16'hff5d; 
        10'b0001100101: data <= 16'hffae; 
        10'b0001100110: data <= 16'h000c; 
        10'b0001100111: data <= 16'h001a; 
        10'b0001101000: data <= 16'h002f; 
        10'b0001101001: data <= 16'h0046; 
        10'b0001101010: data <= 16'h0012; 
        10'b0001101011: data <= 16'h0013; 
        10'b0001101100: data <= 16'h0044; 
        10'b0001101101: data <= 16'h0041; 
        10'b0001101110: data <= 16'h0014; 
        10'b0001101111: data <= 16'h0026; 
        10'b0001110000: data <= 16'h0042; 
        10'b0001110001: data <= 16'h002c; 
        10'b0001110010: data <= 16'h0031; 
        10'b0001110011: data <= 16'h0030; 
        10'b0001110100: data <= 16'h001c; 
        10'b0001110101: data <= 16'h0036; 
        10'b0001110110: data <= 16'hffd7; 
        10'b0001110111: data <= 16'hfff7; 
        10'b0001111000: data <= 16'hffad; 
        10'b0001111001: data <= 16'hffba; 
        10'b0001111010: data <= 16'hff39; 
        10'b0001111011: data <= 16'hff43; 
        10'b0001111100: data <= 16'hfefd; 
        10'b0001111101: data <= 16'hff29; 
        10'b0001111110: data <= 16'hfef8; 
        10'b0001111111: data <= 16'hff1e; 
        10'b0010000000: data <= 16'hff92; 
        10'b0010000001: data <= 16'hff9e; 
        10'b0010000010: data <= 16'hffc6; 
        10'b0010000011: data <= 16'h0038; 
        10'b0010000100: data <= 16'h004d; 
        10'b0010000101: data <= 16'h0058; 
        10'b0010000110: data <= 16'h0054; 
        10'b0010000111: data <= 16'h0070; 
        10'b0010001000: data <= 16'h001f; 
        10'b0010001001: data <= 16'h003f; 
        10'b0010001010: data <= 16'h0010; 
        10'b0010001011: data <= 16'h000a; 
        10'b0010001100: data <= 16'h0043; 
        10'b0010001101: data <= 16'h0013; 
        10'b0010001110: data <= 16'h002f; 
        10'b0010001111: data <= 16'h000f; 
        10'b0010010000: data <= 16'h002b; 
        10'b0010010001: data <= 16'h0009; 
        10'b0010010010: data <= 16'h001f; 
        10'b0010010011: data <= 16'hffdb; 
        10'b0010010100: data <= 16'h000a; 
        10'b0010010101: data <= 16'hffd5; 
        10'b0010010110: data <= 16'hff6f; 
        10'b0010010111: data <= 16'hffa0; 
        10'b0010011000: data <= 16'hff5b; 
        10'b0010011001: data <= 16'hff33; 
        10'b0010011010: data <= 16'hff71; 
        10'b0010011011: data <= 16'hff8a; 
        10'b0010011100: data <= 16'hffec; 
        10'b0010011101: data <= 16'h0012; 
        10'b0010011110: data <= 16'hffe4; 
        10'b0010011111: data <= 16'h0030; 
        10'b0010100000: data <= 16'h003b; 
        10'b0010100001: data <= 16'h004f; 
        10'b0010100010: data <= 16'h00b8; 
        10'b0010100011: data <= 16'h00d0; 
        10'b0010100100: data <= 16'h0071; 
        10'b0010100101: data <= 16'hfff5; 
        10'b0010100110: data <= 16'h0013; 
        10'b0010100111: data <= 16'h000b; 
        10'b0010101000: data <= 16'h003e; 
        10'b0010101001: data <= 16'h0045; 
        10'b0010101010: data <= 16'h0014; 
        10'b0010101011: data <= 16'h0036; 
        10'b0010101100: data <= 16'h003b; 
        10'b0010101101: data <= 16'h0030; 
        10'b0010101110: data <= 16'h0030; 
        10'b0010101111: data <= 16'hfffc; 
        10'b0010110000: data <= 16'hfff5; 
        10'b0010110001: data <= 16'hffc7; 
        10'b0010110010: data <= 16'hff8d; 
        10'b0010110011: data <= 16'hff35; 
        10'b0010110100: data <= 16'hfecc; 
        10'b0010110101: data <= 16'hfe94; 
        10'b0010110110: data <= 16'hfe84; 
        10'b0010110111: data <= 16'hfeb6; 
        10'b0010111000: data <= 16'hfeae; 
        10'b0010111001: data <= 16'hff3a; 
        10'b0010111010: data <= 16'hff33; 
        10'b0010111011: data <= 16'hffa4; 
        10'b0010111100: data <= 16'hffc3; 
        10'b0010111101: data <= 16'hfffb; 
        10'b0010111110: data <= 16'h0108; 
        10'b0010111111: data <= 16'h0115; 
        10'b0011000000: data <= 16'h006b; 
        10'b0011000001: data <= 16'h0054; 
        10'b0011000010: data <= 16'h003c; 
        10'b0011000011: data <= 16'h0003; 
        10'b0011000100: data <= 16'h001d; 
        10'b0011000101: data <= 16'h000f; 
        10'b0011000110: data <= 16'h0015; 
        10'b0011000111: data <= 16'h0025; 
        10'b0011001000: data <= 16'h0015; 
        10'b0011001001: data <= 16'h0032; 
        10'b0011001010: data <= 16'hffe1; 
        10'b0011001011: data <= 16'hfffa; 
        10'b0011001100: data <= 16'hffde; 
        10'b0011001101: data <= 16'hffb2; 
        10'b0011001110: data <= 16'hff3b; 
        10'b0011001111: data <= 16'hfecd; 
        10'b0011010000: data <= 16'hfe71; 
        10'b0011010001: data <= 16'hfee6; 
        10'b0011010010: data <= 16'hfe9f; 
        10'b0011010011: data <= 16'hfe9d; 
        10'b0011010100: data <= 16'hfe93; 
        10'b0011010101: data <= 16'hff17; 
        10'b0011010110: data <= 16'hff11; 
        10'b0011010111: data <= 16'hff5a; 
        10'b0011011000: data <= 16'hff40; 
        10'b0011011001: data <= 16'hffa8; 
        10'b0011011010: data <= 16'h00a3; 
        10'b0011011011: data <= 16'h00dd; 
        10'b0011011100: data <= 16'h0076; 
        10'b0011011101: data <= 16'h0042; 
        10'b0011011110: data <= 16'h003e; 
        10'b0011011111: data <= 16'h0025; 
        10'b0011100000: data <= 16'h003c; 
        10'b0011100001: data <= 16'h0032; 
        10'b0011100010: data <= 16'h0042; 
        10'b0011100011: data <= 16'h000d; 
        10'b0011100100: data <= 16'h0014; 
        10'b0011100101: data <= 16'h001b; 
        10'b0011100110: data <= 16'h0012; 
        10'b0011100111: data <= 16'hfff0; 
        10'b0011101000: data <= 16'hff6b; 
        10'b0011101001: data <= 16'hffb4; 
        10'b0011101010: data <= 16'hff9d; 
        10'b0011101011: data <= 16'hff39; 
        10'b0011101100: data <= 16'hfedd; 
        10'b0011101101: data <= 16'hff46; 
        10'b0011101110: data <= 16'hfe5b; 
        10'b0011101111: data <= 16'hfe4f; 
        10'b0011110000: data <= 16'hfeb0; 
        10'b0011110001: data <= 16'hff2d; 
        10'b0011110010: data <= 16'hff43; 
        10'b0011110011: data <= 16'hffc4; 
        10'b0011110100: data <= 16'hff8d; 
        10'b0011110101: data <= 16'hff8f; 
        10'b0011110110: data <= 16'h004b; 
        10'b0011110111: data <= 16'h0074; 
        10'b0011111000: data <= 16'h0058; 
        10'b0011111001: data <= 16'h0012; 
        10'b0011111010: data <= 16'h0018; 
        10'b0011111011: data <= 16'h002b; 
        10'b0011111100: data <= 16'h0047; 
        10'b0011111101: data <= 16'h003c; 
        10'b0011111110: data <= 16'h0038; 
        10'b0011111111: data <= 16'h000c; 
        10'b0100000000: data <= 16'hffdb; 
        10'b0100000001: data <= 16'h0001; 
        10'b0100000010: data <= 16'hffa4; 
        10'b0100000011: data <= 16'hffbe; 
        10'b0100000100: data <= 16'hffd5; 
        10'b0100000101: data <= 16'hfff2; 
        10'b0100000110: data <= 16'hffcd; 
        10'b0100000111: data <= 16'hffc3; 
        10'b0100001000: data <= 16'hffc1; 
        10'b0100001001: data <= 16'hff58; 
        10'b0100001010: data <= 16'hfda1; 
        10'b0100001011: data <= 16'hfe3a; 
        10'b0100001100: data <= 16'hff92; 
        10'b0100001101: data <= 16'hffaf; 
        10'b0100001110: data <= 16'hffe7; 
        10'b0100001111: data <= 16'h000d; 
        10'b0100010000: data <= 16'hffc0; 
        10'b0100010001: data <= 16'hffc2; 
        10'b0100010010: data <= 16'h001f; 
        10'b0100010011: data <= 16'h0007; 
        10'b0100010100: data <= 16'hffb8; 
        10'b0100010101: data <= 16'hffb5; 
        10'b0100010110: data <= 16'hffdf; 
        10'b0100010111: data <= 16'h0030; 
        10'b0100011000: data <= 16'h0026; 
        10'b0100011001: data <= 16'h001b; 
        10'b0100011010: data <= 16'h001b; 
        10'b0100011011: data <= 16'h0007; 
        10'b0100011100: data <= 16'h001c; 
        10'b0100011101: data <= 16'hffae; 
        10'b0100011110: data <= 16'hff79; 
        10'b0100011111: data <= 16'hffbe; 
        10'b0100100000: data <= 16'h0014; 
        10'b0100100001: data <= 16'h00ad; 
        10'b0100100010: data <= 16'h0069; 
        10'b0100100011: data <= 16'h004e; 
        10'b0100100100: data <= 16'h005e; 
        10'b0100100101: data <= 16'hff18; 
        10'b0100100110: data <= 16'hfd7f; 
        10'b0100100111: data <= 16'hff3d; 
        10'b0100101000: data <= 16'h0016; 
        10'b0100101001: data <= 16'hffe3; 
        10'b0100101010: data <= 16'hffea; 
        10'b0100101011: data <= 16'h0017; 
        10'b0100101100: data <= 16'hff80; 
        10'b0100101101: data <= 16'hffab; 
        10'b0100101110: data <= 16'hfff0; 
        10'b0100101111: data <= 16'hff75; 
        10'b0100110000: data <= 16'hffb1; 
        10'b0100110001: data <= 16'hffce; 
        10'b0100110010: data <= 16'h0028; 
        10'b0100110011: data <= 16'h0042; 
        10'b0100110100: data <= 16'h002c; 
        10'b0100110101: data <= 16'h002e; 
        10'b0100110110: data <= 16'h0027; 
        10'b0100110111: data <= 16'hffe8; 
        10'b0100111000: data <= 16'hfff7; 
        10'b0100111001: data <= 16'hffd2; 
        10'b0100111010: data <= 16'hffd0; 
        10'b0100111011: data <= 16'h0029; 
        10'b0100111100: data <= 16'h0083; 
        10'b0100111101: data <= 16'h00dd; 
        10'b0100111110: data <= 16'h0130; 
        10'b0100111111: data <= 16'h00c1; 
        10'b0101000000: data <= 16'h00da; 
        10'b0101000001: data <= 16'hfe9c; 
        10'b0101000010: data <= 16'hfe1d; 
        10'b0101000011: data <= 16'h003f; 
        10'b0101000100: data <= 16'h00fa; 
        10'b0101000101: data <= 16'h002a; 
        10'b0101000110: data <= 16'hfff2; 
        10'b0101000111: data <= 16'hffd8; 
        10'b0101001000: data <= 16'hff77; 
        10'b0101001001: data <= 16'hff8b; 
        10'b0101001010: data <= 16'hffc4; 
        10'b0101001011: data <= 16'hff94; 
        10'b0101001100: data <= 16'hff88; 
        10'b0101001101: data <= 16'hfff9; 
        10'b0101001110: data <= 16'hfffc; 
        10'b0101001111: data <= 16'h0011; 
        10'b0101010000: data <= 16'h0032; 
        10'b0101010001: data <= 16'h002b; 
        10'b0101010010: data <= 16'h0015; 
        10'b0101010011: data <= 16'h001e; 
        10'b0101010100: data <= 16'hfffd; 
        10'b0101010101: data <= 16'hffd3; 
        10'b0101010110: data <= 16'h0080; 
        10'b0101010111: data <= 16'h00d4; 
        10'b0101011000: data <= 16'h0148; 
        10'b0101011001: data <= 16'h011f; 
        10'b0101011010: data <= 16'h01de; 
        10'b0101011011: data <= 16'h021d; 
        10'b0101011100: data <= 16'h0200; 
        10'b0101011101: data <= 16'hfff8; 
        10'b0101011110: data <= 16'hff01; 
        10'b0101011111: data <= 16'h00c8; 
        10'b0101100000: data <= 16'h0145; 
        10'b0101100001: data <= 16'h0025; 
        10'b0101100010: data <= 16'h000e; 
        10'b0101100011: data <= 16'h002c; 
        10'b0101100100: data <= 16'hfff8; 
        10'b0101100101: data <= 16'h000a; 
        10'b0101100110: data <= 16'hfff1; 
        10'b0101100111: data <= 16'hffb8; 
        10'b0101101000: data <= 16'hffc0; 
        10'b0101101001: data <= 16'hffee; 
        10'b0101101010: data <= 16'h0047; 
        10'b0101101011: data <= 16'h0029; 
        10'b0101101100: data <= 16'h0008; 
        10'b0101101101: data <= 16'h002f; 
        10'b0101101110: data <= 16'h0006; 
        10'b0101101111: data <= 16'h0013; 
        10'b0101110000: data <= 16'h0037; 
        10'b0101110001: data <= 16'h009b; 
        10'b0101110010: data <= 16'h013b; 
        10'b0101110011: data <= 16'h016e; 
        10'b0101110100: data <= 16'h01a5; 
        10'b0101110101: data <= 16'h015f; 
        10'b0101110110: data <= 16'h019a; 
        10'b0101110111: data <= 16'h029c; 
        10'b0101111000: data <= 16'h01fb; 
        10'b0101111001: data <= 16'h0008; 
        10'b0101111010: data <= 16'hffb8; 
        10'b0101111011: data <= 16'h00eb; 
        10'b0101111100: data <= 16'h00f1; 
        10'b0101111101: data <= 16'h010c; 
        10'b0101111110: data <= 16'h00b9; 
        10'b0101111111: data <= 16'h0053; 
        10'b0110000000: data <= 16'h00b9; 
        10'b0110000001: data <= 16'h0088; 
        10'b0110000010: data <= 16'h0041; 
        10'b0110000011: data <= 16'hffda; 
        10'b0110000100: data <= 16'hffdf; 
        10'b0110000101: data <= 16'h0004; 
        10'b0110000110: data <= 16'h0039; 
        10'b0110000111: data <= 16'h0029; 
        10'b0110001000: data <= 16'h0007; 
        10'b0110001001: data <= 16'h003a; 
        10'b0110001010: data <= 16'h0005; 
        10'b0110001011: data <= 16'h0044; 
        10'b0110001100: data <= 16'h0089; 
        10'b0110001101: data <= 16'h0114; 
        10'b0110001110: data <= 16'h0180; 
        10'b0110001111: data <= 16'h01a4; 
        10'b0110010000: data <= 16'h013a; 
        10'b0110010001: data <= 16'h012c; 
        10'b0110010010: data <= 16'h0169; 
        10'b0110010011: data <= 16'h01b6; 
        10'b0110010100: data <= 16'h013f; 
        10'b0110010101: data <= 16'h001a; 
        10'b0110010110: data <= 16'hffd2; 
        10'b0110010111: data <= 16'h0055; 
        10'b0110011000: data <= 16'h010c; 
        10'b0110011001: data <= 16'h01b9; 
        10'b0110011010: data <= 16'h012c; 
        10'b0110011011: data <= 16'h0113; 
        10'b0110011100: data <= 16'h009a; 
        10'b0110011101: data <= 16'h0067; 
        10'b0110011110: data <= 16'h0022; 
        10'b0110011111: data <= 16'h0013; 
        10'b0110100000: data <= 16'hfff5; 
        10'b0110100001: data <= 16'h0012; 
        10'b0110100010: data <= 16'h0023; 
        10'b0110100011: data <= 16'h0010; 
        10'b0110100100: data <= 16'h0030; 
        10'b0110100101: data <= 16'h0045; 
        10'b0110100110: data <= 16'h002c; 
        10'b0110100111: data <= 16'h0039; 
        10'b0110101000: data <= 16'h007c; 
        10'b0110101001: data <= 16'h008d; 
        10'b0110101010: data <= 16'h00db; 
        10'b0110101011: data <= 16'h00c9; 
        10'b0110101100: data <= 16'h0144; 
        10'b0110101101: data <= 16'h0116; 
        10'b0110101110: data <= 16'h00c2; 
        10'b0110101111: data <= 16'h008d; 
        10'b0110110000: data <= 16'h00a6; 
        10'b0110110001: data <= 16'h0021; 
        10'b0110110010: data <= 16'h0085; 
        10'b0110110011: data <= 16'h00ba; 
        10'b0110110100: data <= 16'h0183; 
        10'b0110110101: data <= 16'h0158; 
        10'b0110110110: data <= 16'h00f6; 
        10'b0110110111: data <= 16'h0092; 
        10'b0110111000: data <= 16'hffd9; 
        10'b0110111001: data <= 16'h0036; 
        10'b0110111010: data <= 16'h0062; 
        10'b0110111011: data <= 16'h000a; 
        10'b0110111100: data <= 16'hffc5; 
        10'b0110111101: data <= 16'h001f; 
        10'b0110111110: data <= 16'h0008; 
        10'b0110111111: data <= 16'h0014; 
        10'b0111000000: data <= 16'h0015; 
        10'b0111000001: data <= 16'h0000; 
        10'b0111000010: data <= 16'h0003; 
        10'b0111000011: data <= 16'hfff7; 
        10'b0111000100: data <= 16'h0022; 
        10'b0111000101: data <= 16'h0053; 
        10'b0111000110: data <= 16'h0087; 
        10'b0111000111: data <= 16'h00ec; 
        10'b0111001000: data <= 16'h0158; 
        10'b0111001001: data <= 16'h00f5; 
        10'b0111001010: data <= 16'h0042; 
        10'b0111001011: data <= 16'hfff7; 
        10'b0111001100: data <= 16'h0043; 
        10'b0111001101: data <= 16'h0054; 
        10'b0111001110: data <= 16'h013b; 
        10'b0111001111: data <= 16'h01b4; 
        10'b0111010000: data <= 16'h01c1; 
        10'b0111010001: data <= 16'h0175; 
        10'b0111010010: data <= 16'h00fd; 
        10'b0111010011: data <= 16'h0020; 
        10'b0111010100: data <= 16'h006a; 
        10'b0111010101: data <= 16'h0097; 
        10'b0111010110: data <= 16'h0023; 
        10'b0111010111: data <= 16'hffe7; 
        10'b0111011000: data <= 16'hfff9; 
        10'b0111011001: data <= 16'h000f; 
        10'b0111011010: data <= 16'h001b; 
        10'b0111011011: data <= 16'h001c; 
        10'b0111011100: data <= 16'h0019; 
        10'b0111011101: data <= 16'h001a; 
        10'b0111011110: data <= 16'h0033; 
        10'b0111011111: data <= 16'hffff; 
        10'b0111100000: data <= 16'hffdc; 
        10'b0111100001: data <= 16'hffb6; 
        10'b0111100010: data <= 16'h002c; 
        10'b0111100011: data <= 16'h00bb; 
        10'b0111100100: data <= 16'h0169; 
        10'b0111100101: data <= 16'h0139; 
        10'b0111100110: data <= 16'h0071; 
        10'b0111100111: data <= 16'h0059; 
        10'b0111101000: data <= 16'h0081; 
        10'b0111101001: data <= 16'h0136; 
        10'b0111101010: data <= 16'h0200; 
        10'b0111101011: data <= 16'h0195; 
        10'b0111101100: data <= 16'h0153; 
        10'b0111101101: data <= 16'h0069; 
        10'b0111101110: data <= 16'h0010; 
        10'b0111101111: data <= 16'hff8f; 
        10'b0111110000: data <= 16'h0022; 
        10'b0111110001: data <= 16'h000c; 
        10'b0111110010: data <= 16'hffbb; 
        10'b0111110011: data <= 16'hffe2; 
        10'b0111110100: data <= 16'hffd3; 
        10'b0111110101: data <= 16'hffe6; 
        10'b0111110110: data <= 16'h002e; 
        10'b0111110111: data <= 16'h0038; 
        10'b0111111000: data <= 16'h001c; 
        10'b0111111001: data <= 16'h002b; 
        10'b0111111010: data <= 16'h0025; 
        10'b0111111011: data <= 16'h0006; 
        10'b0111111100: data <= 16'hffd4; 
        10'b0111111101: data <= 16'hffa4; 
        10'b0111111110: data <= 16'hff95; 
        10'b0111111111: data <= 16'hfffe; 
        10'b1000000000: data <= 16'h005c; 
        10'b1000000001: data <= 16'h0015; 
        10'b1000000010: data <= 16'hffb5; 
        10'b1000000011: data <= 16'hffd4; 
        10'b1000000100: data <= 16'h0076; 
        10'b1000000101: data <= 16'h0085; 
        10'b1000000110: data <= 16'h00e1; 
        10'b1000000111: data <= 16'h00c0; 
        10'b1000001000: data <= 16'h0065; 
        10'b1000001001: data <= 16'hff64; 
        10'b1000001010: data <= 16'hff6d; 
        10'b1000001011: data <= 16'hff28; 
        10'b1000001100: data <= 16'hff80; 
        10'b1000001101: data <= 16'hff7b; 
        10'b1000001110: data <= 16'hff4f; 
        10'b1000001111: data <= 16'hff77; 
        10'b1000010000: data <= 16'hffdc; 
        10'b1000010001: data <= 16'hffed; 
        10'b1000010010: data <= 16'h0010; 
        10'b1000010011: data <= 16'h0002; 
        10'b1000010100: data <= 16'h001b; 
        10'b1000010101: data <= 16'h0032; 
        10'b1000010110: data <= 16'h0013; 
        10'b1000010111: data <= 16'h000b; 
        10'b1000011000: data <= 16'hff9d; 
        10'b1000011001: data <= 16'hff85; 
        10'b1000011010: data <= 16'hff5e; 
        10'b1000011011: data <= 16'hff0c; 
        10'b1000011100: data <= 16'hfeed; 
        10'b1000011101: data <= 16'hfedb; 
        10'b1000011110: data <= 16'hfea6; 
        10'b1000011111: data <= 16'hfeb5; 
        10'b1000100000: data <= 16'hfedb; 
        10'b1000100001: data <= 16'hff54; 
        10'b1000100010: data <= 16'hffcd; 
        10'b1000100011: data <= 16'h002d; 
        10'b1000100100: data <= 16'hff7b; 
        10'b1000100101: data <= 16'hff8d; 
        10'b1000100110: data <= 16'hff73; 
        10'b1000100111: data <= 16'hff3d; 
        10'b1000101000: data <= 16'hff26; 
        10'b1000101001: data <= 16'hff37; 
        10'b1000101010: data <= 16'hff34; 
        10'b1000101011: data <= 16'hff76; 
        10'b1000101100: data <= 16'hffdc; 
        10'b1000101101: data <= 16'h001b; 
        10'b1000101110: data <= 16'h0030; 
        10'b1000101111: data <= 16'h002c; 
        10'b1000110000: data <= 16'h0048; 
        10'b1000110001: data <= 16'h0043; 
        10'b1000110010: data <= 16'h0013; 
        10'b1000110011: data <= 16'h000b; 
        10'b1000110100: data <= 16'hffb0; 
        10'b1000110101: data <= 16'hff77; 
        10'b1000110110: data <= 16'hff38; 
        10'b1000110111: data <= 16'hfebb; 
        10'b1000111000: data <= 16'hfe7e; 
        10'b1000111001: data <= 16'hfe67; 
        10'b1000111010: data <= 16'hfe5f; 
        10'b1000111011: data <= 16'hfecf; 
        10'b1000111100: data <= 16'hff09; 
        10'b1000111101: data <= 16'hfeec; 
        10'b1000111110: data <= 16'hff53; 
        10'b1000111111: data <= 16'hffa6; 
        10'b1001000000: data <= 16'hffe1; 
        10'b1001000001: data <= 16'hffef; 
        10'b1001000010: data <= 16'hffb8; 
        10'b1001000011: data <= 16'hff65; 
        10'b1001000100: data <= 16'hff98; 
        10'b1001000101: data <= 16'hff8a; 
        10'b1001000110: data <= 16'hff71; 
        10'b1001000111: data <= 16'hffb7; 
        10'b1001001000: data <= 16'hffba; 
        10'b1001001001: data <= 16'h0005; 
        10'b1001001010: data <= 16'h0011; 
        10'b1001001011: data <= 16'h0030; 
        10'b1001001100: data <= 16'h000d; 
        10'b1001001101: data <= 16'h0015; 
        10'b1001001110: data <= 16'h0005; 
        10'b1001001111: data <= 16'h000a; 
        10'b1001010000: data <= 16'hffff; 
        10'b1001010001: data <= 16'hffb2; 
        10'b1001010010: data <= 16'hff3b; 
        10'b1001010011: data <= 16'hfeec; 
        10'b1001010100: data <= 16'hff08; 
        10'b1001010101: data <= 16'hfee6; 
        10'b1001010110: data <= 16'hff0a; 
        10'b1001010111: data <= 16'hff4a; 
        10'b1001011000: data <= 16'hff68; 
        10'b1001011001: data <= 16'hff74; 
        10'b1001011010: data <= 16'hff5f; 
        10'b1001011011: data <= 16'hffb6; 
        10'b1001011100: data <= 16'hff9d; 
        10'b1001011101: data <= 16'h0012; 
        10'b1001011110: data <= 16'hffe2; 
        10'b1001011111: data <= 16'h0005; 
        10'b1001100000: data <= 16'hfff3; 
        10'b1001100001: data <= 16'hff9f; 
        10'b1001100010: data <= 16'hffae; 
        10'b1001100011: data <= 16'hfff1; 
        10'b1001100100: data <= 16'hfffd; 
        10'b1001100101: data <= 16'h001e; 
        10'b1001100110: data <= 16'h0028; 
        10'b1001100111: data <= 16'h0027; 
        10'b1001101000: data <= 16'h0023; 
        10'b1001101001: data <= 16'h0028; 
        10'b1001101010: data <= 16'h0010; 
        10'b1001101011: data <= 16'h002c; 
        10'b1001101100: data <= 16'hfff6; 
        10'b1001101101: data <= 16'hffd6; 
        10'b1001101110: data <= 16'hffaf; 
        10'b1001101111: data <= 16'hff7a; 
        10'b1001110000: data <= 16'hff4b; 
        10'b1001110001: data <= 16'hff92; 
        10'b1001110010: data <= 16'hff8f; 
        10'b1001110011: data <= 16'hffb1; 
        10'b1001110100: data <= 16'hffad; 
        10'b1001110101: data <= 16'hffb9; 
        10'b1001110110: data <= 16'hffa7; 
        10'b1001110111: data <= 16'hffc9; 
        10'b1001111000: data <= 16'hffcc; 
        10'b1001111001: data <= 16'h0013; 
        10'b1001111010: data <= 16'h0050; 
        10'b1001111011: data <= 16'h0083; 
        10'b1001111100: data <= 16'h0065; 
        10'b1001111101: data <= 16'h0042; 
        10'b1001111110: data <= 16'hffd4; 
        10'b1001111111: data <= 16'hffd5; 
        10'b1010000000: data <= 16'hfffe; 
        10'b1010000001: data <= 16'h001d; 
        10'b1010000010: data <= 16'h0005; 
        10'b1010000011: data <= 16'h0016; 
        10'b1010000100: data <= 16'h0016; 
        10'b1010000101: data <= 16'h0002; 
        10'b1010000110: data <= 16'h0014; 
        10'b1010000111: data <= 16'h0027; 
        10'b1010001000: data <= 16'h0016; 
        10'b1010001001: data <= 16'h001b; 
        10'b1010001010: data <= 16'hffd5; 
        10'b1010001011: data <= 16'hffd0; 
        10'b1010001100: data <= 16'hffbf; 
        10'b1010001101: data <= 16'h001e; 
        10'b1010001110: data <= 16'hffba; 
        10'b1010001111: data <= 16'h000b; 
        10'b1010010000: data <= 16'hffb8; 
        10'b1010010001: data <= 16'hffc7; 
        10'b1010010010: data <= 16'hffc8; 
        10'b1010010011: data <= 16'hfffc; 
        10'b1010010100: data <= 16'h0013; 
        10'b1010010101: data <= 16'h0031; 
        10'b1010010110: data <= 16'h0097; 
        10'b1010010111: data <= 16'h0093; 
        10'b1010011000: data <= 16'h007d; 
        10'b1010011001: data <= 16'h0038; 
        10'b1010011010: data <= 16'hffeb; 
        10'b1010011011: data <= 16'h0011; 
        10'b1010011100: data <= 16'h0021; 
        10'b1010011101: data <= 16'h002e; 
        10'b1010011110: data <= 16'h000f; 
        10'b1010011111: data <= 16'h0039; 
        10'b1010100000: data <= 16'h002b; 
        10'b1010100001: data <= 16'h003d; 
        10'b1010100010: data <= 16'h001d; 
        10'b1010100011: data <= 16'h0030; 
        10'b1010100100: data <= 16'h000b; 
        10'b1010100101: data <= 16'h0025; 
        10'b1010100110: data <= 16'h000e; 
        10'b1010100111: data <= 16'hffbb; 
        10'b1010101000: data <= 16'hffba; 
        10'b1010101001: data <= 16'hffea; 
        10'b1010101010: data <= 16'hffb5; 
        10'b1010101011: data <= 16'hfff4; 
        10'b1010101100: data <= 16'hffca; 
        10'b1010101101: data <= 16'hffcf; 
        10'b1010101110: data <= 16'hffa5; 
        10'b1010101111: data <= 16'hff9a; 
        10'b1010110000: data <= 16'hffd4; 
        10'b1010110001: data <= 16'hffe9; 
        10'b1010110010: data <= 16'h0008; 
        10'b1010110011: data <= 16'h004f; 
        10'b1010110100: data <= 16'h003a; 
        10'b1010110101: data <= 16'hffe8; 
        10'b1010110110: data <= 16'hfff9; 
        10'b1010110111: data <= 16'h001f; 
        10'b1010111000: data <= 16'h0032; 
        10'b1010111001: data <= 16'h0008; 
        10'b1010111010: data <= 16'h000d; 
        10'b1010111011: data <= 16'h002c; 
        10'b1010111100: data <= 16'h0040; 
        10'b1010111101: data <= 16'h003e; 
        10'b1010111110: data <= 16'h0039; 
        10'b1010111111: data <= 16'h000d; 
        10'b1011000000: data <= 16'h0039; 
        10'b1011000001: data <= 16'h0003; 
        10'b1011000010: data <= 16'hffd7; 
        10'b1011000011: data <= 16'hffbe; 
        10'b1011000100: data <= 16'hff9c; 
        10'b1011000101: data <= 16'hff97; 
        10'b1011000110: data <= 16'hff53; 
        10'b1011000111: data <= 16'hff3d; 
        10'b1011001000: data <= 16'hff48; 
        10'b1011001001: data <= 16'hff49; 
        10'b1011001010: data <= 16'hff65; 
        10'b1011001011: data <= 16'hff5b; 
        10'b1011001100: data <= 16'hff2b; 
        10'b1011001101: data <= 16'hff0d; 
        10'b1011001110: data <= 16'hff26; 
        10'b1011001111: data <= 16'hff89; 
        10'b1011010000: data <= 16'hff93; 
        10'b1011010001: data <= 16'hffd9; 
        10'b1011010010: data <= 16'h0002; 
        10'b1011010011: data <= 16'h002a; 
        10'b1011010100: data <= 16'h0003; 
        10'b1011010101: data <= 16'h003a; 
        10'b1011010110: data <= 16'h0017; 
        10'b1011010111: data <= 16'h0015; 
        10'b1011011000: data <= 16'h001e; 
        10'b1011011001: data <= 16'h002b; 
        10'b1011011010: data <= 16'h000a; 
        10'b1011011011: data <= 16'h001d; 
        10'b1011011100: data <= 16'hfffd; 
        10'b1011011101: data <= 16'hfff6; 
        10'b1011011110: data <= 16'h0011; 
        10'b1011011111: data <= 16'h000d; 
        10'b1011100000: data <= 16'hfff3; 
        10'b1011100001: data <= 16'hffc4; 
        10'b1011100010: data <= 16'hff6e; 
        10'b1011100011: data <= 16'hff81; 
        10'b1011100100: data <= 16'hff6e; 
        10'b1011100101: data <= 16'hff3a; 
        10'b1011100110: data <= 16'hff28; 
        10'b1011100111: data <= 16'hff58; 
        10'b1011101000: data <= 16'hff41; 
        10'b1011101001: data <= 16'hff5d; 
        10'b1011101010: data <= 16'hff7b; 
        10'b1011101011: data <= 16'hffb0; 
        10'b1011101100: data <= 16'hffe3; 
        10'b1011101101: data <= 16'h002b; 
        10'b1011101110: data <= 16'h002b; 
        10'b1011101111: data <= 16'h0005; 
        10'b1011110000: data <= 16'h001c; 
        10'b1011110001: data <= 16'h0005; 
        10'b1011110010: data <= 16'h0045; 
        10'b1011110011: data <= 16'h001e; 
        10'b1011110100: data <= 16'h002a; 
        10'b1011110101: data <= 16'h0006; 
        10'b1011110110: data <= 16'h0009; 
        10'b1011110111: data <= 16'h0042; 
        10'b1011111000: data <= 16'h0019; 
        10'b1011111001: data <= 16'h0037; 
        10'b1011111010: data <= 16'h0019; 
        10'b1011111011: data <= 16'h0043; 
        10'b1011111100: data <= 16'h0000; 
        10'b1011111101: data <= 16'h001d; 
        10'b1011111110: data <= 16'h000f; 
        10'b1011111111: data <= 16'hfff7; 
        10'b1100000000: data <= 16'hfff9; 
        10'b1100000001: data <= 16'h0002; 
        10'b1100000010: data <= 16'hffe4; 
        10'b1100000011: data <= 16'h0035; 
        10'b1100000100: data <= 16'hfff2; 
        10'b1100000101: data <= 16'hfff0; 
        10'b1100000110: data <= 16'hfffb; 
        10'b1100000111: data <= 16'h001c; 
        10'b1100001000: data <= 16'h0016; 
        10'b1100001001: data <= 16'h0015; 
        10'b1100001010: data <= 16'h0017; 
        10'b1100001011: data <= 16'h0027; 
        10'b1100001100: data <= 16'h0025; 
        10'b1100001101: data <= 16'h0031; 
        10'b1100001110: data <= 16'h0023; 
        10'b1100001111: data <= 16'h0017; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 11) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 17'h00000; 
        10'b0000000001: data <= 17'h00012; 
        10'b0000000010: data <= 17'h00079; 
        10'b0000000011: data <= 17'h00079; 
        10'b0000000100: data <= 17'h00002; 
        10'b0000000101: data <= 17'h00002; 
        10'b0000000110: data <= 17'h0005f; 
        10'b0000000111: data <= 17'h0001a; 
        10'b0000001000: data <= 17'h00008; 
        10'b0000001001: data <= 17'h00012; 
        10'b0000001010: data <= 17'h00003; 
        10'b0000001011: data <= 17'h00057; 
        10'b0000001100: data <= 17'h00072; 
        10'b0000001101: data <= 17'h00041; 
        10'b0000001110: data <= 17'h00054; 
        10'b0000001111: data <= 17'h00009; 
        10'b0000010000: data <= 17'h0004f; 
        10'b0000010001: data <= 17'h0006c; 
        10'b0000010010: data <= 17'h00017; 
        10'b0000010011: data <= 17'h00057; 
        10'b0000010100: data <= 17'h00007; 
        10'b0000010101: data <= 17'h00034; 
        10'b0000010110: data <= 17'h00074; 
        10'b0000010111: data <= 17'h0000c; 
        10'b0000011000: data <= 17'h00074; 
        10'b0000011001: data <= 17'h00012; 
        10'b0000011010: data <= 17'h0007f; 
        10'b0000011011: data <= 17'h00034; 
        10'b0000011100: data <= 17'h00021; 
        10'b0000011101: data <= 17'h0003c; 
        10'b0000011110: data <= 17'h1ffff; 
        10'b0000011111: data <= 17'h0000a; 
        10'b0000100000: data <= 17'h0003a; 
        10'b0000100001: data <= 17'h0008c; 
        10'b0000100010: data <= 17'h0001d; 
        10'b0000100011: data <= 17'h1ffe9; 
        10'b0000100100: data <= 17'h0004e; 
        10'b0000100101: data <= 17'h00003; 
        10'b0000100110: data <= 17'h00034; 
        10'b0000100111: data <= 17'h1ffd7; 
        10'b0000101000: data <= 17'h00024; 
        10'b0000101001: data <= 17'h1ffc8; 
        10'b0000101010: data <= 17'h00003; 
        10'b0000101011: data <= 17'h0004d; 
        10'b0000101100: data <= 17'h0005b; 
        10'b0000101101: data <= 17'h0001b; 
        10'b0000101110: data <= 17'h00001; 
        10'b0000101111: data <= 17'h00017; 
        10'b0000110000: data <= 17'h00062; 
        10'b0000110001: data <= 17'h1fffe; 
        10'b0000110010: data <= 17'h1fffd; 
        10'b0000110011: data <= 17'h00008; 
        10'b0000110100: data <= 17'h00057; 
        10'b0000110101: data <= 17'h0005c; 
        10'b0000110110: data <= 17'h00016; 
        10'b0000110111: data <= 17'h0005b; 
        10'b0000111000: data <= 17'h00069; 
        10'b0000111001: data <= 17'h00044; 
        10'b0000111010: data <= 17'h00068; 
        10'b0000111011: data <= 17'h0006a; 
        10'b0000111100: data <= 17'h00065; 
        10'b0000111101: data <= 17'h0005a; 
        10'b0000111110: data <= 17'h00077; 
        10'b0000111111: data <= 17'h1ffda; 
        10'b0001000000: data <= 17'h1ffd7; 
        10'b0001000001: data <= 17'h00016; 
        10'b0001000010: data <= 17'h1fff2; 
        10'b0001000011: data <= 17'h1ffb9; 
        10'b0001000100: data <= 17'h1feef; 
        10'b0001000101: data <= 17'h1ff92; 
        10'b0001000110: data <= 17'h1ff7c; 
        10'b0001000111: data <= 17'h1ff45; 
        10'b0001001000: data <= 17'h1ff78; 
        10'b0001001001: data <= 17'h1ffe5; 
        10'b0001001010: data <= 17'h00022; 
        10'b0001001011: data <= 17'h00060; 
        10'b0001001100: data <= 17'h0007d; 
        10'b0001001101: data <= 17'h00048; 
        10'b0001001110: data <= 17'h00076; 
        10'b0001001111: data <= 17'h00020; 
        10'b0001010000: data <= 17'h0002d; 
        10'b0001010001: data <= 17'h00050; 
        10'b0001010010: data <= 17'h00005; 
        10'b0001010011: data <= 17'h00037; 
        10'b0001010100: data <= 17'h0006a; 
        10'b0001010101: data <= 17'h0005f; 
        10'b0001010110: data <= 17'h00025; 
        10'b0001010111: data <= 17'h0003c; 
        10'b0001011000: data <= 17'h0003e; 
        10'b0001011001: data <= 17'h00001; 
        10'b0001011010: data <= 17'h0004f; 
        10'b0001011011: data <= 17'h1ffba; 
        10'b0001011100: data <= 17'h1ff99; 
        10'b0001011101: data <= 17'h1ffc8; 
        10'b0001011110: data <= 17'h1ff15; 
        10'b0001011111: data <= 17'h1feea; 
        10'b0001100000: data <= 17'h1fe44; 
        10'b0001100001: data <= 17'h1fe59; 
        10'b0001100010: data <= 17'h1fe6d; 
        10'b0001100011: data <= 17'h1fe17; 
        10'b0001100100: data <= 17'h1feba; 
        10'b0001100101: data <= 17'h1ff5d; 
        10'b0001100110: data <= 17'h00018; 
        10'b0001100111: data <= 17'h00034; 
        10'b0001101000: data <= 17'h0005f; 
        10'b0001101001: data <= 17'h0008c; 
        10'b0001101010: data <= 17'h00025; 
        10'b0001101011: data <= 17'h00025; 
        10'b0001101100: data <= 17'h00088; 
        10'b0001101101: data <= 17'h00082; 
        10'b0001101110: data <= 17'h00028; 
        10'b0001101111: data <= 17'h0004d; 
        10'b0001110000: data <= 17'h00084; 
        10'b0001110001: data <= 17'h00058; 
        10'b0001110010: data <= 17'h00063; 
        10'b0001110011: data <= 17'h00060; 
        10'b0001110100: data <= 17'h00039; 
        10'b0001110101: data <= 17'h0006c; 
        10'b0001110110: data <= 17'h1ffaf; 
        10'b0001110111: data <= 17'h1ffee; 
        10'b0001111000: data <= 17'h1ff5b; 
        10'b0001111001: data <= 17'h1ff74; 
        10'b0001111010: data <= 17'h1fe72; 
        10'b0001111011: data <= 17'h1fe86; 
        10'b0001111100: data <= 17'h1fdfb; 
        10'b0001111101: data <= 17'h1fe52; 
        10'b0001111110: data <= 17'h1fdf0; 
        10'b0001111111: data <= 17'h1fe3c; 
        10'b0010000000: data <= 17'h1ff25; 
        10'b0010000001: data <= 17'h1ff3d; 
        10'b0010000010: data <= 17'h1ff8b; 
        10'b0010000011: data <= 17'h00070; 
        10'b0010000100: data <= 17'h0009b; 
        10'b0010000101: data <= 17'h000b1; 
        10'b0010000110: data <= 17'h000a8; 
        10'b0010000111: data <= 17'h000df; 
        10'b0010001000: data <= 17'h0003e; 
        10'b0010001001: data <= 17'h0007d; 
        10'b0010001010: data <= 17'h00020; 
        10'b0010001011: data <= 17'h00015; 
        10'b0010001100: data <= 17'h00086; 
        10'b0010001101: data <= 17'h00026; 
        10'b0010001110: data <= 17'h0005f; 
        10'b0010001111: data <= 17'h0001f; 
        10'b0010010000: data <= 17'h00057; 
        10'b0010010001: data <= 17'h00012; 
        10'b0010010010: data <= 17'h0003d; 
        10'b0010010011: data <= 17'h1ffb5; 
        10'b0010010100: data <= 17'h00014; 
        10'b0010010101: data <= 17'h1ffaa; 
        10'b0010010110: data <= 17'h1fedd; 
        10'b0010010111: data <= 17'h1ff3f; 
        10'b0010011000: data <= 17'h1feb5; 
        10'b0010011001: data <= 17'h1fe66; 
        10'b0010011010: data <= 17'h1fee1; 
        10'b0010011011: data <= 17'h1ff13; 
        10'b0010011100: data <= 17'h1ffd8; 
        10'b0010011101: data <= 17'h00024; 
        10'b0010011110: data <= 17'h1ffc7; 
        10'b0010011111: data <= 17'h00060; 
        10'b0010100000: data <= 17'h00075; 
        10'b0010100001: data <= 17'h0009e; 
        10'b0010100010: data <= 17'h00171; 
        10'b0010100011: data <= 17'h001a0; 
        10'b0010100100: data <= 17'h000e2; 
        10'b0010100101: data <= 17'h1ffea; 
        10'b0010100110: data <= 17'h00025; 
        10'b0010100111: data <= 17'h00016; 
        10'b0010101000: data <= 17'h0007d; 
        10'b0010101001: data <= 17'h0008a; 
        10'b0010101010: data <= 17'h00029; 
        10'b0010101011: data <= 17'h0006c; 
        10'b0010101100: data <= 17'h00076; 
        10'b0010101101: data <= 17'h00061; 
        10'b0010101110: data <= 17'h00060; 
        10'b0010101111: data <= 17'h1fff8; 
        10'b0010110000: data <= 17'h1ffea; 
        10'b0010110001: data <= 17'h1ff8e; 
        10'b0010110010: data <= 17'h1ff19; 
        10'b0010110011: data <= 17'h1fe6a; 
        10'b0010110100: data <= 17'h1fd99; 
        10'b0010110101: data <= 17'h1fd29; 
        10'b0010110110: data <= 17'h1fd09; 
        10'b0010110111: data <= 17'h1fd6d; 
        10'b0010111000: data <= 17'h1fd5d; 
        10'b0010111001: data <= 17'h1fe74; 
        10'b0010111010: data <= 17'h1fe67; 
        10'b0010111011: data <= 17'h1ff48; 
        10'b0010111100: data <= 17'h1ff87; 
        10'b0010111101: data <= 17'h1fff7; 
        10'b0010111110: data <= 17'h00210; 
        10'b0010111111: data <= 17'h0022b; 
        10'b0011000000: data <= 17'h000d5; 
        10'b0011000001: data <= 17'h000a7; 
        10'b0011000010: data <= 17'h00078; 
        10'b0011000011: data <= 17'h00005; 
        10'b0011000100: data <= 17'h0003b; 
        10'b0011000101: data <= 17'h0001f; 
        10'b0011000110: data <= 17'h0002a; 
        10'b0011000111: data <= 17'h0004b; 
        10'b0011001000: data <= 17'h0002b; 
        10'b0011001001: data <= 17'h00064; 
        10'b0011001010: data <= 17'h1ffc2; 
        10'b0011001011: data <= 17'h1fff5; 
        10'b0011001100: data <= 17'h1ffbb; 
        10'b0011001101: data <= 17'h1ff64; 
        10'b0011001110: data <= 17'h1fe76; 
        10'b0011001111: data <= 17'h1fd9a; 
        10'b0011010000: data <= 17'h1fce2; 
        10'b0011010001: data <= 17'h1fdcc; 
        10'b0011010010: data <= 17'h1fd3f; 
        10'b0011010011: data <= 17'h1fd39; 
        10'b0011010100: data <= 17'h1fd25; 
        10'b0011010101: data <= 17'h1fe2e; 
        10'b0011010110: data <= 17'h1fe23; 
        10'b0011010111: data <= 17'h1feb4; 
        10'b0011011000: data <= 17'h1fe80; 
        10'b0011011001: data <= 17'h1ff51; 
        10'b0011011010: data <= 17'h00146; 
        10'b0011011011: data <= 17'h001b9; 
        10'b0011011100: data <= 17'h000eb; 
        10'b0011011101: data <= 17'h00085; 
        10'b0011011110: data <= 17'h0007c; 
        10'b0011011111: data <= 17'h0004a; 
        10'b0011100000: data <= 17'h00078; 
        10'b0011100001: data <= 17'h00065; 
        10'b0011100010: data <= 17'h00084; 
        10'b0011100011: data <= 17'h0001a; 
        10'b0011100100: data <= 17'h00028; 
        10'b0011100101: data <= 17'h00037; 
        10'b0011100110: data <= 17'h00025; 
        10'b0011100111: data <= 17'h1ffe0; 
        10'b0011101000: data <= 17'h1fed7; 
        10'b0011101001: data <= 17'h1ff69; 
        10'b0011101010: data <= 17'h1ff3b; 
        10'b0011101011: data <= 17'h1fe73; 
        10'b0011101100: data <= 17'h1fdbb; 
        10'b0011101101: data <= 17'h1fe8c; 
        10'b0011101110: data <= 17'h1fcb5; 
        10'b0011101111: data <= 17'h1fc9f; 
        10'b0011110000: data <= 17'h1fd5f; 
        10'b0011110001: data <= 17'h1fe5b; 
        10'b0011110010: data <= 17'h1fe86; 
        10'b0011110011: data <= 17'h1ff89; 
        10'b0011110100: data <= 17'h1ff19; 
        10'b0011110101: data <= 17'h1ff1d; 
        10'b0011110110: data <= 17'h00096; 
        10'b0011110111: data <= 17'h000e7; 
        10'b0011111000: data <= 17'h000b0; 
        10'b0011111001: data <= 17'h00023; 
        10'b0011111010: data <= 17'h00030; 
        10'b0011111011: data <= 17'h00056; 
        10'b0011111100: data <= 17'h0008e; 
        10'b0011111101: data <= 17'h00078; 
        10'b0011111110: data <= 17'h00070; 
        10'b0011111111: data <= 17'h00017; 
        10'b0100000000: data <= 17'h1ffb6; 
        10'b0100000001: data <= 17'h00002; 
        10'b0100000010: data <= 17'h1ff49; 
        10'b0100000011: data <= 17'h1ff7d; 
        10'b0100000100: data <= 17'h1ffab; 
        10'b0100000101: data <= 17'h1ffe4; 
        10'b0100000110: data <= 17'h1ff9a; 
        10'b0100000111: data <= 17'h1ff86; 
        10'b0100001000: data <= 17'h1ff82; 
        10'b0100001001: data <= 17'h1feb1; 
        10'b0100001010: data <= 17'h1fb42; 
        10'b0100001011: data <= 17'h1fc73; 
        10'b0100001100: data <= 17'h1ff24; 
        10'b0100001101: data <= 17'h1ff5d; 
        10'b0100001110: data <= 17'h1ffce; 
        10'b0100001111: data <= 17'h0001b; 
        10'b0100010000: data <= 17'h1ff80; 
        10'b0100010001: data <= 17'h1ff83; 
        10'b0100010010: data <= 17'h0003f; 
        10'b0100010011: data <= 17'h0000e; 
        10'b0100010100: data <= 17'h1ff6f; 
        10'b0100010101: data <= 17'h1ff6a; 
        10'b0100010110: data <= 17'h1ffbf; 
        10'b0100010111: data <= 17'h00060; 
        10'b0100011000: data <= 17'h0004c; 
        10'b0100011001: data <= 17'h00036; 
        10'b0100011010: data <= 17'h00036; 
        10'b0100011011: data <= 17'h0000f; 
        10'b0100011100: data <= 17'h00039; 
        10'b0100011101: data <= 17'h1ff5c; 
        10'b0100011110: data <= 17'h1fef2; 
        10'b0100011111: data <= 17'h1ff7d; 
        10'b0100100000: data <= 17'h00027; 
        10'b0100100001: data <= 17'h0015a; 
        10'b0100100010: data <= 17'h000d1; 
        10'b0100100011: data <= 17'h0009d; 
        10'b0100100100: data <= 17'h000bb; 
        10'b0100100101: data <= 17'h1fe30; 
        10'b0100100110: data <= 17'h1fafe; 
        10'b0100100111: data <= 17'h1fe79; 
        10'b0100101000: data <= 17'h0002d; 
        10'b0100101001: data <= 17'h1ffc6; 
        10'b0100101010: data <= 17'h1ffd4; 
        10'b0100101011: data <= 17'h0002d; 
        10'b0100101100: data <= 17'h1ff00; 
        10'b0100101101: data <= 17'h1ff57; 
        10'b0100101110: data <= 17'h1ffe0; 
        10'b0100101111: data <= 17'h1fee9; 
        10'b0100110000: data <= 17'h1ff62; 
        10'b0100110001: data <= 17'h1ff9c; 
        10'b0100110010: data <= 17'h00050; 
        10'b0100110011: data <= 17'h00084; 
        10'b0100110100: data <= 17'h00059; 
        10'b0100110101: data <= 17'h0005d; 
        10'b0100110110: data <= 17'h0004e; 
        10'b0100110111: data <= 17'h1ffcf; 
        10'b0100111000: data <= 17'h1ffee; 
        10'b0100111001: data <= 17'h1ffa5; 
        10'b0100111010: data <= 17'h1ff9f; 
        10'b0100111011: data <= 17'h00052; 
        10'b0100111100: data <= 17'h00106; 
        10'b0100111101: data <= 17'h001b9; 
        10'b0100111110: data <= 17'h00260; 
        10'b0100111111: data <= 17'h00183; 
        10'b0101000000: data <= 17'h001b5; 
        10'b0101000001: data <= 17'h1fd39; 
        10'b0101000010: data <= 17'h1fc3a; 
        10'b0101000011: data <= 17'h0007d; 
        10'b0101000100: data <= 17'h001f3; 
        10'b0101000101: data <= 17'h00054; 
        10'b0101000110: data <= 17'h1ffe3; 
        10'b0101000111: data <= 17'h1ffb0; 
        10'b0101001000: data <= 17'h1feef; 
        10'b0101001001: data <= 17'h1ff16; 
        10'b0101001010: data <= 17'h1ff89; 
        10'b0101001011: data <= 17'h1ff28; 
        10'b0101001100: data <= 17'h1ff10; 
        10'b0101001101: data <= 17'h1fff2; 
        10'b0101001110: data <= 17'h1fff8; 
        10'b0101001111: data <= 17'h00021; 
        10'b0101010000: data <= 17'h00063; 
        10'b0101010001: data <= 17'h00057; 
        10'b0101010010: data <= 17'h00029; 
        10'b0101010011: data <= 17'h0003c; 
        10'b0101010100: data <= 17'h1fffa; 
        10'b0101010101: data <= 17'h1ffa7; 
        10'b0101010110: data <= 17'h00101; 
        10'b0101010111: data <= 17'h001a7; 
        10'b0101011000: data <= 17'h00290; 
        10'b0101011001: data <= 17'h0023f; 
        10'b0101011010: data <= 17'h003bc; 
        10'b0101011011: data <= 17'h0043b; 
        10'b0101011100: data <= 17'h00400; 
        10'b0101011101: data <= 17'h1ffef; 
        10'b0101011110: data <= 17'h1fe03; 
        10'b0101011111: data <= 17'h00191; 
        10'b0101100000: data <= 17'h0028b; 
        10'b0101100001: data <= 17'h0004a; 
        10'b0101100010: data <= 17'h0001b; 
        10'b0101100011: data <= 17'h00059; 
        10'b0101100100: data <= 17'h1fff0; 
        10'b0101100101: data <= 17'h00013; 
        10'b0101100110: data <= 17'h1ffe3; 
        10'b0101100111: data <= 17'h1ff71; 
        10'b0101101000: data <= 17'h1ff80; 
        10'b0101101001: data <= 17'h1ffdc; 
        10'b0101101010: data <= 17'h0008d; 
        10'b0101101011: data <= 17'h00052; 
        10'b0101101100: data <= 17'h0000f; 
        10'b0101101101: data <= 17'h0005d; 
        10'b0101101110: data <= 17'h0000d; 
        10'b0101101111: data <= 17'h00027; 
        10'b0101110000: data <= 17'h0006e; 
        10'b0101110001: data <= 17'h00136; 
        10'b0101110010: data <= 17'h00277; 
        10'b0101110011: data <= 17'h002dc; 
        10'b0101110100: data <= 17'h00349; 
        10'b0101110101: data <= 17'h002bf; 
        10'b0101110110: data <= 17'h00334; 
        10'b0101110111: data <= 17'h00538; 
        10'b0101111000: data <= 17'h003f5; 
        10'b0101111001: data <= 17'h0000f; 
        10'b0101111010: data <= 17'h1ff70; 
        10'b0101111011: data <= 17'h001d5; 
        10'b0101111100: data <= 17'h001e2; 
        10'b0101111101: data <= 17'h00218; 
        10'b0101111110: data <= 17'h00171; 
        10'b0101111111: data <= 17'h000a6; 
        10'b0110000000: data <= 17'h00172; 
        10'b0110000001: data <= 17'h00110; 
        10'b0110000010: data <= 17'h00082; 
        10'b0110000011: data <= 17'h1ffb4; 
        10'b0110000100: data <= 17'h1ffbe; 
        10'b0110000101: data <= 17'h00007; 
        10'b0110000110: data <= 17'h00071; 
        10'b0110000111: data <= 17'h00051; 
        10'b0110001000: data <= 17'h0000e; 
        10'b0110001001: data <= 17'h00074; 
        10'b0110001010: data <= 17'h00009; 
        10'b0110001011: data <= 17'h00088; 
        10'b0110001100: data <= 17'h00112; 
        10'b0110001101: data <= 17'h00228; 
        10'b0110001110: data <= 17'h00300; 
        10'b0110001111: data <= 17'h00348; 
        10'b0110010000: data <= 17'h00274; 
        10'b0110010001: data <= 17'h00258; 
        10'b0110010010: data <= 17'h002d3; 
        10'b0110010011: data <= 17'h0036c; 
        10'b0110010100: data <= 17'h0027e; 
        10'b0110010101: data <= 17'h00035; 
        10'b0110010110: data <= 17'h1ffa3; 
        10'b0110010111: data <= 17'h000aa; 
        10'b0110011000: data <= 17'h00219; 
        10'b0110011001: data <= 17'h00372; 
        10'b0110011010: data <= 17'h00257; 
        10'b0110011011: data <= 17'h00227; 
        10'b0110011100: data <= 17'h00134; 
        10'b0110011101: data <= 17'h000cf; 
        10'b0110011110: data <= 17'h00043; 
        10'b0110011111: data <= 17'h00026; 
        10'b0110100000: data <= 17'h1ffea; 
        10'b0110100001: data <= 17'h00025; 
        10'b0110100010: data <= 17'h00045; 
        10'b0110100011: data <= 17'h00021; 
        10'b0110100100: data <= 17'h00060; 
        10'b0110100101: data <= 17'h00089; 
        10'b0110100110: data <= 17'h00058; 
        10'b0110100111: data <= 17'h00072; 
        10'b0110101000: data <= 17'h000f8; 
        10'b0110101001: data <= 17'h00119; 
        10'b0110101010: data <= 17'h001b5; 
        10'b0110101011: data <= 17'h00193; 
        10'b0110101100: data <= 17'h00288; 
        10'b0110101101: data <= 17'h0022c; 
        10'b0110101110: data <= 17'h00183; 
        10'b0110101111: data <= 17'h00119; 
        10'b0110110000: data <= 17'h0014c; 
        10'b0110110001: data <= 17'h00042; 
        10'b0110110010: data <= 17'h0010b; 
        10'b0110110011: data <= 17'h00175; 
        10'b0110110100: data <= 17'h00306; 
        10'b0110110101: data <= 17'h002b0; 
        10'b0110110110: data <= 17'h001ec; 
        10'b0110110111: data <= 17'h00123; 
        10'b0110111000: data <= 17'h1ffb2; 
        10'b0110111001: data <= 17'h0006c; 
        10'b0110111010: data <= 17'h000c3; 
        10'b0110111011: data <= 17'h00015; 
        10'b0110111100: data <= 17'h1ff8a; 
        10'b0110111101: data <= 17'h0003e; 
        10'b0110111110: data <= 17'h00010; 
        10'b0110111111: data <= 17'h00027; 
        10'b0111000000: data <= 17'h0002b; 
        10'b0111000001: data <= 17'h00001; 
        10'b0111000010: data <= 17'h00005; 
        10'b0111000011: data <= 17'h1ffef; 
        10'b0111000100: data <= 17'h00043; 
        10'b0111000101: data <= 17'h000a6; 
        10'b0111000110: data <= 17'h0010e; 
        10'b0111000111: data <= 17'h001d8; 
        10'b0111001000: data <= 17'h002b0; 
        10'b0111001001: data <= 17'h001ea; 
        10'b0111001010: data <= 17'h00083; 
        10'b0111001011: data <= 17'h1ffee; 
        10'b0111001100: data <= 17'h00087; 
        10'b0111001101: data <= 17'h000a8; 
        10'b0111001110: data <= 17'h00277; 
        10'b0111001111: data <= 17'h00369; 
        10'b0111010000: data <= 17'h00383; 
        10'b0111010001: data <= 17'h002eb; 
        10'b0111010010: data <= 17'h001f9; 
        10'b0111010011: data <= 17'h0003f; 
        10'b0111010100: data <= 17'h000d4; 
        10'b0111010101: data <= 17'h0012d; 
        10'b0111010110: data <= 17'h00046; 
        10'b0111010111: data <= 17'h1ffce; 
        10'b0111011000: data <= 17'h1fff2; 
        10'b0111011001: data <= 17'h0001d; 
        10'b0111011010: data <= 17'h00036; 
        10'b0111011011: data <= 17'h00039; 
        10'b0111011100: data <= 17'h00033; 
        10'b0111011101: data <= 17'h00034; 
        10'b0111011110: data <= 17'h00067; 
        10'b0111011111: data <= 17'h1fffe; 
        10'b0111100000: data <= 17'h1ffb8; 
        10'b0111100001: data <= 17'h1ff6c; 
        10'b0111100010: data <= 17'h00058; 
        10'b0111100011: data <= 17'h00177; 
        10'b0111100100: data <= 17'h002d2; 
        10'b0111100101: data <= 17'h00272; 
        10'b0111100110: data <= 17'h000e3; 
        10'b0111100111: data <= 17'h000b2; 
        10'b0111101000: data <= 17'h00102; 
        10'b0111101001: data <= 17'h0026c; 
        10'b0111101010: data <= 17'h00400; 
        10'b0111101011: data <= 17'h0032a; 
        10'b0111101100: data <= 17'h002a6; 
        10'b0111101101: data <= 17'h000d1; 
        10'b0111101110: data <= 17'h00020; 
        10'b0111101111: data <= 17'h1ff1d; 
        10'b0111110000: data <= 17'h00044; 
        10'b0111110001: data <= 17'h00019; 
        10'b0111110010: data <= 17'h1ff75; 
        10'b0111110011: data <= 17'h1ffc4; 
        10'b0111110100: data <= 17'h1ffa6; 
        10'b0111110101: data <= 17'h1ffcc; 
        10'b0111110110: data <= 17'h0005b; 
        10'b0111110111: data <= 17'h0006f; 
        10'b0111111000: data <= 17'h00038; 
        10'b0111111001: data <= 17'h00055; 
        10'b0111111010: data <= 17'h0004b; 
        10'b0111111011: data <= 17'h0000b; 
        10'b0111111100: data <= 17'h1ffa9; 
        10'b0111111101: data <= 17'h1ff48; 
        10'b0111111110: data <= 17'h1ff2b; 
        10'b0111111111: data <= 17'h1fffc; 
        10'b1000000000: data <= 17'h000b9; 
        10'b1000000001: data <= 17'h0002a; 
        10'b1000000010: data <= 17'h1ff6a; 
        10'b1000000011: data <= 17'h1ffa7; 
        10'b1000000100: data <= 17'h000ec; 
        10'b1000000101: data <= 17'h0010a; 
        10'b1000000110: data <= 17'h001c2; 
        10'b1000000111: data <= 17'h00181; 
        10'b1000001000: data <= 17'h000c9; 
        10'b1000001001: data <= 17'h1fec9; 
        10'b1000001010: data <= 17'h1fed9; 
        10'b1000001011: data <= 17'h1fe50; 
        10'b1000001100: data <= 17'h1feff; 
        10'b1000001101: data <= 17'h1fef6; 
        10'b1000001110: data <= 17'h1fe9e; 
        10'b1000001111: data <= 17'h1feed; 
        10'b1000010000: data <= 17'h1ffb8; 
        10'b1000010001: data <= 17'h1ffda; 
        10'b1000010010: data <= 17'h00021; 
        10'b1000010011: data <= 17'h00005; 
        10'b1000010100: data <= 17'h00036; 
        10'b1000010101: data <= 17'h00064; 
        10'b1000010110: data <= 17'h00026; 
        10'b1000010111: data <= 17'h00017; 
        10'b1000011000: data <= 17'h1ff3a; 
        10'b1000011001: data <= 17'h1ff0a; 
        10'b1000011010: data <= 17'h1febb; 
        10'b1000011011: data <= 17'h1fe18; 
        10'b1000011100: data <= 17'h1fdd9; 
        10'b1000011101: data <= 17'h1fdb5; 
        10'b1000011110: data <= 17'h1fd4c; 
        10'b1000011111: data <= 17'h1fd6a; 
        10'b1000100000: data <= 17'h1fdb5; 
        10'b1000100001: data <= 17'h1fea8; 
        10'b1000100010: data <= 17'h1ff9a; 
        10'b1000100011: data <= 17'h00059; 
        10'b1000100100: data <= 17'h1fef5; 
        10'b1000100101: data <= 17'h1ff1a; 
        10'b1000100110: data <= 17'h1fee5; 
        10'b1000100111: data <= 17'h1fe7a; 
        10'b1000101000: data <= 17'h1fe4c; 
        10'b1000101001: data <= 17'h1fe6e; 
        10'b1000101010: data <= 17'h1fe68; 
        10'b1000101011: data <= 17'h1feec; 
        10'b1000101100: data <= 17'h1ffb7; 
        10'b1000101101: data <= 17'h00037; 
        10'b1000101110: data <= 17'h00061; 
        10'b1000101111: data <= 17'h00058; 
        10'b1000110000: data <= 17'h00090; 
        10'b1000110001: data <= 17'h00085; 
        10'b1000110010: data <= 17'h00027; 
        10'b1000110011: data <= 17'h00017; 
        10'b1000110100: data <= 17'h1ff5f; 
        10'b1000110101: data <= 17'h1feed; 
        10'b1000110110: data <= 17'h1fe71; 
        10'b1000110111: data <= 17'h1fd76; 
        10'b1000111000: data <= 17'h1fcfc; 
        10'b1000111001: data <= 17'h1fcce; 
        10'b1000111010: data <= 17'h1fcbf; 
        10'b1000111011: data <= 17'h1fd9e; 
        10'b1000111100: data <= 17'h1fe13; 
        10'b1000111101: data <= 17'h1fdd8; 
        10'b1000111110: data <= 17'h1fea5; 
        10'b1000111111: data <= 17'h1ff4b; 
        10'b1001000000: data <= 17'h1ffc2; 
        10'b1001000001: data <= 17'h1ffdd; 
        10'b1001000010: data <= 17'h1ff71; 
        10'b1001000011: data <= 17'h1fec9; 
        10'b1001000100: data <= 17'h1ff2f; 
        10'b1001000101: data <= 17'h1ff14; 
        10'b1001000110: data <= 17'h1fee3; 
        10'b1001000111: data <= 17'h1ff6e; 
        10'b1001001000: data <= 17'h1ff74; 
        10'b1001001001: data <= 17'h0000a; 
        10'b1001001010: data <= 17'h00022; 
        10'b1001001011: data <= 17'h00060; 
        10'b1001001100: data <= 17'h0001b; 
        10'b1001001101: data <= 17'h0002a; 
        10'b1001001110: data <= 17'h0000b; 
        10'b1001001111: data <= 17'h00013; 
        10'b1001010000: data <= 17'h1fffe; 
        10'b1001010001: data <= 17'h1ff63; 
        10'b1001010010: data <= 17'h1fe77; 
        10'b1001010011: data <= 17'h1fdd9; 
        10'b1001010100: data <= 17'h1fe10; 
        10'b1001010101: data <= 17'h1fdcc; 
        10'b1001010110: data <= 17'h1fe15; 
        10'b1001010111: data <= 17'h1fe93; 
        10'b1001011000: data <= 17'h1fed1; 
        10'b1001011001: data <= 17'h1fee7; 
        10'b1001011010: data <= 17'h1febe; 
        10'b1001011011: data <= 17'h1ff6b; 
        10'b1001011100: data <= 17'h1ff39; 
        10'b1001011101: data <= 17'h00024; 
        10'b1001011110: data <= 17'h1ffc5; 
        10'b1001011111: data <= 17'h0000b; 
        10'b1001100000: data <= 17'h1ffe6; 
        10'b1001100001: data <= 17'h1ff3f; 
        10'b1001100010: data <= 17'h1ff5c; 
        10'b1001100011: data <= 17'h1ffe2; 
        10'b1001100100: data <= 17'h1fffb; 
        10'b1001100101: data <= 17'h0003c; 
        10'b1001100110: data <= 17'h00050; 
        10'b1001100111: data <= 17'h0004d; 
        10'b1001101000: data <= 17'h00045; 
        10'b1001101001: data <= 17'h00051; 
        10'b1001101010: data <= 17'h00020; 
        10'b1001101011: data <= 17'h00058; 
        10'b1001101100: data <= 17'h1ffeb; 
        10'b1001101101: data <= 17'h1ffad; 
        10'b1001101110: data <= 17'h1ff5e; 
        10'b1001101111: data <= 17'h1fef4; 
        10'b1001110000: data <= 17'h1fe96; 
        10'b1001110001: data <= 17'h1ff24; 
        10'b1001110010: data <= 17'h1ff1d; 
        10'b1001110011: data <= 17'h1ff63; 
        10'b1001110100: data <= 17'h1ff5a; 
        10'b1001110101: data <= 17'h1ff72; 
        10'b1001110110: data <= 17'h1ff4e; 
        10'b1001110111: data <= 17'h1ff93; 
        10'b1001111000: data <= 17'h1ff97; 
        10'b1001111001: data <= 17'h00026; 
        10'b1001111010: data <= 17'h000a1; 
        10'b1001111011: data <= 17'h00106; 
        10'b1001111100: data <= 17'h000c9; 
        10'b1001111101: data <= 17'h00084; 
        10'b1001111110: data <= 17'h1ffa9; 
        10'b1001111111: data <= 17'h1ffaa; 
        10'b1010000000: data <= 17'h1fffd; 
        10'b1010000001: data <= 17'h0003a; 
        10'b1010000010: data <= 17'h00009; 
        10'b1010000011: data <= 17'h0002c; 
        10'b1010000100: data <= 17'h0002d; 
        10'b1010000101: data <= 17'h00003; 
        10'b1010000110: data <= 17'h00028; 
        10'b1010000111: data <= 17'h0004f; 
        10'b1010001000: data <= 17'h0002c; 
        10'b1010001001: data <= 17'h00037; 
        10'b1010001010: data <= 17'h1ffaa; 
        10'b1010001011: data <= 17'h1ffa0; 
        10'b1010001100: data <= 17'h1ff7e; 
        10'b1010001101: data <= 17'h0003d; 
        10'b1010001110: data <= 17'h1ff74; 
        10'b1010001111: data <= 17'h00017; 
        10'b1010010000: data <= 17'h1ff6f; 
        10'b1010010001: data <= 17'h1ff8e; 
        10'b1010010010: data <= 17'h1ff91; 
        10'b1010010011: data <= 17'h1fff8; 
        10'b1010010100: data <= 17'h00025; 
        10'b1010010101: data <= 17'h00062; 
        10'b1010010110: data <= 17'h0012e; 
        10'b1010010111: data <= 17'h00126; 
        10'b1010011000: data <= 17'h000fb; 
        10'b1010011001: data <= 17'h00070; 
        10'b1010011010: data <= 17'h1ffd7; 
        10'b1010011011: data <= 17'h00022; 
        10'b1010011100: data <= 17'h00042; 
        10'b1010011101: data <= 17'h0005b; 
        10'b1010011110: data <= 17'h0001e; 
        10'b1010011111: data <= 17'h00071; 
        10'b1010100000: data <= 17'h00056; 
        10'b1010100001: data <= 17'h0007a; 
        10'b1010100010: data <= 17'h0003a; 
        10'b1010100011: data <= 17'h00061; 
        10'b1010100100: data <= 17'h00017; 
        10'b1010100101: data <= 17'h0004a; 
        10'b1010100110: data <= 17'h0001c; 
        10'b1010100111: data <= 17'h1ff76; 
        10'b1010101000: data <= 17'h1ff73; 
        10'b1010101001: data <= 17'h1ffd3; 
        10'b1010101010: data <= 17'h1ff6b; 
        10'b1010101011: data <= 17'h1ffe8; 
        10'b1010101100: data <= 17'h1ff95; 
        10'b1010101101: data <= 17'h1ff9d; 
        10'b1010101110: data <= 17'h1ff4a; 
        10'b1010101111: data <= 17'h1ff34; 
        10'b1010110000: data <= 17'h1ffa8; 
        10'b1010110001: data <= 17'h1ffd2; 
        10'b1010110010: data <= 17'h00010; 
        10'b1010110011: data <= 17'h0009f; 
        10'b1010110100: data <= 17'h00074; 
        10'b1010110101: data <= 17'h1ffd1; 
        10'b1010110110: data <= 17'h1fff2; 
        10'b1010110111: data <= 17'h0003d; 
        10'b1010111000: data <= 17'h00065; 
        10'b1010111001: data <= 17'h00010; 
        10'b1010111010: data <= 17'h0001a; 
        10'b1010111011: data <= 17'h00057; 
        10'b1010111100: data <= 17'h00080; 
        10'b1010111101: data <= 17'h0007c; 
        10'b1010111110: data <= 17'h00072; 
        10'b1010111111: data <= 17'h00019; 
        10'b1011000000: data <= 17'h00072; 
        10'b1011000001: data <= 17'h00005; 
        10'b1011000010: data <= 17'h1ffae; 
        10'b1011000011: data <= 17'h1ff7b; 
        10'b1011000100: data <= 17'h1ff38; 
        10'b1011000101: data <= 17'h1ff2e; 
        10'b1011000110: data <= 17'h1fea7; 
        10'b1011000111: data <= 17'h1fe7a; 
        10'b1011001000: data <= 17'h1fe90; 
        10'b1011001001: data <= 17'h1fe92; 
        10'b1011001010: data <= 17'h1fec9; 
        10'b1011001011: data <= 17'h1feb7; 
        10'b1011001100: data <= 17'h1fe56; 
        10'b1011001101: data <= 17'h1fe1b; 
        10'b1011001110: data <= 17'h1fe4c; 
        10'b1011001111: data <= 17'h1ff11; 
        10'b1011010000: data <= 17'h1ff26; 
        10'b1011010001: data <= 17'h1ffb1; 
        10'b1011010010: data <= 17'h00005; 
        10'b1011010011: data <= 17'h00054; 
        10'b1011010100: data <= 17'h00006; 
        10'b1011010101: data <= 17'h00074; 
        10'b1011010110: data <= 17'h0002e; 
        10'b1011010111: data <= 17'h0002a; 
        10'b1011011000: data <= 17'h0003c; 
        10'b1011011001: data <= 17'h00056; 
        10'b1011011010: data <= 17'h00014; 
        10'b1011011011: data <= 17'h0003a; 
        10'b1011011100: data <= 17'h1fffa; 
        10'b1011011101: data <= 17'h1ffec; 
        10'b1011011110: data <= 17'h00023; 
        10'b1011011111: data <= 17'h00019; 
        10'b1011100000: data <= 17'h1ffe6; 
        10'b1011100001: data <= 17'h1ff87; 
        10'b1011100010: data <= 17'h1fedc; 
        10'b1011100011: data <= 17'h1ff02; 
        10'b1011100100: data <= 17'h1fedd; 
        10'b1011100101: data <= 17'h1fe75; 
        10'b1011100110: data <= 17'h1fe50; 
        10'b1011100111: data <= 17'h1feb0; 
        10'b1011101000: data <= 17'h1fe81; 
        10'b1011101001: data <= 17'h1febb; 
        10'b1011101010: data <= 17'h1fef5; 
        10'b1011101011: data <= 17'h1ff61; 
        10'b1011101100: data <= 17'h1ffc6; 
        10'b1011101101: data <= 17'h00056; 
        10'b1011101110: data <= 17'h00055; 
        10'b1011101111: data <= 17'h0000b; 
        10'b1011110000: data <= 17'h00038; 
        10'b1011110001: data <= 17'h00009; 
        10'b1011110010: data <= 17'h00089; 
        10'b1011110011: data <= 17'h0003c; 
        10'b1011110100: data <= 17'h00053; 
        10'b1011110101: data <= 17'h0000c; 
        10'b1011110110: data <= 17'h00013; 
        10'b1011110111: data <= 17'h00084; 
        10'b1011111000: data <= 17'h00032; 
        10'b1011111001: data <= 17'h0006e; 
        10'b1011111010: data <= 17'h00033; 
        10'b1011111011: data <= 17'h00087; 
        10'b1011111100: data <= 17'h00000; 
        10'b1011111101: data <= 17'h0003a; 
        10'b1011111110: data <= 17'h0001e; 
        10'b1011111111: data <= 17'h1ffed; 
        10'b1100000000: data <= 17'h1fff2; 
        10'b1100000001: data <= 17'h00005; 
        10'b1100000010: data <= 17'h1ffc8; 
        10'b1100000011: data <= 17'h0006b; 
        10'b1100000100: data <= 17'h1ffe5; 
        10'b1100000101: data <= 17'h1ffe1; 
        10'b1100000110: data <= 17'h1fff5; 
        10'b1100000111: data <= 17'h00038; 
        10'b1100001000: data <= 17'h0002b; 
        10'b1100001001: data <= 17'h0002b; 
        10'b1100001010: data <= 17'h0002e; 
        10'b1100001011: data <= 17'h0004e; 
        10'b1100001100: data <= 17'h0004b; 
        10'b1100001101: data <= 17'h00063; 
        10'b1100001110: data <= 17'h00047; 
        10'b1100001111: data <= 17'h0002f; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 12) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 18'h00000; 
        10'b0000000001: data <= 18'h00024; 
        10'b0000000010: data <= 18'h000f2; 
        10'b0000000011: data <= 18'h000f2; 
        10'b0000000100: data <= 18'h00004; 
        10'b0000000101: data <= 18'h00005; 
        10'b0000000110: data <= 18'h000bd; 
        10'b0000000111: data <= 18'h00034; 
        10'b0000001000: data <= 18'h00010; 
        10'b0000001001: data <= 18'h00024; 
        10'b0000001010: data <= 18'h00007; 
        10'b0000001011: data <= 18'h000ae; 
        10'b0000001100: data <= 18'h000e5; 
        10'b0000001101: data <= 18'h00082; 
        10'b0000001110: data <= 18'h000a8; 
        10'b0000001111: data <= 18'h00013; 
        10'b0000010000: data <= 18'h0009e; 
        10'b0000010001: data <= 18'h000d8; 
        10'b0000010010: data <= 18'h0002d; 
        10'b0000010011: data <= 18'h000ae; 
        10'b0000010100: data <= 18'h0000d; 
        10'b0000010101: data <= 18'h00068; 
        10'b0000010110: data <= 18'h000e9; 
        10'b0000010111: data <= 18'h00017; 
        10'b0000011000: data <= 18'h000e9; 
        10'b0000011001: data <= 18'h00025; 
        10'b0000011010: data <= 18'h000ff; 
        10'b0000011011: data <= 18'h00069; 
        10'b0000011100: data <= 18'h00043; 
        10'b0000011101: data <= 18'h00077; 
        10'b0000011110: data <= 18'h3fffe; 
        10'b0000011111: data <= 18'h00014; 
        10'b0000100000: data <= 18'h00074; 
        10'b0000100001: data <= 18'h00119; 
        10'b0000100010: data <= 18'h0003a; 
        10'b0000100011: data <= 18'h3ffd3; 
        10'b0000100100: data <= 18'h0009c; 
        10'b0000100101: data <= 18'h00006; 
        10'b0000100110: data <= 18'h00069; 
        10'b0000100111: data <= 18'h3ffae; 
        10'b0000101000: data <= 18'h00048; 
        10'b0000101001: data <= 18'h3ff8f; 
        10'b0000101010: data <= 18'h00006; 
        10'b0000101011: data <= 18'h0009a; 
        10'b0000101100: data <= 18'h000b6; 
        10'b0000101101: data <= 18'h00035; 
        10'b0000101110: data <= 18'h00003; 
        10'b0000101111: data <= 18'h0002e; 
        10'b0000110000: data <= 18'h000c4; 
        10'b0000110001: data <= 18'h3fffb; 
        10'b0000110010: data <= 18'h3fff9; 
        10'b0000110011: data <= 18'h00010; 
        10'b0000110100: data <= 18'h000ad; 
        10'b0000110101: data <= 18'h000b7; 
        10'b0000110110: data <= 18'h0002b; 
        10'b0000110111: data <= 18'h000b7; 
        10'b0000111000: data <= 18'h000d2; 
        10'b0000111001: data <= 18'h00088; 
        10'b0000111010: data <= 18'h000cf; 
        10'b0000111011: data <= 18'h000d4; 
        10'b0000111100: data <= 18'h000c9; 
        10'b0000111101: data <= 18'h000b3; 
        10'b0000111110: data <= 18'h000ee; 
        10'b0000111111: data <= 18'h3ffb4; 
        10'b0001000000: data <= 18'h3ffae; 
        10'b0001000001: data <= 18'h0002b; 
        10'b0001000010: data <= 18'h3ffe4; 
        10'b0001000011: data <= 18'h3ff73; 
        10'b0001000100: data <= 18'h3fdde; 
        10'b0001000101: data <= 18'h3ff23; 
        10'b0001000110: data <= 18'h3fef8; 
        10'b0001000111: data <= 18'h3fe8a; 
        10'b0001001000: data <= 18'h3feef; 
        10'b0001001001: data <= 18'h3ffca; 
        10'b0001001010: data <= 18'h00044; 
        10'b0001001011: data <= 18'h000c0; 
        10'b0001001100: data <= 18'h000fa; 
        10'b0001001101: data <= 18'h00090; 
        10'b0001001110: data <= 18'h000eb; 
        10'b0001001111: data <= 18'h0003f; 
        10'b0001010000: data <= 18'h00059; 
        10'b0001010001: data <= 18'h0009f; 
        10'b0001010010: data <= 18'h0000a; 
        10'b0001010011: data <= 18'h0006f; 
        10'b0001010100: data <= 18'h000d4; 
        10'b0001010101: data <= 18'h000be; 
        10'b0001010110: data <= 18'h00049; 
        10'b0001010111: data <= 18'h00078; 
        10'b0001011000: data <= 18'h0007c; 
        10'b0001011001: data <= 18'h00002; 
        10'b0001011010: data <= 18'h0009f; 
        10'b0001011011: data <= 18'h3ff73; 
        10'b0001011100: data <= 18'h3ff32; 
        10'b0001011101: data <= 18'h3ff90; 
        10'b0001011110: data <= 18'h3fe2a; 
        10'b0001011111: data <= 18'h3fdd4; 
        10'b0001100000: data <= 18'h3fc89; 
        10'b0001100001: data <= 18'h3fcb2; 
        10'b0001100010: data <= 18'h3fcda; 
        10'b0001100011: data <= 18'h3fc2e; 
        10'b0001100100: data <= 18'h3fd73; 
        10'b0001100101: data <= 18'h3feba; 
        10'b0001100110: data <= 18'h00030; 
        10'b0001100111: data <= 18'h00069; 
        10'b0001101000: data <= 18'h000bd; 
        10'b0001101001: data <= 18'h00117; 
        10'b0001101010: data <= 18'h00049; 
        10'b0001101011: data <= 18'h0004b; 
        10'b0001101100: data <= 18'h0010f; 
        10'b0001101101: data <= 18'h00105; 
        10'b0001101110: data <= 18'h00051; 
        10'b0001101111: data <= 18'h00099; 
        10'b0001110000: data <= 18'h00108; 
        10'b0001110001: data <= 18'h000af; 
        10'b0001110010: data <= 18'h000c5; 
        10'b0001110011: data <= 18'h000bf; 
        10'b0001110100: data <= 18'h00072; 
        10'b0001110101: data <= 18'h000d8; 
        10'b0001110110: data <= 18'h3ff5e; 
        10'b0001110111: data <= 18'h3ffdc; 
        10'b0001111000: data <= 18'h3feb5; 
        10'b0001111001: data <= 18'h3fee8; 
        10'b0001111010: data <= 18'h3fce5; 
        10'b0001111011: data <= 18'h3fd0b; 
        10'b0001111100: data <= 18'h3fbf5; 
        10'b0001111101: data <= 18'h3fca5; 
        10'b0001111110: data <= 18'h3fbe1; 
        10'b0001111111: data <= 18'h3fc79; 
        10'b0010000000: data <= 18'h3fe49; 
        10'b0010000001: data <= 18'h3fe7a; 
        10'b0010000010: data <= 18'h3ff17; 
        10'b0010000011: data <= 18'h000e0; 
        10'b0010000100: data <= 18'h00135; 
        10'b0010000101: data <= 18'h00161; 
        10'b0010000110: data <= 18'h00150; 
        10'b0010000111: data <= 18'h001be; 
        10'b0010001000: data <= 18'h0007c; 
        10'b0010001001: data <= 18'h000fb; 
        10'b0010001010: data <= 18'h00040; 
        10'b0010001011: data <= 18'h00029; 
        10'b0010001100: data <= 18'h0010c; 
        10'b0010001101: data <= 18'h0004b; 
        10'b0010001110: data <= 18'h000bd; 
        10'b0010001111: data <= 18'h0003e; 
        10'b0010010000: data <= 18'h000ae; 
        10'b0010010001: data <= 18'h00023; 
        10'b0010010010: data <= 18'h0007b; 
        10'b0010010011: data <= 18'h3ff6b; 
        10'b0010010100: data <= 18'h00028; 
        10'b0010010101: data <= 18'h3ff54; 
        10'b0010010110: data <= 18'h3fdba; 
        10'b0010010111: data <= 18'h3fe7f; 
        10'b0010011000: data <= 18'h3fd6b; 
        10'b0010011001: data <= 18'h3fccc; 
        10'b0010011010: data <= 18'h3fdc2; 
        10'b0010011011: data <= 18'h3fe26; 
        10'b0010011100: data <= 18'h3ffb1; 
        10'b0010011101: data <= 18'h00049; 
        10'b0010011110: data <= 18'h3ff8f; 
        10'b0010011111: data <= 18'h000bf; 
        10'b0010100000: data <= 18'h000ea; 
        10'b0010100001: data <= 18'h0013d; 
        10'b0010100010: data <= 18'h002e2; 
        10'b0010100011: data <= 18'h00341; 
        10'b0010100100: data <= 18'h001c5; 
        10'b0010100101: data <= 18'h3ffd4; 
        10'b0010100110: data <= 18'h0004a; 
        10'b0010100111: data <= 18'h0002d; 
        10'b0010101000: data <= 18'h000f9; 
        10'b0010101001: data <= 18'h00113; 
        10'b0010101010: data <= 18'h00052; 
        10'b0010101011: data <= 18'h000d9; 
        10'b0010101100: data <= 18'h000ec; 
        10'b0010101101: data <= 18'h000c2; 
        10'b0010101110: data <= 18'h000c0; 
        10'b0010101111: data <= 18'h3fff1; 
        10'b0010110000: data <= 18'h3ffd5; 
        10'b0010110001: data <= 18'h3ff1c; 
        10'b0010110010: data <= 18'h3fe32; 
        10'b0010110011: data <= 18'h3fcd4; 
        10'b0010110100: data <= 18'h3fb32; 
        10'b0010110101: data <= 18'h3fa52; 
        10'b0010110110: data <= 18'h3fa11; 
        10'b0010110111: data <= 18'h3fad9; 
        10'b0010111000: data <= 18'h3fab9; 
        10'b0010111001: data <= 18'h3fce8; 
        10'b0010111010: data <= 18'h3fcce; 
        10'b0010111011: data <= 18'h3fe90; 
        10'b0010111100: data <= 18'h3ff0e; 
        10'b0010111101: data <= 18'h3ffed; 
        10'b0010111110: data <= 18'h00420; 
        10'b0010111111: data <= 18'h00456; 
        10'b0011000000: data <= 18'h001ab; 
        10'b0011000001: data <= 18'h0014f; 
        10'b0011000010: data <= 18'h000ef; 
        10'b0011000011: data <= 18'h0000a; 
        10'b0011000100: data <= 18'h00076; 
        10'b0011000101: data <= 18'h0003e; 
        10'b0011000110: data <= 18'h00055; 
        10'b0011000111: data <= 18'h00096; 
        10'b0011001000: data <= 18'h00056; 
        10'b0011001001: data <= 18'h000c8; 
        10'b0011001010: data <= 18'h3ff84; 
        10'b0011001011: data <= 18'h3ffe9; 
        10'b0011001100: data <= 18'h3ff77; 
        10'b0011001101: data <= 18'h3fec8; 
        10'b0011001110: data <= 18'h3fcec; 
        10'b0011001111: data <= 18'h3fb33; 
        10'b0011010000: data <= 18'h3f9c4; 
        10'b0011010001: data <= 18'h3fb98; 
        10'b0011010010: data <= 18'h3fa7d; 
        10'b0011010011: data <= 18'h3fa73; 
        10'b0011010100: data <= 18'h3fa4a; 
        10'b0011010101: data <= 18'h3fc5c; 
        10'b0011010110: data <= 18'h3fc45; 
        10'b0011010111: data <= 18'h3fd67; 
        10'b0011011000: data <= 18'h3fd00; 
        10'b0011011001: data <= 18'h3fea2; 
        10'b0011011010: data <= 18'h0028c; 
        10'b0011011011: data <= 18'h00373; 
        10'b0011011100: data <= 18'h001d7; 
        10'b0011011101: data <= 18'h00109; 
        10'b0011011110: data <= 18'h000f9; 
        10'b0011011111: data <= 18'h00094; 
        10'b0011100000: data <= 18'h000f0; 
        10'b0011100001: data <= 18'h000c9; 
        10'b0011100010: data <= 18'h00109; 
        10'b0011100011: data <= 18'h00033; 
        10'b0011100100: data <= 18'h00050; 
        10'b0011100101: data <= 18'h0006d; 
        10'b0011100110: data <= 18'h00049; 
        10'b0011100111: data <= 18'h3ffc0; 
        10'b0011101000: data <= 18'h3fdae; 
        10'b0011101001: data <= 18'h3fed2; 
        10'b0011101010: data <= 18'h3fe75; 
        10'b0011101011: data <= 18'h3fce6; 
        10'b0011101100: data <= 18'h3fb75; 
        10'b0011101101: data <= 18'h3fd19; 
        10'b0011101110: data <= 18'h3f96b; 
        10'b0011101111: data <= 18'h3f93d; 
        10'b0011110000: data <= 18'h3fabe; 
        10'b0011110001: data <= 18'h3fcb5; 
        10'b0011110010: data <= 18'h3fd0c; 
        10'b0011110011: data <= 18'h3ff12; 
        10'b0011110100: data <= 18'h3fe32; 
        10'b0011110101: data <= 18'h3fe3a; 
        10'b0011110110: data <= 18'h0012d; 
        10'b0011110111: data <= 18'h001cf; 
        10'b0011111000: data <= 18'h00161; 
        10'b0011111001: data <= 18'h00046; 
        10'b0011111010: data <= 18'h0005f; 
        10'b0011111011: data <= 18'h000ad; 
        10'b0011111100: data <= 18'h0011d; 
        10'b0011111101: data <= 18'h000f0; 
        10'b0011111110: data <= 18'h000e0; 
        10'b0011111111: data <= 18'h0002f; 
        10'b0100000000: data <= 18'h3ff6b; 
        10'b0100000001: data <= 18'h00004; 
        10'b0100000010: data <= 18'h3fe92; 
        10'b0100000011: data <= 18'h3fef9; 
        10'b0100000100: data <= 18'h3ff55; 
        10'b0100000101: data <= 18'h3ffc8; 
        10'b0100000110: data <= 18'h3ff35; 
        10'b0100000111: data <= 18'h3ff0b; 
        10'b0100001000: data <= 18'h3ff04; 
        10'b0100001001: data <= 18'h3fd61; 
        10'b0100001010: data <= 18'h3f683; 
        10'b0100001011: data <= 18'h3f8e7; 
        10'b0100001100: data <= 18'h3fe47; 
        10'b0100001101: data <= 18'h3feba; 
        10'b0100001110: data <= 18'h3ff9b; 
        10'b0100001111: data <= 18'h00036; 
        10'b0100010000: data <= 18'h3ff01; 
        10'b0100010001: data <= 18'h3ff07; 
        10'b0100010010: data <= 18'h0007e; 
        10'b0100010011: data <= 18'h0001d; 
        10'b0100010100: data <= 18'h3fedf; 
        10'b0100010101: data <= 18'h3fed3; 
        10'b0100010110: data <= 18'h3ff7e; 
        10'b0100010111: data <= 18'h000c1; 
        10'b0100011000: data <= 18'h00098; 
        10'b0100011001: data <= 18'h0006c; 
        10'b0100011010: data <= 18'h0006d; 
        10'b0100011011: data <= 18'h0001e; 
        10'b0100011100: data <= 18'h00071; 
        10'b0100011101: data <= 18'h3feb9; 
        10'b0100011110: data <= 18'h3fde3; 
        10'b0100011111: data <= 18'h3fef9; 
        10'b0100100000: data <= 18'h0004e; 
        10'b0100100001: data <= 18'h002b4; 
        10'b0100100010: data <= 18'h001a3; 
        10'b0100100011: data <= 18'h00139; 
        10'b0100100100: data <= 18'h00177; 
        10'b0100100101: data <= 18'h3fc5f; 
        10'b0100100110: data <= 18'h3f5fb; 
        10'b0100100111: data <= 18'h3fcf2; 
        10'b0100101000: data <= 18'h00059; 
        10'b0100101001: data <= 18'h3ff8d; 
        10'b0100101010: data <= 18'h3ffa8; 
        10'b0100101011: data <= 18'h0005b; 
        10'b0100101100: data <= 18'h3fe00; 
        10'b0100101101: data <= 18'h3feae; 
        10'b0100101110: data <= 18'h3ffc0; 
        10'b0100101111: data <= 18'h3fdd3; 
        10'b0100110000: data <= 18'h3fec4; 
        10'b0100110001: data <= 18'h3ff38; 
        10'b0100110010: data <= 18'h000a0; 
        10'b0100110011: data <= 18'h00108; 
        10'b0100110100: data <= 18'h000b2; 
        10'b0100110101: data <= 18'h000b9; 
        10'b0100110110: data <= 18'h0009c; 
        10'b0100110111: data <= 18'h3ff9e; 
        10'b0100111000: data <= 18'h3ffdc; 
        10'b0100111001: data <= 18'h3ff49; 
        10'b0100111010: data <= 18'h3ff3f; 
        10'b0100111011: data <= 18'h000a4; 
        10'b0100111100: data <= 18'h0020c; 
        10'b0100111101: data <= 18'h00372; 
        10'b0100111110: data <= 18'h004c0; 
        10'b0100111111: data <= 18'h00306; 
        10'b0101000000: data <= 18'h00369; 
        10'b0101000001: data <= 18'h3fa71; 
        10'b0101000010: data <= 18'h3f874; 
        10'b0101000011: data <= 18'h000fb; 
        10'b0101000100: data <= 18'h003e7; 
        10'b0101000101: data <= 18'h000a8; 
        10'b0101000110: data <= 18'h3ffc6; 
        10'b0101000111: data <= 18'h3ff60; 
        10'b0101001000: data <= 18'h3fdde; 
        10'b0101001001: data <= 18'h3fe2d; 
        10'b0101001010: data <= 18'h3ff12; 
        10'b0101001011: data <= 18'h3fe50; 
        10'b0101001100: data <= 18'h3fe20; 
        10'b0101001101: data <= 18'h3ffe5; 
        10'b0101001110: data <= 18'h3fff0; 
        10'b0101001111: data <= 18'h00042; 
        10'b0101010000: data <= 18'h000c6; 
        10'b0101010001: data <= 18'h000ae; 
        10'b0101010010: data <= 18'h00052; 
        10'b0101010011: data <= 18'h00077; 
        10'b0101010100: data <= 18'h3fff4; 
        10'b0101010101: data <= 18'h3ff4d; 
        10'b0101010110: data <= 18'h00202; 
        10'b0101010111: data <= 18'h0034f; 
        10'b0101011000: data <= 18'h00520; 
        10'b0101011001: data <= 18'h0047d; 
        10'b0101011010: data <= 18'h00778; 
        10'b0101011011: data <= 18'h00876; 
        10'b0101011100: data <= 18'h007ff; 
        10'b0101011101: data <= 18'h3ffde; 
        10'b0101011110: data <= 18'h3fc06; 
        10'b0101011111: data <= 18'h00321; 
        10'b0101100000: data <= 18'h00515; 
        10'b0101100001: data <= 18'h00094; 
        10'b0101100010: data <= 18'h00037; 
        10'b0101100011: data <= 18'h000b2; 
        10'b0101100100: data <= 18'h3ffe1; 
        10'b0101100101: data <= 18'h00026; 
        10'b0101100110: data <= 18'h3ffc6; 
        10'b0101100111: data <= 18'h3fee1; 
        10'b0101101000: data <= 18'h3ff00; 
        10'b0101101001: data <= 18'h3ffb8; 
        10'b0101101010: data <= 18'h0011b; 
        10'b0101101011: data <= 18'h000a3; 
        10'b0101101100: data <= 18'h0001f; 
        10'b0101101101: data <= 18'h000ba; 
        10'b0101101110: data <= 18'h0001a; 
        10'b0101101111: data <= 18'h0004e; 
        10'b0101110000: data <= 18'h000dc; 
        10'b0101110001: data <= 18'h0026c; 
        10'b0101110010: data <= 18'h004ed; 
        10'b0101110011: data <= 18'h005b7; 
        10'b0101110100: data <= 18'h00692; 
        10'b0101110101: data <= 18'h0057d; 
        10'b0101110110: data <= 18'h00668; 
        10'b0101110111: data <= 18'h00a71; 
        10'b0101111000: data <= 18'h007ea; 
        10'b0101111001: data <= 18'h0001e; 
        10'b0101111010: data <= 18'h3fee0; 
        10'b0101111011: data <= 18'h003ab; 
        10'b0101111100: data <= 18'h003c4; 
        10'b0101111101: data <= 18'h0042f; 
        10'b0101111110: data <= 18'h002e3; 
        10'b0101111111: data <= 18'h0014c; 
        10'b0110000000: data <= 18'h002e4; 
        10'b0110000001: data <= 18'h00220; 
        10'b0110000010: data <= 18'h00103; 
        10'b0110000011: data <= 18'h3ff69; 
        10'b0110000100: data <= 18'h3ff7b; 
        10'b0110000101: data <= 18'h0000f; 
        10'b0110000110: data <= 18'h000e3; 
        10'b0110000111: data <= 18'h000a2; 
        10'b0110001000: data <= 18'h0001d; 
        10'b0110001001: data <= 18'h000e8; 
        10'b0110001010: data <= 18'h00013; 
        10'b0110001011: data <= 18'h00111; 
        10'b0110001100: data <= 18'h00225; 
        10'b0110001101: data <= 18'h00450; 
        10'b0110001110: data <= 18'h005ff; 
        10'b0110001111: data <= 18'h00690; 
        10'b0110010000: data <= 18'h004e7; 
        10'b0110010001: data <= 18'h004b0; 
        10'b0110010010: data <= 18'h005a6; 
        10'b0110010011: data <= 18'h006d8; 
        10'b0110010100: data <= 18'h004fc; 
        10'b0110010101: data <= 18'h0006a; 
        10'b0110010110: data <= 18'h3ff46; 
        10'b0110010111: data <= 18'h00153; 
        10'b0110011000: data <= 18'h00432; 
        10'b0110011001: data <= 18'h006e5; 
        10'b0110011010: data <= 18'h004af; 
        10'b0110011011: data <= 18'h0044e; 
        10'b0110011100: data <= 18'h00267; 
        10'b0110011101: data <= 18'h0019e; 
        10'b0110011110: data <= 18'h00086; 
        10'b0110011111: data <= 18'h0004c; 
        10'b0110100000: data <= 18'h3ffd4; 
        10'b0110100001: data <= 18'h0004a; 
        10'b0110100010: data <= 18'h0008a; 
        10'b0110100011: data <= 18'h00041; 
        10'b0110100100: data <= 18'h000c0; 
        10'b0110100101: data <= 18'h00113; 
        10'b0110100110: data <= 18'h000b0; 
        10'b0110100111: data <= 18'h000e3; 
        10'b0110101000: data <= 18'h001f0; 
        10'b0110101001: data <= 18'h00232; 
        10'b0110101010: data <= 18'h0036a; 
        10'b0110101011: data <= 18'h00325; 
        10'b0110101100: data <= 18'h0050f; 
        10'b0110101101: data <= 18'h00459; 
        10'b0110101110: data <= 18'h00306; 
        10'b0110101111: data <= 18'h00232; 
        10'b0110110000: data <= 18'h00298; 
        10'b0110110001: data <= 18'h00083; 
        10'b0110110010: data <= 18'h00215; 
        10'b0110110011: data <= 18'h002ea; 
        10'b0110110100: data <= 18'h0060c; 
        10'b0110110101: data <= 18'h0055f; 
        10'b0110110110: data <= 18'h003d7; 
        10'b0110110111: data <= 18'h00246; 
        10'b0110111000: data <= 18'h3ff63; 
        10'b0110111001: data <= 18'h000d8; 
        10'b0110111010: data <= 18'h00187; 
        10'b0110111011: data <= 18'h00029; 
        10'b0110111100: data <= 18'h3ff15; 
        10'b0110111101: data <= 18'h0007c; 
        10'b0110111110: data <= 18'h00020; 
        10'b0110111111: data <= 18'h0004e; 
        10'b0111000000: data <= 18'h00055; 
        10'b0111000001: data <= 18'h00002; 
        10'b0111000010: data <= 18'h0000a; 
        10'b0111000011: data <= 18'h3ffde; 
        10'b0111000100: data <= 18'h00087; 
        10'b0111000101: data <= 18'h0014c; 
        10'b0111000110: data <= 18'h0021d; 
        10'b0111000111: data <= 18'h003b1; 
        10'b0111001000: data <= 18'h0055f; 
        10'b0111001001: data <= 18'h003d4; 
        10'b0111001010: data <= 18'h00106; 
        10'b0111001011: data <= 18'h3ffdc; 
        10'b0111001100: data <= 18'h0010d; 
        10'b0111001101: data <= 18'h00150; 
        10'b0111001110: data <= 18'h004ee; 
        10'b0111001111: data <= 18'h006d1; 
        10'b0111010000: data <= 18'h00705; 
        10'b0111010001: data <= 18'h005d5; 
        10'b0111010010: data <= 18'h003f3; 
        10'b0111010011: data <= 18'h0007f; 
        10'b0111010100: data <= 18'h001a8; 
        10'b0111010101: data <= 18'h0025a; 
        10'b0111010110: data <= 18'h0008d; 
        10'b0111010111: data <= 18'h3ff9d; 
        10'b0111011000: data <= 18'h3ffe5; 
        10'b0111011001: data <= 18'h0003b; 
        10'b0111011010: data <= 18'h0006d; 
        10'b0111011011: data <= 18'h00072; 
        10'b0111011100: data <= 18'h00065; 
        10'b0111011101: data <= 18'h00067; 
        10'b0111011110: data <= 18'h000ce; 
        10'b0111011111: data <= 18'h3fffd; 
        10'b0111100000: data <= 18'h3ff70; 
        10'b0111100001: data <= 18'h3fed7; 
        10'b0111100010: data <= 18'h000b0; 
        10'b0111100011: data <= 18'h002ed; 
        10'b0111100100: data <= 18'h005a5; 
        10'b0111100101: data <= 18'h004e4; 
        10'b0111100110: data <= 18'h001c6; 
        10'b0111100111: data <= 18'h00165; 
        10'b0111101000: data <= 18'h00205; 
        10'b0111101001: data <= 18'h004d7; 
        10'b0111101010: data <= 18'h007ff; 
        10'b0111101011: data <= 18'h00654; 
        10'b0111101100: data <= 18'h0054b; 
        10'b0111101101: data <= 18'h001a3; 
        10'b0111101110: data <= 18'h00041; 
        10'b0111101111: data <= 18'h3fe3a; 
        10'b0111110000: data <= 18'h00088; 
        10'b0111110001: data <= 18'h00032; 
        10'b0111110010: data <= 18'h3feeb; 
        10'b0111110011: data <= 18'h3ff89; 
        10'b0111110100: data <= 18'h3ff4b; 
        10'b0111110101: data <= 18'h3ff99; 
        10'b0111110110: data <= 18'h000b6; 
        10'b0111110111: data <= 18'h000df; 
        10'b0111111000: data <= 18'h00070; 
        10'b0111111001: data <= 18'h000ab; 
        10'b0111111010: data <= 18'h00096; 
        10'b0111111011: data <= 18'h00016; 
        10'b0111111100: data <= 18'h3ff52; 
        10'b0111111101: data <= 18'h3fe91; 
        10'b0111111110: data <= 18'h3fe56; 
        10'b0111111111: data <= 18'h3fff8; 
        10'b1000000000: data <= 18'h00172; 
        10'b1000000001: data <= 18'h00054; 
        10'b1000000010: data <= 18'h3fed3; 
        10'b1000000011: data <= 18'h3ff4e; 
        10'b1000000100: data <= 18'h001d8; 
        10'b1000000101: data <= 18'h00215; 
        10'b1000000110: data <= 18'h00384; 
        10'b1000000111: data <= 18'h00302; 
        10'b1000001000: data <= 18'h00192; 
        10'b1000001001: data <= 18'h3fd91; 
        10'b1000001010: data <= 18'h3fdb2; 
        10'b1000001011: data <= 18'h3fc9f; 
        10'b1000001100: data <= 18'h3fdff; 
        10'b1000001101: data <= 18'h3fdec; 
        10'b1000001110: data <= 18'h3fd3b; 
        10'b1000001111: data <= 18'h3fddb; 
        10'b1000010000: data <= 18'h3ff71; 
        10'b1000010001: data <= 18'h3ffb4; 
        10'b1000010010: data <= 18'h00042; 
        10'b1000010011: data <= 18'h00009; 
        10'b1000010100: data <= 18'h0006c; 
        10'b1000010101: data <= 18'h000c8; 
        10'b1000010110: data <= 18'h0004c; 
        10'b1000010111: data <= 18'h0002e; 
        10'b1000011000: data <= 18'h3fe74; 
        10'b1000011001: data <= 18'h3fe14; 
        10'b1000011010: data <= 18'h3fd76; 
        10'b1000011011: data <= 18'h3fc30; 
        10'b1000011100: data <= 18'h3fbb3; 
        10'b1000011101: data <= 18'h3fb6a; 
        10'b1000011110: data <= 18'h3fa97; 
        10'b1000011111: data <= 18'h3fad3; 
        10'b1000100000: data <= 18'h3fb6b; 
        10'b1000100001: data <= 18'h3fd50; 
        10'b1000100010: data <= 18'h3ff34; 
        10'b1000100011: data <= 18'h000b3; 
        10'b1000100100: data <= 18'h3fdeb; 
        10'b1000100101: data <= 18'h3fe35; 
        10'b1000100110: data <= 18'h3fdcb; 
        10'b1000100111: data <= 18'h3fcf4; 
        10'b1000101000: data <= 18'h3fc98; 
        10'b1000101001: data <= 18'h3fcdd; 
        10'b1000101010: data <= 18'h3fccf; 
        10'b1000101011: data <= 18'h3fdd8; 
        10'b1000101100: data <= 18'h3ff6e; 
        10'b1000101101: data <= 18'h0006d; 
        10'b1000101110: data <= 18'h000c1; 
        10'b1000101111: data <= 18'h000b1; 
        10'b1000110000: data <= 18'h00120; 
        10'b1000110001: data <= 18'h0010a; 
        10'b1000110010: data <= 18'h0004d; 
        10'b1000110011: data <= 18'h0002e; 
        10'b1000110100: data <= 18'h3febf; 
        10'b1000110101: data <= 18'h3fdda; 
        10'b1000110110: data <= 18'h3fce1; 
        10'b1000110111: data <= 18'h3faec; 
        10'b1000111000: data <= 18'h3f9f7; 
        10'b1000111001: data <= 18'h3f99b; 
        10'b1000111010: data <= 18'h3f97d; 
        10'b1000111011: data <= 18'h3fb3c; 
        10'b1000111100: data <= 18'h3fc25; 
        10'b1000111101: data <= 18'h3fbb1; 
        10'b1000111110: data <= 18'h3fd4b; 
        10'b1000111111: data <= 18'h3fe97; 
        10'b1001000000: data <= 18'h3ff83; 
        10'b1001000001: data <= 18'h3ffba; 
        10'b1001000010: data <= 18'h3fee1; 
        10'b1001000011: data <= 18'h3fd93; 
        10'b1001000100: data <= 18'h3fe5e; 
        10'b1001000101: data <= 18'h3fe27; 
        10'b1001000110: data <= 18'h3fdc6; 
        10'b1001000111: data <= 18'h3fedc; 
        10'b1001001000: data <= 18'h3fee7; 
        10'b1001001001: data <= 18'h00015; 
        10'b1001001010: data <= 18'h00044; 
        10'b1001001011: data <= 18'h000c0; 
        10'b1001001100: data <= 18'h00035; 
        10'b1001001101: data <= 18'h00054; 
        10'b1001001110: data <= 18'h00016; 
        10'b1001001111: data <= 18'h00026; 
        10'b1001010000: data <= 18'h3fffd; 
        10'b1001010001: data <= 18'h3fec7; 
        10'b1001010010: data <= 18'h3fced; 
        10'b1001010011: data <= 18'h3fbb2; 
        10'b1001010100: data <= 18'h3fc20; 
        10'b1001010101: data <= 18'h3fb98; 
        10'b1001010110: data <= 18'h3fc2a; 
        10'b1001010111: data <= 18'h3fd26; 
        10'b1001011000: data <= 18'h3fda1; 
        10'b1001011001: data <= 18'h3fdce; 
        10'b1001011010: data <= 18'h3fd7c; 
        10'b1001011011: data <= 18'h3fed6; 
        10'b1001011100: data <= 18'h3fe73; 
        10'b1001011101: data <= 18'h00048; 
        10'b1001011110: data <= 18'h3ff8a; 
        10'b1001011111: data <= 18'h00015; 
        10'b1001100000: data <= 18'h3ffcc; 
        10'b1001100001: data <= 18'h3fe7e; 
        10'b1001100010: data <= 18'h3feb9; 
        10'b1001100011: data <= 18'h3ffc4; 
        10'b1001100100: data <= 18'h3fff5; 
        10'b1001100101: data <= 18'h00077; 
        10'b1001100110: data <= 18'h000a0; 
        10'b1001100111: data <= 18'h0009a; 
        10'b1001101000: data <= 18'h0008b; 
        10'b1001101001: data <= 18'h000a1; 
        10'b1001101010: data <= 18'h00040; 
        10'b1001101011: data <= 18'h000b1; 
        10'b1001101100: data <= 18'h3ffd6; 
        10'b1001101101: data <= 18'h3ff59; 
        10'b1001101110: data <= 18'h3febb; 
        10'b1001101111: data <= 18'h3fde8; 
        10'b1001110000: data <= 18'h3fd2c; 
        10'b1001110001: data <= 18'h3fe48; 
        10'b1001110010: data <= 18'h3fe3b; 
        10'b1001110011: data <= 18'h3fec6; 
        10'b1001110100: data <= 18'h3feb4; 
        10'b1001110101: data <= 18'h3fee3; 
        10'b1001110110: data <= 18'h3fe9c; 
        10'b1001110111: data <= 18'h3ff26; 
        10'b1001111000: data <= 18'h3ff2e; 
        10'b1001111001: data <= 18'h0004b; 
        10'b1001111010: data <= 18'h00141; 
        10'b1001111011: data <= 18'h0020c; 
        10'b1001111100: data <= 18'h00192; 
        10'b1001111101: data <= 18'h00108; 
        10'b1001111110: data <= 18'h3ff52; 
        10'b1001111111: data <= 18'h3ff54; 
        10'b1010000000: data <= 18'h3fffa; 
        10'b1010000001: data <= 18'h00073; 
        10'b1010000010: data <= 18'h00012; 
        10'b1010000011: data <= 18'h00058; 
        10'b1010000100: data <= 18'h0005a; 
        10'b1010000101: data <= 18'h00006; 
        10'b1010000110: data <= 18'h00050; 
        10'b1010000111: data <= 18'h0009d; 
        10'b1010001000: data <= 18'h00059; 
        10'b1010001001: data <= 18'h0006d; 
        10'b1010001010: data <= 18'h3ff53; 
        10'b1010001011: data <= 18'h3ff40; 
        10'b1010001100: data <= 18'h3fefc; 
        10'b1010001101: data <= 18'h00079; 
        10'b1010001110: data <= 18'h3fee8; 
        10'b1010001111: data <= 18'h0002d; 
        10'b1010010000: data <= 18'h3fede; 
        10'b1010010001: data <= 18'h3ff1d; 
        10'b1010010010: data <= 18'h3ff22; 
        10'b1010010011: data <= 18'h3fff0; 
        10'b1010010100: data <= 18'h0004a; 
        10'b1010010101: data <= 18'h000c4; 
        10'b1010010110: data <= 18'h0025b; 
        10'b1010010111: data <= 18'h0024c; 
        10'b1010011000: data <= 18'h001f6; 
        10'b1010011001: data <= 18'h000df; 
        10'b1010011010: data <= 18'h3ffad; 
        10'b1010011011: data <= 18'h00044; 
        10'b1010011100: data <= 18'h00085; 
        10'b1010011101: data <= 18'h000b6; 
        10'b1010011110: data <= 18'h0003b; 
        10'b1010011111: data <= 18'h000e3; 
        10'b1010100000: data <= 18'h000ab; 
        10'b1010100001: data <= 18'h000f5; 
        10'b1010100010: data <= 18'h00074; 
        10'b1010100011: data <= 18'h000c2; 
        10'b1010100100: data <= 18'h0002e; 
        10'b1010100101: data <= 18'h00095; 
        10'b1010100110: data <= 18'h00038; 
        10'b1010100111: data <= 18'h3feec; 
        10'b1010101000: data <= 18'h3fee7; 
        10'b1010101001: data <= 18'h3ffa6; 
        10'b1010101010: data <= 18'h3fed6; 
        10'b1010101011: data <= 18'h3ffcf; 
        10'b1010101100: data <= 18'h3ff29; 
        10'b1010101101: data <= 18'h3ff3a; 
        10'b1010101110: data <= 18'h3fe94; 
        10'b1010101111: data <= 18'h3fe68; 
        10'b1010110000: data <= 18'h3ff50; 
        10'b1010110001: data <= 18'h3ffa4; 
        10'b1010110010: data <= 18'h00020; 
        10'b1010110011: data <= 18'h0013d; 
        10'b1010110100: data <= 18'h000e7; 
        10'b1010110101: data <= 18'h3ffa1; 
        10'b1010110110: data <= 18'h3ffe5; 
        10'b1010110111: data <= 18'h0007a; 
        10'b1010111000: data <= 18'h000ca; 
        10'b1010111001: data <= 18'h00020; 
        10'b1010111010: data <= 18'h00034; 
        10'b1010111011: data <= 18'h000ae; 
        10'b1010111100: data <= 18'h00100; 
        10'b1010111101: data <= 18'h000f8; 
        10'b1010111110: data <= 18'h000e3; 
        10'b1010111111: data <= 18'h00033; 
        10'b1011000000: data <= 18'h000e4; 
        10'b1011000001: data <= 18'h0000b; 
        10'b1011000010: data <= 18'h3ff5d; 
        10'b1011000011: data <= 18'h3fef6; 
        10'b1011000100: data <= 18'h3fe70; 
        10'b1011000101: data <= 18'h3fe5b; 
        10'b1011000110: data <= 18'h3fd4d; 
        10'b1011000111: data <= 18'h3fcf5; 
        10'b1011001000: data <= 18'h3fd20; 
        10'b1011001001: data <= 18'h3fd24; 
        10'b1011001010: data <= 18'h3fd92; 
        10'b1011001011: data <= 18'h3fd6e; 
        10'b1011001100: data <= 18'h3fcac; 
        10'b1011001101: data <= 18'h3fc35; 
        10'b1011001110: data <= 18'h3fc98; 
        10'b1011001111: data <= 18'h3fe22; 
        10'b1011010000: data <= 18'h3fe4b; 
        10'b1011010001: data <= 18'h3ff62; 
        10'b1011010010: data <= 18'h0000a; 
        10'b1011010011: data <= 18'h000a7; 
        10'b1011010100: data <= 18'h0000c; 
        10'b1011010101: data <= 18'h000e8; 
        10'b1011010110: data <= 18'h0005d; 
        10'b1011010111: data <= 18'h00054; 
        10'b1011011000: data <= 18'h00078; 
        10'b1011011001: data <= 18'h000ad; 
        10'b1011011010: data <= 18'h00027; 
        10'b1011011011: data <= 18'h00073; 
        10'b1011011100: data <= 18'h3fff4; 
        10'b1011011101: data <= 18'h3ffd8; 
        10'b1011011110: data <= 18'h00045; 
        10'b1011011111: data <= 18'h00032; 
        10'b1011100000: data <= 18'h3ffcb; 
        10'b1011100001: data <= 18'h3ff0e; 
        10'b1011100010: data <= 18'h3fdb9; 
        10'b1011100011: data <= 18'h3fe03; 
        10'b1011100100: data <= 18'h3fdba; 
        10'b1011100101: data <= 18'h3fce9; 
        10'b1011100110: data <= 18'h3fca0; 
        10'b1011100111: data <= 18'h3fd60; 
        10'b1011101000: data <= 18'h3fd02; 
        10'b1011101001: data <= 18'h3fd76; 
        10'b1011101010: data <= 18'h3fdea; 
        10'b1011101011: data <= 18'h3fec2; 
        10'b1011101100: data <= 18'h3ff8c; 
        10'b1011101101: data <= 18'h000ac; 
        10'b1011101110: data <= 18'h000ab; 
        10'b1011101111: data <= 18'h00016; 
        10'b1011110000: data <= 18'h00070; 
        10'b1011110001: data <= 18'h00012; 
        10'b1011110010: data <= 18'h00113; 
        10'b1011110011: data <= 18'h00078; 
        10'b1011110100: data <= 18'h000a7; 
        10'b1011110101: data <= 18'h00018; 
        10'b1011110110: data <= 18'h00025; 
        10'b1011110111: data <= 18'h00108; 
        10'b1011111000: data <= 18'h00063; 
        10'b1011111001: data <= 18'h000dc; 
        10'b1011111010: data <= 18'h00065; 
        10'b1011111011: data <= 18'h0010d; 
        10'b1011111100: data <= 18'h3ffff; 
        10'b1011111101: data <= 18'h00074; 
        10'b1011111110: data <= 18'h0003b; 
        10'b1011111111: data <= 18'h3ffdb; 
        10'b1100000000: data <= 18'h3ffe5; 
        10'b1100000001: data <= 18'h0000a; 
        10'b1100000010: data <= 18'h3ff90; 
        10'b1100000011: data <= 18'h000d6; 
        10'b1100000100: data <= 18'h3ffc9; 
        10'b1100000101: data <= 18'h3ffc1; 
        10'b1100000110: data <= 18'h3ffeb; 
        10'b1100000111: data <= 18'h00070; 
        10'b1100001000: data <= 18'h00056; 
        10'b1100001001: data <= 18'h00056; 
        10'b1100001010: data <= 18'h0005b; 
        10'b1100001011: data <= 18'h0009c; 
        10'b1100001100: data <= 18'h00095; 
        10'b1100001101: data <= 18'h000c5; 
        10'b1100001110: data <= 18'h0008d; 
        10'b1100001111: data <= 18'h0005e; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 13) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 19'h00000; 
        10'b0000000001: data <= 19'h00048; 
        10'b0000000010: data <= 19'h001e4; 
        10'b0000000011: data <= 19'h001e3; 
        10'b0000000100: data <= 19'h00009; 
        10'b0000000101: data <= 19'h00009; 
        10'b0000000110: data <= 19'h0017b; 
        10'b0000000111: data <= 19'h00067; 
        10'b0000001000: data <= 19'h00020; 
        10'b0000001001: data <= 19'h00047; 
        10'b0000001010: data <= 19'h0000e; 
        10'b0000001011: data <= 19'h0015c; 
        10'b0000001100: data <= 19'h001ca; 
        10'b0000001101: data <= 19'h00105; 
        10'b0000001110: data <= 19'h00151; 
        10'b0000001111: data <= 19'h00025; 
        10'b0000010000: data <= 19'h0013b; 
        10'b0000010001: data <= 19'h001b0; 
        10'b0000010010: data <= 19'h0005b; 
        10'b0000010011: data <= 19'h0015d; 
        10'b0000010100: data <= 19'h0001a; 
        10'b0000010101: data <= 19'h000cf; 
        10'b0000010110: data <= 19'h001d2; 
        10'b0000010111: data <= 19'h0002e; 
        10'b0000011000: data <= 19'h001d2; 
        10'b0000011001: data <= 19'h0004a; 
        10'b0000011010: data <= 19'h001fd; 
        10'b0000011011: data <= 19'h000d2; 
        10'b0000011100: data <= 19'h00085; 
        10'b0000011101: data <= 19'h000ee; 
        10'b0000011110: data <= 19'h7fffc; 
        10'b0000011111: data <= 19'h00028; 
        10'b0000100000: data <= 19'h000e9; 
        10'b0000100001: data <= 19'h00232; 
        10'b0000100010: data <= 19'h00074; 
        10'b0000100011: data <= 19'h7ffa6; 
        10'b0000100100: data <= 19'h00138; 
        10'b0000100101: data <= 19'h0000b; 
        10'b0000100110: data <= 19'h000d1; 
        10'b0000100111: data <= 19'h7ff5c; 
        10'b0000101000: data <= 19'h00090; 
        10'b0000101001: data <= 19'h7ff1f; 
        10'b0000101010: data <= 19'h0000c; 
        10'b0000101011: data <= 19'h00135; 
        10'b0000101100: data <= 19'h0016c; 
        10'b0000101101: data <= 19'h0006b; 
        10'b0000101110: data <= 19'h00006; 
        10'b0000101111: data <= 19'h0005b; 
        10'b0000110000: data <= 19'h00187; 
        10'b0000110001: data <= 19'h7fff7; 
        10'b0000110010: data <= 19'h7fff3; 
        10'b0000110011: data <= 19'h00020; 
        10'b0000110100: data <= 19'h0015b; 
        10'b0000110101: data <= 19'h0016f; 
        10'b0000110110: data <= 19'h00057; 
        10'b0000110111: data <= 19'h0016e; 
        10'b0000111000: data <= 19'h001a3; 
        10'b0000111001: data <= 19'h00111; 
        10'b0000111010: data <= 19'h0019e; 
        10'b0000111011: data <= 19'h001a9; 
        10'b0000111100: data <= 19'h00192; 
        10'b0000111101: data <= 19'h00167; 
        10'b0000111110: data <= 19'h001dc; 
        10'b0000111111: data <= 19'h7ff68; 
        10'b0001000000: data <= 19'h7ff5c; 
        10'b0001000001: data <= 19'h00057; 
        10'b0001000010: data <= 19'h7ffc8; 
        10'b0001000011: data <= 19'h7fee5; 
        10'b0001000100: data <= 19'h7fbbb; 
        10'b0001000101: data <= 19'h7fe47; 
        10'b0001000110: data <= 19'h7fdef; 
        10'b0001000111: data <= 19'h7fd13; 
        10'b0001001000: data <= 19'h7fddf; 
        10'b0001001001: data <= 19'h7ff95; 
        10'b0001001010: data <= 19'h00088; 
        10'b0001001011: data <= 19'h00181; 
        10'b0001001100: data <= 19'h001f3; 
        10'b0001001101: data <= 19'h00120; 
        10'b0001001110: data <= 19'h001d7; 
        10'b0001001111: data <= 19'h0007f; 
        10'b0001010000: data <= 19'h000b2; 
        10'b0001010001: data <= 19'h0013e; 
        10'b0001010010: data <= 19'h00014; 
        10'b0001010011: data <= 19'h000de; 
        10'b0001010100: data <= 19'h001a7; 
        10'b0001010101: data <= 19'h0017c; 
        10'b0001010110: data <= 19'h00093; 
        10'b0001010111: data <= 19'h000ef; 
        10'b0001011000: data <= 19'h000f8; 
        10'b0001011001: data <= 19'h00003; 
        10'b0001011010: data <= 19'h0013e; 
        10'b0001011011: data <= 19'h7fee7; 
        10'b0001011100: data <= 19'h7fe65; 
        10'b0001011101: data <= 19'h7ff20; 
        10'b0001011110: data <= 19'h7fc54; 
        10'b0001011111: data <= 19'h7fba8; 
        10'b0001100000: data <= 19'h7f912; 
        10'b0001100001: data <= 19'h7f963; 
        10'b0001100010: data <= 19'h7f9b4; 
        10'b0001100011: data <= 19'h7f85c; 
        10'b0001100100: data <= 19'h7fae6; 
        10'b0001100101: data <= 19'h7fd74; 
        10'b0001100110: data <= 19'h00060; 
        10'b0001100111: data <= 19'h000d1; 
        10'b0001101000: data <= 19'h0017b; 
        10'b0001101001: data <= 19'h0022e; 
        10'b0001101010: data <= 19'h00092; 
        10'b0001101011: data <= 19'h00095; 
        10'b0001101100: data <= 19'h0021f; 
        10'b0001101101: data <= 19'h0020a; 
        10'b0001101110: data <= 19'h000a1; 
        10'b0001101111: data <= 19'h00132; 
        10'b0001110000: data <= 19'h00210; 
        10'b0001110001: data <= 19'h0015e; 
        10'b0001110010: data <= 19'h0018a; 
        10'b0001110011: data <= 19'h0017e; 
        10'b0001110100: data <= 19'h000e4; 
        10'b0001110101: data <= 19'h001b0; 
        10'b0001110110: data <= 19'h7febc; 
        10'b0001110111: data <= 19'h7ffb8; 
        10'b0001111000: data <= 19'h7fd6a; 
        10'b0001111001: data <= 19'h7fdd0; 
        10'b0001111010: data <= 19'h7f9c9; 
        10'b0001111011: data <= 19'h7fa17; 
        10'b0001111100: data <= 19'h7f7ea; 
        10'b0001111101: data <= 19'h7f949; 
        10'b0001111110: data <= 19'h7f7c2; 
        10'b0001111111: data <= 19'h7f8f1; 
        10'b0010000000: data <= 19'h7fc92; 
        10'b0010000001: data <= 19'h7fcf4; 
        10'b0010000010: data <= 19'h7fe2d; 
        10'b0010000011: data <= 19'h001c1; 
        10'b0010000100: data <= 19'h0026a; 
        10'b0010000101: data <= 19'h002c2; 
        10'b0010000110: data <= 19'h002a1; 
        10'b0010000111: data <= 19'h0037c; 
        10'b0010001000: data <= 19'h000f7; 
        10'b0010001001: data <= 19'h001f5; 
        10'b0010001010: data <= 19'h00080; 
        10'b0010001011: data <= 19'h00052; 
        10'b0010001100: data <= 19'h00219; 
        10'b0010001101: data <= 19'h00096; 
        10'b0010001110: data <= 19'h0017b; 
        10'b0010001111: data <= 19'h0007c; 
        10'b0010010000: data <= 19'h0015b; 
        10'b0010010001: data <= 19'h00046; 
        10'b0010010010: data <= 19'h000f6; 
        10'b0010010011: data <= 19'h7fed6; 
        10'b0010010100: data <= 19'h00050; 
        10'b0010010101: data <= 19'h7fea7; 
        10'b0010010110: data <= 19'h7fb74; 
        10'b0010010111: data <= 19'h7fcfd; 
        10'b0010011000: data <= 19'h7fad6; 
        10'b0010011001: data <= 19'h7f997; 
        10'b0010011010: data <= 19'h7fb84; 
        10'b0010011011: data <= 19'h7fc4d; 
        10'b0010011100: data <= 19'h7ff61; 
        10'b0010011101: data <= 19'h00091; 
        10'b0010011110: data <= 19'h7ff1d; 
        10'b0010011111: data <= 19'h0017e; 
        10'b0010100000: data <= 19'h001d5; 
        10'b0010100001: data <= 19'h00279; 
        10'b0010100010: data <= 19'h005c4; 
        10'b0010100011: data <= 19'h00681; 
        10'b0010100100: data <= 19'h0038a; 
        10'b0010100101: data <= 19'h7ffa7; 
        10'b0010100110: data <= 19'h00095; 
        10'b0010100111: data <= 19'h0005a; 
        10'b0010101000: data <= 19'h001f2; 
        10'b0010101001: data <= 19'h00227; 
        10'b0010101010: data <= 19'h000a4; 
        10'b0010101011: data <= 19'h001b1; 
        10'b0010101100: data <= 19'h001d7; 
        10'b0010101101: data <= 19'h00183; 
        10'b0010101110: data <= 19'h00180; 
        10'b0010101111: data <= 19'h7ffe2; 
        10'b0010110000: data <= 19'h7ffa9; 
        10'b0010110001: data <= 19'h7fe37; 
        10'b0010110010: data <= 19'h7fc65; 
        10'b0010110011: data <= 19'h7f9a8; 
        10'b0010110100: data <= 19'h7f664; 
        10'b0010110101: data <= 19'h7f4a3; 
        10'b0010110110: data <= 19'h7f422; 
        10'b0010110111: data <= 19'h7f5b3; 
        10'b0010111000: data <= 19'h7f572; 
        10'b0010111001: data <= 19'h7f9d0; 
        10'b0010111010: data <= 19'h7f99b; 
        10'b0010111011: data <= 19'h7fd20; 
        10'b0010111100: data <= 19'h7fe1c; 
        10'b0010111101: data <= 19'h7ffdb; 
        10'b0010111110: data <= 19'h00840; 
        10'b0010111111: data <= 19'h008ab; 
        10'b0011000000: data <= 19'h00356; 
        10'b0011000001: data <= 19'h0029d; 
        10'b0011000010: data <= 19'h001de; 
        10'b0011000011: data <= 19'h00014; 
        10'b0011000100: data <= 19'h000eb; 
        10'b0011000101: data <= 19'h0007b; 
        10'b0011000110: data <= 19'h000a9; 
        10'b0011000111: data <= 19'h0012c; 
        10'b0011001000: data <= 19'h000ac; 
        10'b0011001001: data <= 19'h00191; 
        10'b0011001010: data <= 19'h7ff08; 
        10'b0011001011: data <= 19'h7ffd3; 
        10'b0011001100: data <= 19'h7feed; 
        10'b0011001101: data <= 19'h7fd90; 
        10'b0011001110: data <= 19'h7f9d8; 
        10'b0011001111: data <= 19'h7f666; 
        10'b0011010000: data <= 19'h7f388; 
        10'b0011010001: data <= 19'h7f730; 
        10'b0011010010: data <= 19'h7f4fb; 
        10'b0011010011: data <= 19'h7f4e6; 
        10'b0011010100: data <= 19'h7f495; 
        10'b0011010101: data <= 19'h7f8b8; 
        10'b0011010110: data <= 19'h7f88b; 
        10'b0011010111: data <= 19'h7facf; 
        10'b0011011000: data <= 19'h7fa00; 
        10'b0011011001: data <= 19'h7fd43; 
        10'b0011011010: data <= 19'h00519; 
        10'b0011011011: data <= 19'h006e6; 
        10'b0011011100: data <= 19'h003ae; 
        10'b0011011101: data <= 19'h00213; 
        10'b0011011110: data <= 19'h001f1; 
        10'b0011011111: data <= 19'h00127; 
        10'b0011100000: data <= 19'h001df; 
        10'b0011100001: data <= 19'h00192; 
        10'b0011100010: data <= 19'h00212; 
        10'b0011100011: data <= 19'h00066; 
        10'b0011100100: data <= 19'h0009f; 
        10'b0011100101: data <= 19'h000da; 
        10'b0011100110: data <= 19'h00093; 
        10'b0011100111: data <= 19'h7ff81; 
        10'b0011101000: data <= 19'h7fb5c; 
        10'b0011101001: data <= 19'h7fda4; 
        10'b0011101010: data <= 19'h7fcea; 
        10'b0011101011: data <= 19'h7f9cc; 
        10'b0011101100: data <= 19'h7f6ea; 
        10'b0011101101: data <= 19'h7fa31; 
        10'b0011101110: data <= 19'h7f2d6; 
        10'b0011101111: data <= 19'h7f27a; 
        10'b0011110000: data <= 19'h7f57d; 
        10'b0011110001: data <= 19'h7f96b; 
        10'b0011110010: data <= 19'h7fa17; 
        10'b0011110011: data <= 19'h7fe24; 
        10'b0011110100: data <= 19'h7fc65; 
        10'b0011110101: data <= 19'h7fc75; 
        10'b0011110110: data <= 19'h00259; 
        10'b0011110111: data <= 19'h0039d; 
        10'b0011111000: data <= 19'h002c2; 
        10'b0011111001: data <= 19'h0008c; 
        10'b0011111010: data <= 19'h000be; 
        10'b0011111011: data <= 19'h0015a; 
        10'b0011111100: data <= 19'h0023a; 
        10'b0011111101: data <= 19'h001df; 
        10'b0011111110: data <= 19'h001c0; 
        10'b0011111111: data <= 19'h0005e; 
        10'b0100000000: data <= 19'h7fed7; 
        10'b0100000001: data <= 19'h00009; 
        10'b0100000010: data <= 19'h7fd23; 
        10'b0100000011: data <= 19'h7fdf2; 
        10'b0100000100: data <= 19'h7feab; 
        10'b0100000101: data <= 19'h7ff90; 
        10'b0100000110: data <= 19'h7fe69; 
        10'b0100000111: data <= 19'h7fe17; 
        10'b0100001000: data <= 19'h7fe08; 
        10'b0100001001: data <= 19'h7fac3; 
        10'b0100001010: data <= 19'h7ed06; 
        10'b0100001011: data <= 19'h7f1ce; 
        10'b0100001100: data <= 19'h7fc8e; 
        10'b0100001101: data <= 19'h7fd74; 
        10'b0100001110: data <= 19'h7ff37; 
        10'b0100001111: data <= 19'h0006c; 
        10'b0100010000: data <= 19'h7fe02; 
        10'b0100010001: data <= 19'h7fe0d; 
        10'b0100010010: data <= 19'h000fc; 
        10'b0100010011: data <= 19'h00039; 
        10'b0100010100: data <= 19'h7fdbe; 
        10'b0100010101: data <= 19'h7fda6; 
        10'b0100010110: data <= 19'h7fefb; 
        10'b0100010111: data <= 19'h00181; 
        10'b0100011000: data <= 19'h00130; 
        10'b0100011001: data <= 19'h000d7; 
        10'b0100011010: data <= 19'h000d9; 
        10'b0100011011: data <= 19'h0003c; 
        10'b0100011100: data <= 19'h000e2; 
        10'b0100011101: data <= 19'h7fd72; 
        10'b0100011110: data <= 19'h7fbc6; 
        10'b0100011111: data <= 19'h7fdf3; 
        10'b0100100000: data <= 19'h0009c; 
        10'b0100100001: data <= 19'h00568; 
        10'b0100100010: data <= 19'h00346; 
        10'b0100100011: data <= 19'h00272; 
        10'b0100100100: data <= 19'h002ee; 
        10'b0100100101: data <= 19'h7f8be; 
        10'b0100100110: data <= 19'h7ebf6; 
        10'b0100100111: data <= 19'h7f9e4; 
        10'b0100101000: data <= 19'h000b3; 
        10'b0100101001: data <= 19'h7ff1a; 
        10'b0100101010: data <= 19'h7ff50; 
        10'b0100101011: data <= 19'h000b5; 
        10'b0100101100: data <= 19'h7fc00; 
        10'b0100101101: data <= 19'h7fd5c; 
        10'b0100101110: data <= 19'h7ff80; 
        10'b0100101111: data <= 19'h7fba5; 
        10'b0100110000: data <= 19'h7fd88; 
        10'b0100110001: data <= 19'h7fe6f; 
        10'b0100110010: data <= 19'h0013f; 
        10'b0100110011: data <= 19'h00210; 
        10'b0100110100: data <= 19'h00163; 
        10'b0100110101: data <= 19'h00172; 
        10'b0100110110: data <= 19'h00139; 
        10'b0100110111: data <= 19'h7ff3c; 
        10'b0100111000: data <= 19'h7ffb8; 
        10'b0100111001: data <= 19'h7fe92; 
        10'b0100111010: data <= 19'h7fe7d; 
        10'b0100111011: data <= 19'h00148; 
        10'b0100111100: data <= 19'h00418; 
        10'b0100111101: data <= 19'h006e5; 
        10'b0100111110: data <= 19'h00981; 
        10'b0100111111: data <= 19'h0060b; 
        10'b0101000000: data <= 19'h006d3; 
        10'b0101000001: data <= 19'h7f4e2; 
        10'b0101000010: data <= 19'h7f0e9; 
        10'b0101000011: data <= 19'h001f5; 
        10'b0101000100: data <= 19'h007ce; 
        10'b0101000101: data <= 19'h00151; 
        10'b0101000110: data <= 19'h7ff8c; 
        10'b0101000111: data <= 19'h7fec0; 
        10'b0101001000: data <= 19'h7fbbb; 
        10'b0101001001: data <= 19'h7fc5a; 
        10'b0101001010: data <= 19'h7fe24; 
        10'b0101001011: data <= 19'h7fca0; 
        10'b0101001100: data <= 19'h7fc40; 
        10'b0101001101: data <= 19'h7ffca; 
        10'b0101001110: data <= 19'h7ffdf; 
        10'b0101001111: data <= 19'h00084; 
        10'b0101010000: data <= 19'h0018d; 
        10'b0101010001: data <= 19'h0015c; 
        10'b0101010010: data <= 19'h000a5; 
        10'b0101010011: data <= 19'h000ee; 
        10'b0101010100: data <= 19'h7ffe8; 
        10'b0101010101: data <= 19'h7fe9b; 
        10'b0101010110: data <= 19'h00404; 
        10'b0101010111: data <= 19'h0069e; 
        10'b0101011000: data <= 19'h00a3f; 
        10'b0101011001: data <= 19'h008fb; 
        10'b0101011010: data <= 19'h00eef; 
        10'b0101011011: data <= 19'h010ec; 
        10'b0101011100: data <= 19'h00ffe; 
        10'b0101011101: data <= 19'h7ffbc; 
        10'b0101011110: data <= 19'h7f80b; 
        10'b0101011111: data <= 19'h00642; 
        10'b0101100000: data <= 19'h00a2a; 
        10'b0101100001: data <= 19'h00128; 
        10'b0101100010: data <= 19'h0006e; 
        10'b0101100011: data <= 19'h00163; 
        10'b0101100100: data <= 19'h7ffc1; 
        10'b0101100101: data <= 19'h0004d; 
        10'b0101100110: data <= 19'h7ff8c; 
        10'b0101100111: data <= 19'h7fdc2; 
        10'b0101101000: data <= 19'h7fdff; 
        10'b0101101001: data <= 19'h7ff70; 
        10'b0101101010: data <= 19'h00235; 
        10'b0101101011: data <= 19'h00147; 
        10'b0101101100: data <= 19'h0003e; 
        10'b0101101101: data <= 19'h00174; 
        10'b0101101110: data <= 19'h00034; 
        10'b0101101111: data <= 19'h0009c; 
        10'b0101110000: data <= 19'h001b7; 
        10'b0101110001: data <= 19'h004d7; 
        10'b0101110010: data <= 19'h009da; 
        10'b0101110011: data <= 19'h00b6e; 
        10'b0101110100: data <= 19'h00d24; 
        10'b0101110101: data <= 19'h00afb; 
        10'b0101110110: data <= 19'h00cd0; 
        10'b0101110111: data <= 19'h014e2; 
        10'b0101111000: data <= 19'h00fd4; 
        10'b0101111001: data <= 19'h0003d; 
        10'b0101111010: data <= 19'h7fdc1; 
        10'b0101111011: data <= 19'h00756; 
        10'b0101111100: data <= 19'h00789; 
        10'b0101111101: data <= 19'h0085e; 
        10'b0101111110: data <= 19'h005c5; 
        10'b0101111111: data <= 19'h00299; 
        10'b0110000000: data <= 19'h005c7; 
        10'b0110000001: data <= 19'h00441; 
        10'b0110000010: data <= 19'h00207; 
        10'b0110000011: data <= 19'h7fed2; 
        10'b0110000100: data <= 19'h7fef6; 
        10'b0110000101: data <= 19'h0001e; 
        10'b0110000110: data <= 19'h001c6; 
        10'b0110000111: data <= 19'h00145; 
        10'b0110001000: data <= 19'h0003a; 
        10'b0110001001: data <= 19'h001d0; 
        10'b0110001010: data <= 19'h00025; 
        10'b0110001011: data <= 19'h00222; 
        10'b0110001100: data <= 19'h00449; 
        10'b0110001101: data <= 19'h008a1; 
        10'b0110001110: data <= 19'h00bfe; 
        10'b0110001111: data <= 19'h00d20; 
        10'b0110010000: data <= 19'h009cf; 
        10'b0110010001: data <= 19'h00960; 
        10'b0110010010: data <= 19'h00b4b; 
        10'b0110010011: data <= 19'h00db0; 
        10'b0110010100: data <= 19'h009f7; 
        10'b0110010101: data <= 19'h000d3; 
        10'b0110010110: data <= 19'h7fe8d; 
        10'b0110010111: data <= 19'h002a6; 
        10'b0110011000: data <= 19'h00864; 
        10'b0110011001: data <= 19'h00dca; 
        10'b0110011010: data <= 19'h0095d; 
        10'b0110011011: data <= 19'h0089b; 
        10'b0110011100: data <= 19'h004ce; 
        10'b0110011101: data <= 19'h0033b; 
        10'b0110011110: data <= 19'h0010d; 
        10'b0110011111: data <= 19'h00098; 
        10'b0110100000: data <= 19'h7ffa9; 
        10'b0110100001: data <= 19'h00093; 
        10'b0110100010: data <= 19'h00114; 
        10'b0110100011: data <= 19'h00082; 
        10'b0110100100: data <= 19'h0017f; 
        10'b0110100101: data <= 19'h00226; 
        10'b0110100110: data <= 19'h00161; 
        10'b0110100111: data <= 19'h001c6; 
        10'b0110101000: data <= 19'h003e0; 
        10'b0110101001: data <= 19'h00465; 
        10'b0110101010: data <= 19'h006d4; 
        10'b0110101011: data <= 19'h0064a; 
        10'b0110101100: data <= 19'h00a1f; 
        10'b0110101101: data <= 19'h008b2; 
        10'b0110101110: data <= 19'h0060d; 
        10'b0110101111: data <= 19'h00465; 
        10'b0110110000: data <= 19'h00531; 
        10'b0110110001: data <= 19'h00106; 
        10'b0110110010: data <= 19'h0042a; 
        10'b0110110011: data <= 19'h005d3; 
        10'b0110110100: data <= 19'h00c17; 
        10'b0110110101: data <= 19'h00abe; 
        10'b0110110110: data <= 19'h007ae; 
        10'b0110110111: data <= 19'h0048d; 
        10'b0110111000: data <= 19'h7fec7; 
        10'b0110111001: data <= 19'h001b0; 
        10'b0110111010: data <= 19'h0030d; 
        10'b0110111011: data <= 19'h00052; 
        10'b0110111100: data <= 19'h7fe29; 
        10'b0110111101: data <= 19'h000f8; 
        10'b0110111110: data <= 19'h0003f; 
        10'b0110111111: data <= 19'h0009c; 
        10'b0111000000: data <= 19'h000aa; 
        10'b0111000001: data <= 19'h00003; 
        10'b0111000010: data <= 19'h00014; 
        10'b0111000011: data <= 19'h7ffbc; 
        10'b0111000100: data <= 19'h0010e; 
        10'b0111000101: data <= 19'h00298; 
        10'b0111000110: data <= 19'h0043a; 
        10'b0111000111: data <= 19'h00761; 
        10'b0111001000: data <= 19'h00abe; 
        10'b0111001001: data <= 19'h007a7; 
        10'b0111001010: data <= 19'h0020d; 
        10'b0111001011: data <= 19'h7ffb9; 
        10'b0111001100: data <= 19'h0021b; 
        10'b0111001101: data <= 19'h002a0; 
        10'b0111001110: data <= 19'h009dc; 
        10'b0111001111: data <= 19'h00da2; 
        10'b0111010000: data <= 19'h00e0a; 
        10'b0111010001: data <= 19'h00baa; 
        10'b0111010010: data <= 19'h007e5; 
        10'b0111010011: data <= 19'h000fd; 
        10'b0111010100: data <= 19'h00350; 
        10'b0111010101: data <= 19'h004b4; 
        10'b0111010110: data <= 19'h00119; 
        10'b0111010111: data <= 19'h7ff39; 
        10'b0111011000: data <= 19'h7ffc9; 
        10'b0111011001: data <= 19'h00075; 
        10'b0111011010: data <= 19'h000d9; 
        10'b0111011011: data <= 19'h000e4; 
        10'b0111011100: data <= 19'h000ca; 
        10'b0111011101: data <= 19'h000ce; 
        10'b0111011110: data <= 19'h0019b; 
        10'b0111011111: data <= 19'h7fff9; 
        10'b0111100000: data <= 19'h7fedf; 
        10'b0111100001: data <= 19'h7fdae; 
        10'b0111100010: data <= 19'h0015f; 
        10'b0111100011: data <= 19'h005da; 
        10'b0111100100: data <= 19'h00b49; 
        10'b0111100101: data <= 19'h009c9; 
        10'b0111100110: data <= 19'h0038b; 
        10'b0111100111: data <= 19'h002ca; 
        10'b0111101000: data <= 19'h0040a; 
        10'b0111101001: data <= 19'h009ae; 
        10'b0111101010: data <= 19'h00ffe; 
        10'b0111101011: data <= 19'h00ca8; 
        10'b0111101100: data <= 19'h00a97; 
        10'b0111101101: data <= 19'h00345; 
        10'b0111101110: data <= 19'h00081; 
        10'b0111101111: data <= 19'h7fc75; 
        10'b0111110000: data <= 19'h00110; 
        10'b0111110001: data <= 19'h00063; 
        10'b0111110010: data <= 19'h7fdd6; 
        10'b0111110011: data <= 19'h7ff11; 
        10'b0111110100: data <= 19'h7fe97; 
        10'b0111110101: data <= 19'h7ff31; 
        10'b0111110110: data <= 19'h0016d; 
        10'b0111110111: data <= 19'h001be; 
        10'b0111111000: data <= 19'h000df; 
        10'b0111111001: data <= 19'h00156; 
        10'b0111111010: data <= 19'h0012b; 
        10'b0111111011: data <= 19'h0002d; 
        10'b0111111100: data <= 19'h7fea3; 
        10'b0111111101: data <= 19'h7fd22; 
        10'b0111111110: data <= 19'h7fcac; 
        10'b0111111111: data <= 19'h7ffef; 
        10'b1000000000: data <= 19'h002e3; 
        10'b1000000001: data <= 19'h000a9; 
        10'b1000000010: data <= 19'h7fda6; 
        10'b1000000011: data <= 19'h7fe9c; 
        10'b1000000100: data <= 19'h003b1; 
        10'b1000000101: data <= 19'h00429; 
        10'b1000000110: data <= 19'h00707; 
        10'b1000000111: data <= 19'h00604; 
        10'b1000001000: data <= 19'h00324; 
        10'b1000001001: data <= 19'h7fb23; 
        10'b1000001010: data <= 19'h7fb64; 
        10'b1000001011: data <= 19'h7f93e; 
        10'b1000001100: data <= 19'h7fbfe; 
        10'b1000001101: data <= 19'h7fbd8; 
        10'b1000001110: data <= 19'h7fa76; 
        10'b1000001111: data <= 19'h7fbb5; 
        10'b1000010000: data <= 19'h7fee2; 
        10'b1000010001: data <= 19'h7ff68; 
        10'b1000010010: data <= 19'h00084; 
        10'b1000010011: data <= 19'h00012; 
        10'b1000010100: data <= 19'h000d8; 
        10'b1000010101: data <= 19'h00190; 
        10'b1000010110: data <= 19'h00098; 
        10'b1000010111: data <= 19'h0005b; 
        10'b1000011000: data <= 19'h7fce8; 
        10'b1000011001: data <= 19'h7fc28; 
        10'b1000011010: data <= 19'h7faec; 
        10'b1000011011: data <= 19'h7f85f; 
        10'b1000011100: data <= 19'h7f765; 
        10'b1000011101: data <= 19'h7f6d4; 
        10'b1000011110: data <= 19'h7f52e; 
        10'b1000011111: data <= 19'h7f5a7; 
        10'b1000100000: data <= 19'h7f6d6; 
        10'b1000100001: data <= 19'h7faa1; 
        10'b1000100010: data <= 19'h7fe68; 
        10'b1000100011: data <= 19'h00165; 
        10'b1000100100: data <= 19'h7fbd5; 
        10'b1000100101: data <= 19'h7fc6a; 
        10'b1000100110: data <= 19'h7fb95; 
        10'b1000100111: data <= 19'h7f9e7; 
        10'b1000101000: data <= 19'h7f930; 
        10'b1000101001: data <= 19'h7f9b9; 
        10'b1000101010: data <= 19'h7f99f; 
        10'b1000101011: data <= 19'h7fbb0; 
        10'b1000101100: data <= 19'h7fedd; 
        10'b1000101101: data <= 19'h000db; 
        10'b1000101110: data <= 19'h00183; 
        10'b1000101111: data <= 19'h00161; 
        10'b1000110000: data <= 19'h00240; 
        10'b1000110001: data <= 19'h00215; 
        10'b1000110010: data <= 19'h0009a; 
        10'b1000110011: data <= 19'h0005c; 
        10'b1000110100: data <= 19'h7fd7d; 
        10'b1000110101: data <= 19'h7fbb5; 
        10'b1000110110: data <= 19'h7f9c3; 
        10'b1000110111: data <= 19'h7f5d9; 
        10'b1000111000: data <= 19'h7f3ee; 
        10'b1000111001: data <= 19'h7f336; 
        10'b1000111010: data <= 19'h7f2fa; 
        10'b1000111011: data <= 19'h7f677; 
        10'b1000111100: data <= 19'h7f84a; 
        10'b1000111101: data <= 19'h7f761; 
        10'b1000111110: data <= 19'h7fa95; 
        10'b1000111111: data <= 19'h7fd2d; 
        10'b1001000000: data <= 19'h7ff06; 
        10'b1001000001: data <= 19'h7ff75; 
        10'b1001000010: data <= 19'h7fdc3; 
        10'b1001000011: data <= 19'h7fb26; 
        10'b1001000100: data <= 19'h7fcbd; 
        10'b1001000101: data <= 19'h7fc4f; 
        10'b1001000110: data <= 19'h7fb8b; 
        10'b1001000111: data <= 19'h7fdb7; 
        10'b1001001000: data <= 19'h7fdce; 
        10'b1001001001: data <= 19'h00029; 
        10'b1001001010: data <= 19'h00087; 
        10'b1001001011: data <= 19'h00181; 
        10'b1001001100: data <= 19'h0006a; 
        10'b1001001101: data <= 19'h000a8; 
        10'b1001001110: data <= 19'h0002c; 
        10'b1001001111: data <= 19'h0004d; 
        10'b1001010000: data <= 19'h7fffa; 
        10'b1001010001: data <= 19'h7fd8e; 
        10'b1001010010: data <= 19'h7f9da; 
        10'b1001010011: data <= 19'h7f763; 
        10'b1001010100: data <= 19'h7f83f; 
        10'b1001010101: data <= 19'h7f72f; 
        10'b1001010110: data <= 19'h7f853; 
        10'b1001010111: data <= 19'h7fa4d; 
        10'b1001011000: data <= 19'h7fb43; 
        10'b1001011001: data <= 19'h7fb9c; 
        10'b1001011010: data <= 19'h7faf9; 
        10'b1001011011: data <= 19'h7fdac; 
        10'b1001011100: data <= 19'h7fce6; 
        10'b1001011101: data <= 19'h0008f; 
        10'b1001011110: data <= 19'h7ff13; 
        10'b1001011111: data <= 19'h0002b; 
        10'b1001100000: data <= 19'h7ff99; 
        10'b1001100001: data <= 19'h7fcfb; 
        10'b1001100010: data <= 19'h7fd71; 
        10'b1001100011: data <= 19'h7ff87; 
        10'b1001100100: data <= 19'h7ffeb; 
        10'b1001100101: data <= 19'h000ee; 
        10'b1001100110: data <= 19'h00140; 
        10'b1001100111: data <= 19'h00134; 
        10'b1001101000: data <= 19'h00115; 
        10'b1001101001: data <= 19'h00142; 
        10'b1001101010: data <= 19'h00080; 
        10'b1001101011: data <= 19'h00161; 
        10'b1001101100: data <= 19'h7ffad; 
        10'b1001101101: data <= 19'h7feb2; 
        10'b1001101110: data <= 19'h7fd77; 
        10'b1001101111: data <= 19'h7fbd0; 
        10'b1001110000: data <= 19'h7fa57; 
        10'b1001110001: data <= 19'h7fc90; 
        10'b1001110010: data <= 19'h7fc75; 
        10'b1001110011: data <= 19'h7fd8b; 
        10'b1001110100: data <= 19'h7fd69; 
        10'b1001110101: data <= 19'h7fdc7; 
        10'b1001110110: data <= 19'h7fd39; 
        10'b1001110111: data <= 19'h7fe4b; 
        10'b1001111000: data <= 19'h7fe5d; 
        10'b1001111001: data <= 19'h00097; 
        10'b1001111010: data <= 19'h00283; 
        10'b1001111011: data <= 19'h00418; 
        10'b1001111100: data <= 19'h00325; 
        10'b1001111101: data <= 19'h00210; 
        10'b1001111110: data <= 19'h7fea3; 
        10'b1001111111: data <= 19'h7fea9; 
        10'b1010000000: data <= 19'h7fff3; 
        10'b1010000001: data <= 19'h000e6; 
        10'b1010000010: data <= 19'h00025; 
        10'b1010000011: data <= 19'h000b1; 
        10'b1010000100: data <= 19'h000b4; 
        10'b1010000101: data <= 19'h0000c; 
        10'b1010000110: data <= 19'h0009f; 
        10'b1010000111: data <= 19'h0013a; 
        10'b1010001000: data <= 19'h000b2; 
        10'b1010001001: data <= 19'h000da; 
        10'b1010001010: data <= 19'h7fea6; 
        10'b1010001011: data <= 19'h7fe7f; 
        10'b1010001100: data <= 19'h7fdf8; 
        10'b1010001101: data <= 19'h000f3; 
        10'b1010001110: data <= 19'h7fdd0; 
        10'b1010001111: data <= 19'h0005a; 
        10'b1010010000: data <= 19'h7fdbd; 
        10'b1010010001: data <= 19'h7fe39; 
        10'b1010010010: data <= 19'h7fe43; 
        10'b1010010011: data <= 19'h7ffdf; 
        10'b1010010100: data <= 19'h00094; 
        10'b1010010101: data <= 19'h00187; 
        10'b1010010110: data <= 19'h004b6; 
        10'b1010010111: data <= 19'h00499; 
        10'b1010011000: data <= 19'h003eb; 
        10'b1010011001: data <= 19'h001bf; 
        10'b1010011010: data <= 19'h7ff5a; 
        10'b1010011011: data <= 19'h00088; 
        10'b1010011100: data <= 19'h0010a; 
        10'b1010011101: data <= 19'h0016c; 
        10'b1010011110: data <= 19'h00077; 
        10'b1010011111: data <= 19'h001c5; 
        10'b1010100000: data <= 19'h00157; 
        10'b1010100001: data <= 19'h001e9; 
        10'b1010100010: data <= 19'h000e8; 
        10'b1010100011: data <= 19'h00184; 
        10'b1010100100: data <= 19'h0005b; 
        10'b1010100101: data <= 19'h00129; 
        10'b1010100110: data <= 19'h00071; 
        10'b1010100111: data <= 19'h7fdd9; 
        10'b1010101000: data <= 19'h7fdcd; 
        10'b1010101001: data <= 19'h7ff4d; 
        10'b1010101010: data <= 19'h7fdab; 
        10'b1010101011: data <= 19'h7ff9f; 
        10'b1010101100: data <= 19'h7fe53; 
        10'b1010101101: data <= 19'h7fe75; 
        10'b1010101110: data <= 19'h7fd28; 
        10'b1010101111: data <= 19'h7fccf; 
        10'b1010110000: data <= 19'h7fea0; 
        10'b1010110001: data <= 19'h7ff49; 
        10'b1010110010: data <= 19'h00040; 
        10'b1010110011: data <= 19'h0027a; 
        10'b1010110100: data <= 19'h001cf; 
        10'b1010110101: data <= 19'h7ff42; 
        10'b1010110110: data <= 19'h7ffc9; 
        10'b1010110111: data <= 19'h000f5; 
        10'b1010111000: data <= 19'h00193; 
        10'b1010111001: data <= 19'h00040; 
        10'b1010111010: data <= 19'h00069; 
        10'b1010111011: data <= 19'h0015d; 
        10'b1010111100: data <= 19'h00200; 
        10'b1010111101: data <= 19'h001f1; 
        10'b1010111110: data <= 19'h001c6; 
        10'b1010111111: data <= 19'h00066; 
        10'b1011000000: data <= 19'h001c9; 
        10'b1011000001: data <= 19'h00016; 
        10'b1011000010: data <= 19'h7feb9; 
        10'b1011000011: data <= 19'h7fdec; 
        10'b1011000100: data <= 19'h7fce0; 
        10'b1011000101: data <= 19'h7fcb7; 
        10'b1011000110: data <= 19'h7fa9b; 
        10'b1011000111: data <= 19'h7f9ea; 
        10'b1011001000: data <= 19'h7fa41; 
        10'b1011001001: data <= 19'h7fa48; 
        10'b1011001010: data <= 19'h7fb24; 
        10'b1011001011: data <= 19'h7fadc; 
        10'b1011001100: data <= 19'h7f959; 
        10'b1011001101: data <= 19'h7f86a; 
        10'b1011001110: data <= 19'h7f930; 
        10'b1011001111: data <= 19'h7fc44; 
        10'b1011010000: data <= 19'h7fc96; 
        10'b1011010001: data <= 19'h7fec4; 
        10'b1011010010: data <= 19'h00013; 
        10'b1011010011: data <= 19'h0014e; 
        10'b1011010100: data <= 19'h00019; 
        10'b1011010101: data <= 19'h001d0; 
        10'b1011010110: data <= 19'h000ba; 
        10'b1011010111: data <= 19'h000a9; 
        10'b1011011000: data <= 19'h000f0; 
        10'b1011011001: data <= 19'h0015a; 
        10'b1011011010: data <= 19'h0004e; 
        10'b1011011011: data <= 19'h000e6; 
        10'b1011011100: data <= 19'h7ffe9; 
        10'b1011011101: data <= 19'h7ffb1; 
        10'b1011011110: data <= 19'h0008b; 
        10'b1011011111: data <= 19'h00064; 
        10'b1011100000: data <= 19'h7ff97; 
        10'b1011100001: data <= 19'h7fe1c; 
        10'b1011100010: data <= 19'h7fb72; 
        10'b1011100011: data <= 19'h7fc07; 
        10'b1011100100: data <= 19'h7fb74; 
        10'b1011100101: data <= 19'h7f9d3; 
        10'b1011100110: data <= 19'h7f941; 
        10'b1011100111: data <= 19'h7fac0; 
        10'b1011101000: data <= 19'h7fa05; 
        10'b1011101001: data <= 19'h7faec; 
        10'b1011101010: data <= 19'h7fbd5; 
        10'b1011101011: data <= 19'h7fd84; 
        10'b1011101100: data <= 19'h7ff17; 
        10'b1011101101: data <= 19'h00159; 
        10'b1011101110: data <= 19'h00155; 
        10'b1011101111: data <= 19'h0002b; 
        10'b1011110000: data <= 19'h000e0; 
        10'b1011110001: data <= 19'h00025; 
        10'b1011110010: data <= 19'h00225; 
        10'b1011110011: data <= 19'h000f1; 
        10'b1011110100: data <= 19'h0014d; 
        10'b1011110101: data <= 19'h00031; 
        10'b1011110110: data <= 19'h0004a; 
        10'b1011110111: data <= 19'h00210; 
        10'b1011111000: data <= 19'h000c6; 
        10'b1011111001: data <= 19'h001b8; 
        10'b1011111010: data <= 19'h000cb; 
        10'b1011111011: data <= 19'h0021b; 
        10'b1011111100: data <= 19'h7ffff; 
        10'b1011111101: data <= 19'h000e8; 
        10'b1011111110: data <= 19'h00077; 
        10'b1011111111: data <= 19'h7ffb5; 
        10'b1100000000: data <= 19'h7ffc9; 
        10'b1100000001: data <= 19'h00014; 
        10'b1100000010: data <= 19'h7ff20; 
        10'b1100000011: data <= 19'h001ab; 
        10'b1100000100: data <= 19'h7ff92; 
        10'b1100000101: data <= 19'h7ff83; 
        10'b1100000110: data <= 19'h7ffd6; 
        10'b1100000111: data <= 19'h000e1; 
        10'b1100001000: data <= 19'h000ad; 
        10'b1100001001: data <= 19'h000ac; 
        10'b1100001010: data <= 19'h000b7; 
        10'b1100001011: data <= 19'h00138; 
        10'b1100001100: data <= 19'h0012a; 
        10'b1100001101: data <= 19'h0018a; 
        10'b1100001110: data <= 19'h0011b; 
        10'b1100001111: data <= 19'h000bb; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 14) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 20'hfffff; 
        10'b0000000001: data <= 20'h00090; 
        10'b0000000010: data <= 20'h003c8; 
        10'b0000000011: data <= 20'h003c6; 
        10'b0000000100: data <= 20'h00012; 
        10'b0000000101: data <= 20'h00012; 
        10'b0000000110: data <= 20'h002f6; 
        10'b0000000111: data <= 20'h000cf; 
        10'b0000001000: data <= 20'h00040; 
        10'b0000001001: data <= 20'h0008f; 
        10'b0000001010: data <= 20'h0001c; 
        10'b0000001011: data <= 20'h002b8; 
        10'b0000001100: data <= 20'h00394; 
        10'b0000001101: data <= 20'h00209; 
        10'b0000001110: data <= 20'h002a1; 
        10'b0000001111: data <= 20'h0004b; 
        10'b0000010000: data <= 20'h00276; 
        10'b0000010001: data <= 20'h00360; 
        10'b0000010010: data <= 20'h000b6; 
        10'b0000010011: data <= 20'h002b9; 
        10'b0000010100: data <= 20'h00034; 
        10'b0000010101: data <= 20'h0019e; 
        10'b0000010110: data <= 20'h003a4; 
        10'b0000010111: data <= 20'h0005d; 
        10'b0000011000: data <= 20'h003a4; 
        10'b0000011001: data <= 20'h00094; 
        10'b0000011010: data <= 20'h003fb; 
        10'b0000011011: data <= 20'h001a4; 
        10'b0000011100: data <= 20'h0010b; 
        10'b0000011101: data <= 20'h001dd; 
        10'b0000011110: data <= 20'hffff8; 
        10'b0000011111: data <= 20'h00050; 
        10'b0000100000: data <= 20'h001d2; 
        10'b0000100001: data <= 20'h00464; 
        10'b0000100010: data <= 20'h000e8; 
        10'b0000100011: data <= 20'hfff4c; 
        10'b0000100100: data <= 20'h00270; 
        10'b0000100101: data <= 20'h00016; 
        10'b0000100110: data <= 20'h001a3; 
        10'b0000100111: data <= 20'hffeb9; 
        10'b0000101000: data <= 20'h00120; 
        10'b0000101001: data <= 20'hffe3d; 
        10'b0000101010: data <= 20'h00018; 
        10'b0000101011: data <= 20'h0026a; 
        10'b0000101100: data <= 20'h002d8; 
        10'b0000101101: data <= 20'h000d6; 
        10'b0000101110: data <= 20'h0000b; 
        10'b0000101111: data <= 20'h000b7; 
        10'b0000110000: data <= 20'h0030f; 
        10'b0000110001: data <= 20'hfffed; 
        10'b0000110010: data <= 20'hfffe6; 
        10'b0000110011: data <= 20'h00040; 
        10'b0000110100: data <= 20'h002b5; 
        10'b0000110101: data <= 20'h002de; 
        10'b0000110110: data <= 20'h000ae; 
        10'b0000110111: data <= 20'h002dc; 
        10'b0000111000: data <= 20'h00347; 
        10'b0000111001: data <= 20'h00221; 
        10'b0000111010: data <= 20'h0033c; 
        10'b0000111011: data <= 20'h00351; 
        10'b0000111100: data <= 20'h00324; 
        10'b0000111101: data <= 20'h002cd; 
        10'b0000111110: data <= 20'h003b9; 
        10'b0000111111: data <= 20'hffecf; 
        10'b0001000000: data <= 20'hffeb7; 
        10'b0001000001: data <= 20'h000ae; 
        10'b0001000010: data <= 20'hfff90; 
        10'b0001000011: data <= 20'hffdcb; 
        10'b0001000100: data <= 20'hff776; 
        10'b0001000101: data <= 20'hffc8d; 
        10'b0001000110: data <= 20'hffbde; 
        10'b0001000111: data <= 20'hffa26; 
        10'b0001001000: data <= 20'hffbbd; 
        10'b0001001001: data <= 20'hfff2a; 
        10'b0001001010: data <= 20'h00111; 
        10'b0001001011: data <= 20'h00301; 
        10'b0001001100: data <= 20'h003e7; 
        10'b0001001101: data <= 20'h00240; 
        10'b0001001110: data <= 20'h003ad; 
        10'b0001001111: data <= 20'h000fe; 
        10'b0001010000: data <= 20'h00165; 
        10'b0001010001: data <= 20'h0027d; 
        10'b0001010010: data <= 20'h00027; 
        10'b0001010011: data <= 20'h001bb; 
        10'b0001010100: data <= 20'h0034e; 
        10'b0001010101: data <= 20'h002f9; 
        10'b0001010110: data <= 20'h00126; 
        10'b0001010111: data <= 20'h001df; 
        10'b0001011000: data <= 20'h001f0; 
        10'b0001011001: data <= 20'h00007; 
        10'b0001011010: data <= 20'h0027b; 
        10'b0001011011: data <= 20'hffdcd; 
        10'b0001011100: data <= 20'hffcca; 
        10'b0001011101: data <= 20'hffe3f; 
        10'b0001011110: data <= 20'hff8a9; 
        10'b0001011111: data <= 20'hff750; 
        10'b0001100000: data <= 20'hff224; 
        10'b0001100001: data <= 20'hff2c7; 
        10'b0001100010: data <= 20'hff368; 
        10'b0001100011: data <= 20'hff0b8; 
        10'b0001100100: data <= 20'hff5cc; 
        10'b0001100101: data <= 20'hffae8; 
        10'b0001100110: data <= 20'h000c0; 
        10'b0001100111: data <= 20'h001a2; 
        10'b0001101000: data <= 20'h002f5; 
        10'b0001101001: data <= 20'h0045c; 
        10'b0001101010: data <= 20'h00124; 
        10'b0001101011: data <= 20'h0012a; 
        10'b0001101100: data <= 20'h0043e; 
        10'b0001101101: data <= 20'h00413; 
        10'b0001101110: data <= 20'h00143; 
        10'b0001101111: data <= 20'h00264; 
        10'b0001110000: data <= 20'h0041f; 
        10'b0001110001: data <= 20'h002bc; 
        10'b0001110010: data <= 20'h00314; 
        10'b0001110011: data <= 20'h002fd; 
        10'b0001110100: data <= 20'h001c7; 
        10'b0001110101: data <= 20'h00360; 
        10'b0001110110: data <= 20'hffd78; 
        10'b0001110111: data <= 20'hfff70; 
        10'b0001111000: data <= 20'hffad5; 
        10'b0001111001: data <= 20'hffba1; 
        10'b0001111010: data <= 20'hff392; 
        10'b0001111011: data <= 20'hff42d; 
        10'b0001111100: data <= 20'hfefd4; 
        10'b0001111101: data <= 20'hff292; 
        10'b0001111110: data <= 20'hfef83; 
        10'b0001111111: data <= 20'hff1e3; 
        10'b0010000000: data <= 20'hff924; 
        10'b0010000001: data <= 20'hff9e8; 
        10'b0010000010: data <= 20'hffc5a; 
        10'b0010000011: data <= 20'h00382; 
        10'b0010000100: data <= 20'h004d5; 
        10'b0010000101: data <= 20'h00585; 
        10'b0010000110: data <= 20'h00541; 
        10'b0010000111: data <= 20'h006f8; 
        10'b0010001000: data <= 20'h001ee; 
        10'b0010001001: data <= 20'h003ea; 
        10'b0010001010: data <= 20'h000ff; 
        10'b0010001011: data <= 20'h000a5; 
        10'b0010001100: data <= 20'h00431; 
        10'b0010001101: data <= 20'h0012c; 
        10'b0010001110: data <= 20'h002f6; 
        10'b0010001111: data <= 20'h000f8; 
        10'b0010010000: data <= 20'h002b7; 
        10'b0010010001: data <= 20'h0008c; 
        10'b0010010010: data <= 20'h001eb; 
        10'b0010010011: data <= 20'hffdac; 
        10'b0010010100: data <= 20'h000a0; 
        10'b0010010101: data <= 20'hffd4f; 
        10'b0010010110: data <= 20'hff6e9; 
        10'b0010010111: data <= 20'hff9fb; 
        10'b0010011000: data <= 20'hff5ac; 
        10'b0010011001: data <= 20'hff32e; 
        10'b0010011010: data <= 20'hff709; 
        10'b0010011011: data <= 20'hff89a; 
        10'b0010011100: data <= 20'hffec3; 
        10'b0010011101: data <= 20'h00123; 
        10'b0010011110: data <= 20'hffe3a; 
        10'b0010011111: data <= 20'h002fc; 
        10'b0010100000: data <= 20'h003a9; 
        10'b0010100001: data <= 20'h004f2; 
        10'b0010100010: data <= 20'h00b87; 
        10'b0010100011: data <= 20'h00d02; 
        10'b0010100100: data <= 20'h00714; 
        10'b0010100101: data <= 20'hfff4f; 
        10'b0010100110: data <= 20'h0012a; 
        10'b0010100111: data <= 20'h000b4; 
        10'b0010101000: data <= 20'h003e4; 
        10'b0010101001: data <= 20'h0044e; 
        10'b0010101010: data <= 20'h00148; 
        10'b0010101011: data <= 20'h00362; 
        10'b0010101100: data <= 20'h003af; 
        10'b0010101101: data <= 20'h00306; 
        10'b0010101110: data <= 20'h002ff; 
        10'b0010101111: data <= 20'hfffc3; 
        10'b0010110000: data <= 20'hfff52; 
        10'b0010110001: data <= 20'hffc6e; 
        10'b0010110010: data <= 20'hff8ca; 
        10'b0010110011: data <= 20'hff350; 
        10'b0010110100: data <= 20'hfecc7; 
        10'b0010110101: data <= 20'hfe946; 
        10'b0010110110: data <= 20'hfe844; 
        10'b0010110111: data <= 20'hfeb66; 
        10'b0010111000: data <= 20'hfeae4; 
        10'b0010111001: data <= 20'hff3a0; 
        10'b0010111010: data <= 20'hff336; 
        10'b0010111011: data <= 20'hffa3f; 
        10'b0010111100: data <= 20'hffc37; 
        10'b0010111101: data <= 20'hfffb6; 
        10'b0010111110: data <= 20'h01081; 
        10'b0010111111: data <= 20'h01156; 
        10'b0011000000: data <= 20'h006ac; 
        10'b0011000001: data <= 20'h0053b; 
        10'b0011000010: data <= 20'h003bd; 
        10'b0011000011: data <= 20'h00029; 
        10'b0011000100: data <= 20'h001d7; 
        10'b0011000101: data <= 20'h000f6; 
        10'b0011000110: data <= 20'h00153; 
        10'b0011000111: data <= 20'h00258; 
        10'b0011001000: data <= 20'h00158; 
        10'b0011001001: data <= 20'h00322; 
        10'b0011001010: data <= 20'hffe10; 
        10'b0011001011: data <= 20'hfffa6; 
        10'b0011001100: data <= 20'hffdda; 
        10'b0011001101: data <= 20'hffb21; 
        10'b0011001110: data <= 20'hff3b0; 
        10'b0011001111: data <= 20'hfeccd; 
        10'b0011010000: data <= 20'hfe70f; 
        10'b0011010001: data <= 20'hfee60; 
        10'b0011010010: data <= 20'hfe9f6; 
        10'b0011010011: data <= 20'hfe9cb; 
        10'b0011010100: data <= 20'hfe92a; 
        10'b0011010101: data <= 20'hff171; 
        10'b0011010110: data <= 20'hff116; 
        10'b0011010111: data <= 20'hff59e; 
        10'b0011011000: data <= 20'hff3ff; 
        10'b0011011001: data <= 20'hffa86; 
        10'b0011011010: data <= 20'h00a32; 
        10'b0011011011: data <= 20'h00dcb; 
        10'b0011011100: data <= 20'h0075c; 
        10'b0011011101: data <= 20'h00425; 
        10'b0011011110: data <= 20'h003e3; 
        10'b0011011111: data <= 20'h0024f; 
        10'b0011100000: data <= 20'h003bf; 
        10'b0011100001: data <= 20'h00325; 
        10'b0011100010: data <= 20'h00423; 
        10'b0011100011: data <= 20'h000cd; 
        10'b0011100100: data <= 20'h0013f; 
        10'b0011100101: data <= 20'h001b5; 
        10'b0011100110: data <= 20'h00125; 
        10'b0011100111: data <= 20'hfff01; 
        10'b0011101000: data <= 20'hff6b8; 
        10'b0011101001: data <= 20'hffb47; 
        10'b0011101010: data <= 20'hff9d5; 
        10'b0011101011: data <= 20'hff398; 
        10'b0011101100: data <= 20'hfedd5; 
        10'b0011101101: data <= 20'hff463; 
        10'b0011101110: data <= 20'hfe5ac; 
        10'b0011101111: data <= 20'hfe4f4; 
        10'b0011110000: data <= 20'hfeafa; 
        10'b0011110001: data <= 20'hff2d5; 
        10'b0011110010: data <= 20'hff42f; 
        10'b0011110011: data <= 20'hffc47; 
        10'b0011110100: data <= 20'hff8ca; 
        10'b0011110101: data <= 20'hff8e9; 
        10'b0011110110: data <= 20'h004b2; 
        10'b0011110111: data <= 20'h0073a; 
        10'b0011111000: data <= 20'h00583; 
        10'b0011111001: data <= 20'h00119; 
        10'b0011111010: data <= 20'h0017c; 
        10'b0011111011: data <= 20'h002b3; 
        10'b0011111100: data <= 20'h00474; 
        10'b0011111101: data <= 20'h003bf; 
        10'b0011111110: data <= 20'h0037f; 
        10'b0011111111: data <= 20'h000bc; 
        10'b0100000000: data <= 20'hffdae; 
        10'b0100000001: data <= 20'h00011; 
        10'b0100000010: data <= 20'hffa46; 
        10'b0100000011: data <= 20'hffbe4; 
        10'b0100000100: data <= 20'hffd55; 
        10'b0100000101: data <= 20'hfff1f; 
        10'b0100000110: data <= 20'hffcd2; 
        10'b0100000111: data <= 20'hffc2e; 
        10'b0100001000: data <= 20'hffc10; 
        10'b0100001001: data <= 20'hff586; 
        10'b0100001010: data <= 20'hfda0c; 
        10'b0100001011: data <= 20'hfe39b; 
        10'b0100001100: data <= 20'hff91d; 
        10'b0100001101: data <= 20'hffae9; 
        10'b0100001110: data <= 20'hffe6d; 
        10'b0100001111: data <= 20'h000d7; 
        10'b0100010000: data <= 20'hffc03; 
        10'b0100010001: data <= 20'hffc1b; 
        10'b0100010010: data <= 20'h001f7; 
        10'b0100010011: data <= 20'h00072; 
        10'b0100010100: data <= 20'hffb7b; 
        10'b0100010101: data <= 20'hffb4c; 
        10'b0100010110: data <= 20'hffdf6; 
        10'b0100010111: data <= 20'h00302; 
        10'b0100011000: data <= 20'h00260; 
        10'b0100011001: data <= 20'h001ae; 
        10'b0100011010: data <= 20'h001b3; 
        10'b0100011011: data <= 20'h00077; 
        10'b0100011100: data <= 20'h001c4; 
        10'b0100011101: data <= 20'hffae4; 
        10'b0100011110: data <= 20'hff78d; 
        10'b0100011111: data <= 20'hffbe5; 
        10'b0100100000: data <= 20'h00139; 
        10'b0100100001: data <= 20'h00ad1; 
        10'b0100100010: data <= 20'h0068c; 
        10'b0100100011: data <= 20'h004e5; 
        10'b0100100100: data <= 20'h005dc; 
        10'b0100100101: data <= 20'hff17c; 
        10'b0100100110: data <= 20'hfd7ec; 
        10'b0100100111: data <= 20'hff3c9; 
        10'b0100101000: data <= 20'h00166; 
        10'b0100101001: data <= 20'hffe33; 
        10'b0100101010: data <= 20'hffea1; 
        10'b0100101011: data <= 20'h0016b; 
        10'b0100101100: data <= 20'hff800; 
        10'b0100101101: data <= 20'hffab7; 
        10'b0100101110: data <= 20'hfff01; 
        10'b0100101111: data <= 20'hff74b; 
        10'b0100110000: data <= 20'hffb11; 
        10'b0100110001: data <= 20'hffcdf; 
        10'b0100110010: data <= 20'h0027f; 
        10'b0100110011: data <= 20'h0041f; 
        10'b0100110100: data <= 20'h002c6; 
        10'b0100110101: data <= 20'h002e4; 
        10'b0100110110: data <= 20'h00271; 
        10'b0100110111: data <= 20'hffe78; 
        10'b0100111000: data <= 20'hfff6f; 
        10'b0100111001: data <= 20'hffd25; 
        10'b0100111010: data <= 20'hffcfa; 
        10'b0100111011: data <= 20'h0028f; 
        10'b0100111100: data <= 20'h0082f; 
        10'b0100111101: data <= 20'h00dca; 
        10'b0100111110: data <= 20'h01301; 
        10'b0100111111: data <= 20'h00c17; 
        10'b0101000000: data <= 20'h00da5; 
        10'b0101000001: data <= 20'hfe9c4; 
        10'b0101000010: data <= 20'hfe1d2; 
        10'b0101000011: data <= 20'h003eb; 
        10'b0101000100: data <= 20'h00f9b; 
        10'b0101000101: data <= 20'h002a1; 
        10'b0101000110: data <= 20'hfff19; 
        10'b0101000111: data <= 20'hffd7f; 
        10'b0101001000: data <= 20'hff776; 
        10'b0101001001: data <= 20'hff8b4; 
        10'b0101001010: data <= 20'hffc47; 
        10'b0101001011: data <= 20'hff93f; 
        10'b0101001100: data <= 20'hff87f; 
        10'b0101001101: data <= 20'hfff94; 
        10'b0101001110: data <= 20'hfffbf; 
        10'b0101001111: data <= 20'h00109; 
        10'b0101010000: data <= 20'h00319; 
        10'b0101010001: data <= 20'h002b7; 
        10'b0101010010: data <= 20'h0014a; 
        10'b0101010011: data <= 20'h001dc; 
        10'b0101010100: data <= 20'hfffcf; 
        10'b0101010101: data <= 20'hffd36; 
        10'b0101010110: data <= 20'h00807; 
        10'b0101010111: data <= 20'h00d3b; 
        10'b0101011000: data <= 20'h0147f; 
        10'b0101011001: data <= 20'h011f5; 
        10'b0101011010: data <= 20'h01dde; 
        10'b0101011011: data <= 20'h021d7; 
        10'b0101011100: data <= 20'h01ffd; 
        10'b0101011101: data <= 20'hfff78; 
        10'b0101011110: data <= 20'hff016; 
        10'b0101011111: data <= 20'h00c85; 
        10'b0101100000: data <= 20'h01455; 
        10'b0101100001: data <= 20'h0024f; 
        10'b0101100010: data <= 20'h000db; 
        10'b0101100011: data <= 20'h002c7; 
        10'b0101100100: data <= 20'hfff83; 
        10'b0101100101: data <= 20'h00099; 
        10'b0101100110: data <= 20'hfff18; 
        10'b0101100111: data <= 20'hffb84; 
        10'b0101101000: data <= 20'hffbfe; 
        10'b0101101001: data <= 20'hffedf; 
        10'b0101101010: data <= 20'h0046b; 
        10'b0101101011: data <= 20'h0028e; 
        10'b0101101100: data <= 20'h0007c; 
        10'b0101101101: data <= 20'h002e9; 
        10'b0101101110: data <= 20'h00067; 
        10'b0101101111: data <= 20'h00138; 
        10'b0101110000: data <= 20'h0036f; 
        10'b0101110001: data <= 20'h009af; 
        10'b0101110010: data <= 20'h013b4; 
        10'b0101110011: data <= 20'h016dd; 
        10'b0101110100: data <= 20'h01a49; 
        10'b0101110101: data <= 20'h015f6; 
        10'b0101110110: data <= 20'h019a1; 
        10'b0101110111: data <= 20'h029c3; 
        10'b0101111000: data <= 20'h01fa8; 
        10'b0101111001: data <= 20'h0007a; 
        10'b0101111010: data <= 20'hffb81; 
        10'b0101111011: data <= 20'h00eab; 
        10'b0101111100: data <= 20'h00f11; 
        10'b0101111101: data <= 20'h010bc; 
        10'b0101111110: data <= 20'h00b8a; 
        10'b0101111111: data <= 20'h00531; 
        10'b0110000000: data <= 20'h00b8f; 
        10'b0110000001: data <= 20'h00882; 
        10'b0110000010: data <= 20'h0040e; 
        10'b0110000011: data <= 20'hffda3; 
        10'b0110000100: data <= 20'hffded; 
        10'b0110000101: data <= 20'h0003c; 
        10'b0110000110: data <= 20'h0038c; 
        10'b0110000111: data <= 20'h0028a; 
        10'b0110001000: data <= 20'h00073; 
        10'b0110001001: data <= 20'h003a0; 
        10'b0110001010: data <= 20'h0004a; 
        10'b0110001011: data <= 20'h00444; 
        10'b0110001100: data <= 20'h00892; 
        10'b0110001101: data <= 20'h01142; 
        10'b0110001110: data <= 20'h017fd; 
        10'b0110001111: data <= 20'h01a41; 
        10'b0110010000: data <= 20'h0139d; 
        10'b0110010001: data <= 20'h012bf; 
        10'b0110010010: data <= 20'h01697; 
        10'b0110010011: data <= 20'h01b60; 
        10'b0110010100: data <= 20'h013ee; 
        10'b0110010101: data <= 20'h001a7; 
        10'b0110010110: data <= 20'hffd19; 
        10'b0110010111: data <= 20'h0054c; 
        10'b0110011000: data <= 20'h010c8; 
        10'b0110011001: data <= 20'h01b93; 
        10'b0110011010: data <= 20'h012bb; 
        10'b0110011011: data <= 20'h01137; 
        10'b0110011100: data <= 20'h0099c; 
        10'b0110011101: data <= 20'h00676; 
        10'b0110011110: data <= 20'h0021a; 
        10'b0110011111: data <= 20'h00130; 
        10'b0110100000: data <= 20'hfff51; 
        10'b0110100001: data <= 20'h00127; 
        10'b0110100010: data <= 20'h00229; 
        10'b0110100011: data <= 20'h00105; 
        10'b0110100100: data <= 20'h002fe; 
        10'b0110100101: data <= 20'h0044b; 
        10'b0110100110: data <= 20'h002c2; 
        10'b0110100111: data <= 20'h0038d; 
        10'b0110101000: data <= 20'h007c0; 
        10'b0110101001: data <= 20'h008ca; 
        10'b0110101010: data <= 20'h00da9; 
        10'b0110101011: data <= 20'h00c94; 
        10'b0110101100: data <= 20'h0143e; 
        10'b0110101101: data <= 20'h01164; 
        10'b0110101110: data <= 20'h00c1a; 
        10'b0110101111: data <= 20'h008ca; 
        10'b0110110000: data <= 20'h00a62; 
        10'b0110110001: data <= 20'h0020d; 
        10'b0110110010: data <= 20'h00854; 
        10'b0110110011: data <= 20'h00ba6; 
        10'b0110110100: data <= 20'h0182f; 
        10'b0110110101: data <= 20'h0157d; 
        10'b0110110110: data <= 20'h00f5c; 
        10'b0110110111: data <= 20'h00919; 
        10'b0110111000: data <= 20'hffd8d; 
        10'b0110111001: data <= 20'h00360; 
        10'b0110111010: data <= 20'h0061b; 
        10'b0110111011: data <= 20'h000a5; 
        10'b0110111100: data <= 20'hffc53; 
        10'b0110111101: data <= 20'h001ef; 
        10'b0110111110: data <= 20'h0007f; 
        10'b0110111111: data <= 20'h00138; 
        10'b0111000000: data <= 20'h00154; 
        10'b0111000001: data <= 20'h00007; 
        10'b0111000010: data <= 20'h00028; 
        10'b0111000011: data <= 20'hfff78; 
        10'b0111000100: data <= 20'h0021b; 
        10'b0111000101: data <= 20'h00530; 
        10'b0111000110: data <= 20'h00874; 
        10'b0111000111: data <= 20'h00ec2; 
        10'b0111001000: data <= 20'h0157c; 
        10'b0111001001: data <= 20'h00f4f; 
        10'b0111001010: data <= 20'h00419; 
        10'b0111001011: data <= 20'hfff71; 
        10'b0111001100: data <= 20'h00435; 
        10'b0111001101: data <= 20'h00540; 
        10'b0111001110: data <= 20'h013b8; 
        10'b0111001111: data <= 20'h01b44; 
        10'b0111010000: data <= 20'h01c15; 
        10'b0111010001: data <= 20'h01754; 
        10'b0111010010: data <= 20'h00fcb; 
        10'b0111010011: data <= 20'h001fb; 
        10'b0111010100: data <= 20'h006a0; 
        10'b0111010101: data <= 20'h00968; 
        10'b0111010110: data <= 20'h00233; 
        10'b0111010111: data <= 20'hffe73; 
        10'b0111011000: data <= 20'hfff93; 
        10'b0111011001: data <= 20'h000ea; 
        10'b0111011010: data <= 20'h001b2; 
        10'b0111011011: data <= 20'h001c8; 
        10'b0111011100: data <= 20'h00194; 
        10'b0111011101: data <= 20'h0019d; 
        10'b0111011110: data <= 20'h00337; 
        10'b0111011111: data <= 20'hffff3; 
        10'b0111100000: data <= 20'hffdbf; 
        10'b0111100001: data <= 20'hffb5c; 
        10'b0111100010: data <= 20'h002bf; 
        10'b0111100011: data <= 20'h00bb4; 
        10'b0111100100: data <= 20'h01693; 
        10'b0111100101: data <= 20'h01392; 
        10'b0111100110: data <= 20'h00717; 
        10'b0111100111: data <= 20'h00594; 
        10'b0111101000: data <= 20'h00813; 
        10'b0111101001: data <= 20'h0135d; 
        10'b0111101010: data <= 20'h01ffd; 
        10'b0111101011: data <= 20'h01951; 
        10'b0111101100: data <= 20'h0152d; 
        10'b0111101101: data <= 20'h0068b; 
        10'b0111101110: data <= 20'h00103; 
        10'b0111101111: data <= 20'hff8ea; 
        10'b0111110000: data <= 20'h0021f; 
        10'b0111110001: data <= 20'h000c7; 
        10'b0111110010: data <= 20'hffbab; 
        10'b0111110011: data <= 20'hffe23; 
        10'b0111110100: data <= 20'hffd2e; 
        10'b0111110101: data <= 20'hffe63; 
        10'b0111110110: data <= 20'h002d9; 
        10'b0111110111: data <= 20'h0037b; 
        10'b0111111000: data <= 20'h001bf; 
        10'b0111111001: data <= 20'h002ac; 
        10'b0111111010: data <= 20'h00256; 
        10'b0111111011: data <= 20'h00059; 
        10'b0111111100: data <= 20'hffd46; 
        10'b0111111101: data <= 20'hffa44; 
        10'b0111111110: data <= 20'hff957; 
        10'b0111111111: data <= 20'hfffdf; 
        10'b1000000000: data <= 20'h005c6; 
        10'b1000000001: data <= 20'h00152; 
        10'b1000000010: data <= 20'hffb4c; 
        10'b1000000011: data <= 20'hffd38; 
        10'b1000000100: data <= 20'h00762; 
        10'b1000000101: data <= 20'h00852; 
        10'b1000000110: data <= 20'h00e0f; 
        10'b1000000111: data <= 20'h00c07; 
        10'b1000001000: data <= 20'h00648; 
        10'b1000001001: data <= 20'hff645; 
        10'b1000001010: data <= 20'hff6c9; 
        10'b1000001011: data <= 20'hff27c; 
        10'b1000001100: data <= 20'hff7fc; 
        10'b1000001101: data <= 20'hff7af; 
        10'b1000001110: data <= 20'hff4ed; 
        10'b1000001111: data <= 20'hff76b; 
        10'b1000010000: data <= 20'hffdc3; 
        10'b1000010001: data <= 20'hffed0; 
        10'b1000010010: data <= 20'h00107; 
        10'b1000010011: data <= 20'h00024; 
        10'b1000010100: data <= 20'h001b0; 
        10'b1000010101: data <= 20'h00320; 
        10'b1000010110: data <= 20'h00130; 
        10'b1000010111: data <= 20'h000b7; 
        10'b1000011000: data <= 20'hff9d0; 
        10'b1000011001: data <= 20'hff850; 
        10'b1000011010: data <= 20'hff5d8; 
        10'b1000011011: data <= 20'hff0be; 
        10'b1000011100: data <= 20'hfeeca; 
        10'b1000011101: data <= 20'hfeda9; 
        10'b1000011110: data <= 20'hfea5c; 
        10'b1000011111: data <= 20'hfeb4d; 
        10'b1000100000: data <= 20'hfedac; 
        10'b1000100001: data <= 20'hff542; 
        10'b1000100010: data <= 20'hffccf; 
        10'b1000100011: data <= 20'h002ca; 
        10'b1000100100: data <= 20'hff7ab; 
        10'b1000100101: data <= 20'hff8d4; 
        10'b1000100110: data <= 20'hff72a; 
        10'b1000100111: data <= 20'hff3cf; 
        10'b1000101000: data <= 20'hff25f; 
        10'b1000101001: data <= 20'hff372; 
        10'b1000101010: data <= 20'hff33e; 
        10'b1000101011: data <= 20'hff75f; 
        10'b1000101100: data <= 20'hffdba; 
        10'b1000101101: data <= 20'h001b5; 
        10'b1000101110: data <= 20'h00305; 
        10'b1000101111: data <= 20'h002c3; 
        10'b1000110000: data <= 20'h0047f; 
        10'b1000110001: data <= 20'h0042a; 
        10'b1000110010: data <= 20'h00134; 
        10'b1000110011: data <= 20'h000b7; 
        10'b1000110100: data <= 20'hffafb; 
        10'b1000110101: data <= 20'hff769; 
        10'b1000110110: data <= 20'hff386; 
        10'b1000110111: data <= 20'hfebb1; 
        10'b1000111000: data <= 20'hfe7dc; 
        10'b1000111001: data <= 20'hfe66c; 
        10'b1000111010: data <= 20'hfe5f4; 
        10'b1000111011: data <= 20'hfecee; 
        10'b1000111100: data <= 20'hff095; 
        10'b1000111101: data <= 20'hfeec3; 
        10'b1000111110: data <= 20'hff52b; 
        10'b1000111111: data <= 20'hffa5b; 
        10'b1001000000: data <= 20'hffe0d; 
        10'b1001000001: data <= 20'hffee9; 
        10'b1001000010: data <= 20'hffb86; 
        10'b1001000011: data <= 20'hff64c; 
        10'b1001000100: data <= 20'hff97a; 
        10'b1001000101: data <= 20'hff89e; 
        10'b1001000110: data <= 20'hff717; 
        10'b1001000111: data <= 20'hffb6e; 
        10'b1001001000: data <= 20'hffb9d; 
        10'b1001001001: data <= 20'h00053; 
        10'b1001001010: data <= 20'h0010f; 
        10'b1001001011: data <= 20'h00302; 
        10'b1001001100: data <= 20'h000d5; 
        10'b1001001101: data <= 20'h0014f; 
        10'b1001001110: data <= 20'h00058; 
        10'b1001001111: data <= 20'h00099; 
        10'b1001010000: data <= 20'hffff3; 
        10'b1001010001: data <= 20'hffb1b; 
        10'b1001010010: data <= 20'hff3b5; 
        10'b1001010011: data <= 20'hfeec6; 
        10'b1001010100: data <= 20'hff07f; 
        10'b1001010101: data <= 20'hfee5e; 
        10'b1001010110: data <= 20'hff0a7; 
        10'b1001010111: data <= 20'hff49a; 
        10'b1001011000: data <= 20'hff685; 
        10'b1001011001: data <= 20'hff738; 
        10'b1001011010: data <= 20'hff5f1; 
        10'b1001011011: data <= 20'hffb59; 
        10'b1001011100: data <= 20'hff9cc; 
        10'b1001011101: data <= 20'h0011e; 
        10'b1001011110: data <= 20'hffe26; 
        10'b1001011111: data <= 20'h00056; 
        10'b1001100000: data <= 20'hfff31; 
        10'b1001100001: data <= 20'hff9f6; 
        10'b1001100010: data <= 20'hffae3; 
        10'b1001100011: data <= 20'hfff0f; 
        10'b1001100100: data <= 20'hfffd6; 
        10'b1001100101: data <= 20'h001dc; 
        10'b1001100110: data <= 20'h0027f; 
        10'b1001100111: data <= 20'h00268; 
        10'b1001101000: data <= 20'h0022b; 
        10'b1001101001: data <= 20'h00285; 
        10'b1001101010: data <= 20'h00101; 
        10'b1001101011: data <= 20'h002c2; 
        10'b1001101100: data <= 20'hfff5a; 
        10'b1001101101: data <= 20'hffd64; 
        10'b1001101110: data <= 20'hffaed; 
        10'b1001101111: data <= 20'hff7a0; 
        10'b1001110000: data <= 20'hff4af; 
        10'b1001110001: data <= 20'hff920; 
        10'b1001110010: data <= 20'hff8eb; 
        10'b1001110011: data <= 20'hffb16; 
        10'b1001110100: data <= 20'hffad2; 
        10'b1001110101: data <= 20'hffb8d; 
        10'b1001110110: data <= 20'hffa72; 
        10'b1001110111: data <= 20'hffc96; 
        10'b1001111000: data <= 20'hffcba; 
        10'b1001111001: data <= 20'h0012e; 
        10'b1001111010: data <= 20'h00505; 
        10'b1001111011: data <= 20'h00831; 
        10'b1001111100: data <= 20'h00649; 
        10'b1001111101: data <= 20'h0041f; 
        10'b1001111110: data <= 20'hffd46; 
        10'b1001111111: data <= 20'hffd52; 
        10'b1010000000: data <= 20'hfffe6; 
        10'b1010000001: data <= 20'h001cc; 
        10'b1010000010: data <= 20'h00049; 
        10'b1010000011: data <= 20'h00161; 
        10'b1010000100: data <= 20'h00167; 
        10'b1010000101: data <= 20'h00019; 
        10'b1010000110: data <= 20'h0013e; 
        10'b1010000111: data <= 20'h00274; 
        10'b1010001000: data <= 20'h00163; 
        10'b1010001001: data <= 20'h001b4; 
        10'b1010001010: data <= 20'hffd4c; 
        10'b1010001011: data <= 20'hffcff; 
        10'b1010001100: data <= 20'hffbef; 
        10'b1010001101: data <= 20'h001e5; 
        10'b1010001110: data <= 20'hffba0; 
        10'b1010001111: data <= 20'h000b5; 
        10'b1010010000: data <= 20'hffb7a; 
        10'b1010010001: data <= 20'hffc72; 
        10'b1010010010: data <= 20'hffc87; 
        10'b1010010011: data <= 20'hfffbe; 
        10'b1010010100: data <= 20'h00128; 
        10'b1010010101: data <= 20'h0030f; 
        10'b1010010110: data <= 20'h0096c; 
        10'b1010010111: data <= 20'h00932; 
        10'b1010011000: data <= 20'h007d6; 
        10'b1010011001: data <= 20'h0037e; 
        10'b1010011010: data <= 20'hffeb5; 
        10'b1010011011: data <= 20'h00110; 
        10'b1010011100: data <= 20'h00214; 
        10'b1010011101: data <= 20'h002d8; 
        10'b1010011110: data <= 20'h000ee; 
        10'b1010011111: data <= 20'h0038a; 
        10'b1010100000: data <= 20'h002ad; 
        10'b1010100001: data <= 20'h003d3; 
        10'b1010100010: data <= 20'h001cf; 
        10'b1010100011: data <= 20'h00308; 
        10'b1010100100: data <= 20'h000b6; 
        10'b1010100101: data <= 20'h00252; 
        10'b1010100110: data <= 20'h000e2; 
        10'b1010100111: data <= 20'hffbb1; 
        10'b1010101000: data <= 20'hffb9a; 
        10'b1010101001: data <= 20'hffe99; 
        10'b1010101010: data <= 20'hffb56; 
        10'b1010101011: data <= 20'hfff3d; 
        10'b1010101100: data <= 20'hffca6; 
        10'b1010101101: data <= 20'hffce9; 
        10'b1010101110: data <= 20'hffa50; 
        10'b1010101111: data <= 20'hff99e; 
        10'b1010110000: data <= 20'hffd3f; 
        10'b1010110001: data <= 20'hffe92; 
        10'b1010110010: data <= 20'h00080; 
        10'b1010110011: data <= 20'h004f4; 
        10'b1010110100: data <= 20'h0039e; 
        10'b1010110101: data <= 20'hffe85; 
        10'b1010110110: data <= 20'hfff93; 
        10'b1010110111: data <= 20'h001ea; 
        10'b1010111000: data <= 20'h00326; 
        10'b1010111001: data <= 20'h00081; 
        10'b1010111010: data <= 20'h000d1; 
        10'b1010111011: data <= 20'h002ba; 
        10'b1010111100: data <= 20'h00401; 
        10'b1010111101: data <= 20'h003e2; 
        10'b1010111110: data <= 20'h0038c; 
        10'b1010111111: data <= 20'h000cb; 
        10'b1011000000: data <= 20'h00392; 
        10'b1011000001: data <= 20'h0002b; 
        10'b1011000010: data <= 20'hffd73; 
        10'b1011000011: data <= 20'hffbd9; 
        10'b1011000100: data <= 20'hff9c1; 
        10'b1011000101: data <= 20'hff96e; 
        10'b1011000110: data <= 20'hff536; 
        10'b1011000111: data <= 20'hff3d4; 
        10'b1011001000: data <= 20'hff481; 
        10'b1011001001: data <= 20'hff491; 
        10'b1011001010: data <= 20'hff649; 
        10'b1011001011: data <= 20'hff5b7; 
        10'b1011001100: data <= 20'hff2b1; 
        10'b1011001101: data <= 20'hff0d5; 
        10'b1011001110: data <= 20'hff261; 
        10'b1011001111: data <= 20'hff889; 
        10'b1011010000: data <= 20'hff92c; 
        10'b1011010001: data <= 20'hffd89; 
        10'b1011010010: data <= 20'h00027; 
        10'b1011010011: data <= 20'h0029d; 
        10'b1011010100: data <= 20'h00032; 
        10'b1011010101: data <= 20'h003a1; 
        10'b1011010110: data <= 20'h00174; 
        10'b1011010111: data <= 20'h00151; 
        10'b1011011000: data <= 20'h001df; 
        10'b1011011001: data <= 20'h002b3; 
        10'b1011011010: data <= 20'h0009c; 
        10'b1011011011: data <= 20'h001cc; 
        10'b1011011100: data <= 20'hfffd2; 
        10'b1011011101: data <= 20'hfff62; 
        10'b1011011110: data <= 20'h00115; 
        10'b1011011111: data <= 20'h000c8; 
        10'b1011100000: data <= 20'hfff2d; 
        10'b1011100001: data <= 20'hffc39; 
        10'b1011100010: data <= 20'hff6e4; 
        10'b1011100011: data <= 20'hff80d; 
        10'b1011100100: data <= 20'hff6e8; 
        10'b1011100101: data <= 20'hff3a6; 
        10'b1011100110: data <= 20'hff281; 
        10'b1011100111: data <= 20'hff57f; 
        10'b1011101000: data <= 20'hff40a; 
        10'b1011101001: data <= 20'hff5d8; 
        10'b1011101010: data <= 20'hff7a9; 
        10'b1011101011: data <= 20'hffb08; 
        10'b1011101100: data <= 20'hffe2e; 
        10'b1011101101: data <= 20'h002b1; 
        10'b1011101110: data <= 20'h002ab; 
        10'b1011101111: data <= 20'h00056; 
        10'b1011110000: data <= 20'h001c0; 
        10'b1011110001: data <= 20'h00049; 
        10'b1011110010: data <= 20'h0044b; 
        10'b1011110011: data <= 20'h001e1; 
        10'b1011110100: data <= 20'h0029b; 
        10'b1011110101: data <= 20'h00062; 
        10'b1011110110: data <= 20'h00094; 
        10'b1011110111: data <= 20'h00420; 
        10'b1011111000: data <= 20'h0018c; 
        10'b1011111001: data <= 20'h00370; 
        10'b1011111010: data <= 20'h00195; 
        10'b1011111011: data <= 20'h00435; 
        10'b1011111100: data <= 20'hffffe; 
        10'b1011111101: data <= 20'h001d0; 
        10'b1011111110: data <= 20'h000ee; 
        10'b1011111111: data <= 20'hfff6a; 
        10'b1100000000: data <= 20'hfff92; 
        10'b1100000001: data <= 20'h00027; 
        10'b1100000010: data <= 20'hffe40; 
        10'b1100000011: data <= 20'h00356; 
        10'b1100000100: data <= 20'hfff25; 
        10'b1100000101: data <= 20'hfff06; 
        10'b1100000110: data <= 20'hfffab; 
        10'b1100000111: data <= 20'h001c2; 
        10'b1100001000: data <= 20'h0015a; 
        10'b1100001001: data <= 20'h00158; 
        10'b1100001010: data <= 20'h0016d; 
        10'b1100001011: data <= 20'h00270; 
        10'b1100001100: data <= 20'h00255; 
        10'b1100001101: data <= 20'h00314; 
        10'b1100001110: data <= 20'h00235; 
        10'b1100001111: data <= 20'h00177; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 15) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 21'h1ffffe; 
        10'b0000000001: data <= 21'h000120; 
        10'b0000000010: data <= 21'h00078f; 
        10'b0000000011: data <= 21'h00078d; 
        10'b0000000100: data <= 21'h000023; 
        10'b0000000101: data <= 21'h000025; 
        10'b0000000110: data <= 21'h0005eb; 
        10'b0000000111: data <= 21'h00019e; 
        10'b0000001000: data <= 21'h000080; 
        10'b0000001001: data <= 21'h00011e; 
        10'b0000001010: data <= 21'h000038; 
        10'b0000001011: data <= 21'h00056f; 
        10'b0000001100: data <= 21'h000727; 
        10'b0000001101: data <= 21'h000412; 
        10'b0000001110: data <= 21'h000542; 
        10'b0000001111: data <= 21'h000095; 
        10'b0000010000: data <= 21'h0004ec; 
        10'b0000010001: data <= 21'h0006c0; 
        10'b0000010010: data <= 21'h00016c; 
        10'b0000010011: data <= 21'h000573; 
        10'b0000010100: data <= 21'h000068; 
        10'b0000010101: data <= 21'h00033d; 
        10'b0000010110: data <= 21'h000748; 
        10'b0000010111: data <= 21'h0000ba; 
        10'b0000011000: data <= 21'h000747; 
        10'b0000011001: data <= 21'h000127; 
        10'b0000011010: data <= 21'h0007f6; 
        10'b0000011011: data <= 21'h000347; 
        10'b0000011100: data <= 21'h000215; 
        10'b0000011101: data <= 21'h0003b9; 
        10'b0000011110: data <= 21'h1ffff0; 
        10'b0000011111: data <= 21'h0000a0; 
        10'b0000100000: data <= 21'h0003a4; 
        10'b0000100001: data <= 21'h0008c8; 
        10'b0000100010: data <= 21'h0001d1; 
        10'b0000100011: data <= 21'h1ffe98; 
        10'b0000100100: data <= 21'h0004e0; 
        10'b0000100101: data <= 21'h00002d; 
        10'b0000100110: data <= 21'h000346; 
        10'b0000100111: data <= 21'h1ffd71; 
        10'b0000101000: data <= 21'h000241; 
        10'b0000101001: data <= 21'h1ffc7b; 
        10'b0000101010: data <= 21'h000030; 
        10'b0000101011: data <= 21'h0004d3; 
        10'b0000101100: data <= 21'h0005af; 
        10'b0000101101: data <= 21'h0001ac; 
        10'b0000101110: data <= 21'h000017; 
        10'b0000101111: data <= 21'h00016e; 
        10'b0000110000: data <= 21'h00061e; 
        10'b0000110001: data <= 21'h1fffdb; 
        10'b0000110010: data <= 21'h1fffcc; 
        10'b0000110011: data <= 21'h000080; 
        10'b0000110100: data <= 21'h00056a; 
        10'b0000110101: data <= 21'h0005bb; 
        10'b0000110110: data <= 21'h00015b; 
        10'b0000110111: data <= 21'h0005b7; 
        10'b0000111000: data <= 21'h00068e; 
        10'b0000111001: data <= 21'h000443; 
        10'b0000111010: data <= 21'h000678; 
        10'b0000111011: data <= 21'h0006a2; 
        10'b0000111100: data <= 21'h000649; 
        10'b0000111101: data <= 21'h00059b; 
        10'b0000111110: data <= 21'h000772; 
        10'b0000111111: data <= 21'h1ffd9e; 
        10'b0001000000: data <= 21'h1ffd6f; 
        10'b0001000001: data <= 21'h00015b; 
        10'b0001000010: data <= 21'h1fff20; 
        10'b0001000011: data <= 21'h1ffb96; 
        10'b0001000100: data <= 21'h1feeec; 
        10'b0001000101: data <= 21'h1ff91a; 
        10'b0001000110: data <= 21'h1ff7bc; 
        10'b0001000111: data <= 21'h1ff44c; 
        10'b0001001000: data <= 21'h1ff77b; 
        10'b0001001001: data <= 21'h1ffe53; 
        10'b0001001010: data <= 21'h000222; 
        10'b0001001011: data <= 21'h000602; 
        10'b0001001100: data <= 21'h0007ce; 
        10'b0001001101: data <= 21'h000480; 
        10'b0001001110: data <= 21'h00075a; 
        10'b0001001111: data <= 21'h0001fb; 
        10'b0001010000: data <= 21'h0002c9; 
        10'b0001010001: data <= 21'h0004f9; 
        10'b0001010010: data <= 21'h00004f; 
        10'b0001010011: data <= 21'h000376; 
        10'b0001010100: data <= 21'h00069d; 
        10'b0001010101: data <= 21'h0005f1; 
        10'b0001010110: data <= 21'h00024b; 
        10'b0001010111: data <= 21'h0003bd; 
        10'b0001011000: data <= 21'h0003e0; 
        10'b0001011001: data <= 21'h00000d; 
        10'b0001011010: data <= 21'h0004f6; 
        10'b0001011011: data <= 21'h1ffb9a; 
        10'b0001011100: data <= 21'h1ff993; 
        10'b0001011101: data <= 21'h1ffc7f; 
        10'b0001011110: data <= 21'h1ff151; 
        10'b0001011111: data <= 21'h1feea0; 
        10'b0001100000: data <= 21'h1fe447; 
        10'b0001100001: data <= 21'h1fe58d; 
        10'b0001100010: data <= 21'h1fe6d1; 
        10'b0001100011: data <= 21'h1fe170; 
        10'b0001100100: data <= 21'h1feb99; 
        10'b0001100101: data <= 21'h1ff5cf; 
        10'b0001100110: data <= 21'h00017f; 
        10'b0001100111: data <= 21'h000345; 
        10'b0001101000: data <= 21'h0005eb; 
        10'b0001101001: data <= 21'h0008b8; 
        10'b0001101010: data <= 21'h000248; 
        10'b0001101011: data <= 21'h000254; 
        10'b0001101100: data <= 21'h00087c; 
        10'b0001101101: data <= 21'h000827; 
        10'b0001101110: data <= 21'h000285; 
        10'b0001101111: data <= 21'h0004c8; 
        10'b0001110000: data <= 21'h00083e; 
        10'b0001110001: data <= 21'h000578; 
        10'b0001110010: data <= 21'h000629; 
        10'b0001110011: data <= 21'h0005f9; 
        10'b0001110100: data <= 21'h00038e; 
        10'b0001110101: data <= 21'h0006c1; 
        10'b0001110110: data <= 21'h1ffaef; 
        10'b0001110111: data <= 21'h1ffedf; 
        10'b0001111000: data <= 21'h1ff5aa; 
        10'b0001111001: data <= 21'h1ff742; 
        10'b0001111010: data <= 21'h1fe725; 
        10'b0001111011: data <= 21'h1fe85a; 
        10'b0001111100: data <= 21'h1fdfa9; 
        10'b0001111101: data <= 21'h1fe524; 
        10'b0001111110: data <= 21'h1fdf06; 
        10'b0001111111: data <= 21'h1fe3c6; 
        10'b0010000000: data <= 21'h1ff249; 
        10'b0010000001: data <= 21'h1ff3cf; 
        10'b0010000010: data <= 21'h1ff8b5; 
        10'b0010000011: data <= 21'h000704; 
        10'b0010000100: data <= 21'h0009aa; 
        10'b0010000101: data <= 21'h000b0a; 
        10'b0010000110: data <= 21'h000a82; 
        10'b0010000111: data <= 21'h000df0; 
        10'b0010001000: data <= 21'h0003dd; 
        10'b0010001001: data <= 21'h0007d5; 
        10'b0010001010: data <= 21'h0001fe; 
        10'b0010001011: data <= 21'h000149; 
        10'b0010001100: data <= 21'h000863; 
        10'b0010001101: data <= 21'h000259; 
        10'b0010001110: data <= 21'h0005ec; 
        10'b0010001111: data <= 21'h0001f0; 
        10'b0010010000: data <= 21'h00056d; 
        10'b0010010001: data <= 21'h000118; 
        10'b0010010010: data <= 21'h0003d7; 
        10'b0010010011: data <= 21'h1ffb57; 
        10'b0010010100: data <= 21'h000140; 
        10'b0010010101: data <= 21'h1ffa9e; 
        10'b0010010110: data <= 21'h1fedd2; 
        10'b0010010111: data <= 21'h1ff3f5; 
        10'b0010011000: data <= 21'h1feb58; 
        10'b0010011001: data <= 21'h1fe65d; 
        10'b0010011010: data <= 21'h1fee12; 
        10'b0010011011: data <= 21'h1ff134; 
        10'b0010011100: data <= 21'h1ffd86; 
        10'b0010011101: data <= 21'h000245; 
        10'b0010011110: data <= 21'h1ffc74; 
        10'b0010011111: data <= 21'h0005f8; 
        10'b0010100000: data <= 21'h000753; 
        10'b0010100001: data <= 21'h0009e5; 
        10'b0010100010: data <= 21'h00170f; 
        10'b0010100011: data <= 21'h001a04; 
        10'b0010100100: data <= 21'h000e27; 
        10'b0010100101: data <= 21'h1ffe9d; 
        10'b0010100110: data <= 21'h000253; 
        10'b0010100111: data <= 21'h000167; 
        10'b0010101000: data <= 21'h0007c8; 
        10'b0010101001: data <= 21'h00089b; 
        10'b0010101010: data <= 21'h000290; 
        10'b0010101011: data <= 21'h0006c4; 
        10'b0010101100: data <= 21'h00075d; 
        10'b0010101101: data <= 21'h00060d; 
        10'b0010101110: data <= 21'h0005ff; 
        10'b0010101111: data <= 21'h1fff86; 
        10'b0010110000: data <= 21'h1ffea5; 
        10'b0010110001: data <= 21'h1ff8dc; 
        10'b0010110010: data <= 21'h1ff194; 
        10'b0010110011: data <= 21'h1fe6a0; 
        10'b0010110100: data <= 21'h1fd98e; 
        10'b0010110101: data <= 21'h1fd28d; 
        10'b0010110110: data <= 21'h1fd089; 
        10'b0010110111: data <= 21'h1fd6cc; 
        10'b0010111000: data <= 21'h1fd5c8; 
        10'b0010111001: data <= 21'h1fe740; 
        10'b0010111010: data <= 21'h1fe66c; 
        10'b0010111011: data <= 21'h1ff47f; 
        10'b0010111100: data <= 21'h1ff86e; 
        10'b0010111101: data <= 21'h1fff6c; 
        10'b0010111110: data <= 21'h002101; 
        10'b0010111111: data <= 21'h0022ad; 
        10'b0011000000: data <= 21'h000d57; 
        10'b0011000001: data <= 21'h000a75; 
        10'b0011000010: data <= 21'h000779; 
        10'b0011000011: data <= 21'h000052; 
        10'b0011000100: data <= 21'h0003ae; 
        10'b0011000101: data <= 21'h0001ed; 
        10'b0011000110: data <= 21'h0002a6; 
        10'b0011000111: data <= 21'h0004af; 
        10'b0011001000: data <= 21'h0002af; 
        10'b0011001001: data <= 21'h000644; 
        10'b0011001010: data <= 21'h1ffc20; 
        10'b0011001011: data <= 21'h1fff4b; 
        10'b0011001100: data <= 21'h1ffbb5; 
        10'b0011001101: data <= 21'h1ff642; 
        10'b0011001110: data <= 21'h1fe760; 
        10'b0011001111: data <= 21'h1fd99a; 
        10'b0011010000: data <= 21'h1fce1f; 
        10'b0011010001: data <= 21'h1fdcc0; 
        10'b0011010010: data <= 21'h1fd3eb; 
        10'b0011010011: data <= 21'h1fd397; 
        10'b0011010100: data <= 21'h1fd254; 
        10'b0011010101: data <= 21'h1fe2e1; 
        10'b0011010110: data <= 21'h1fe22c; 
        10'b0011010111: data <= 21'h1feb3c; 
        10'b0011011000: data <= 21'h1fe7ff; 
        10'b0011011001: data <= 21'h1ff50d; 
        10'b0011011010: data <= 21'h001463; 
        10'b0011011011: data <= 21'h001b96; 
        10'b0011011100: data <= 21'h000eb8; 
        10'b0011011101: data <= 21'h00084b; 
        10'b0011011110: data <= 21'h0007c6; 
        10'b0011011111: data <= 21'h00049e; 
        10'b0011100000: data <= 21'h00077e; 
        10'b0011100001: data <= 21'h00064a; 
        10'b0011100010: data <= 21'h000846; 
        10'b0011100011: data <= 21'h00019a; 
        10'b0011100100: data <= 21'h00027e; 
        10'b0011100101: data <= 21'h000369; 
        10'b0011100110: data <= 21'h00024b; 
        10'b0011100111: data <= 21'h1ffe02; 
        10'b0011101000: data <= 21'h1fed6f; 
        10'b0011101001: data <= 21'h1ff68f; 
        10'b0011101010: data <= 21'h1ff3aa; 
        10'b0011101011: data <= 21'h1fe730; 
        10'b0011101100: data <= 21'h1fdba9; 
        10'b0011101101: data <= 21'h1fe8c5; 
        10'b0011101110: data <= 21'h1fcb57; 
        10'b0011101111: data <= 21'h1fc9e8; 
        10'b0011110000: data <= 21'h1fd5f4; 
        10'b0011110001: data <= 21'h1fe5aa; 
        10'b0011110010: data <= 21'h1fe85d; 
        10'b0011110011: data <= 21'h1ff88f; 
        10'b0011110100: data <= 21'h1ff193; 
        10'b0011110101: data <= 21'h1ff1d2; 
        10'b0011110110: data <= 21'h000965; 
        10'b0011110111: data <= 21'h000e75; 
        10'b0011111000: data <= 21'h000b07; 
        10'b0011111001: data <= 21'h000231; 
        10'b0011111010: data <= 21'h0002f9; 
        10'b0011111011: data <= 21'h000567; 
        10'b0011111100: data <= 21'h0008e8; 
        10'b0011111101: data <= 21'h00077e; 
        10'b0011111110: data <= 21'h0006ff; 
        10'b0011111111: data <= 21'h000178; 
        10'b0100000000: data <= 21'h1ffb5b; 
        10'b0100000001: data <= 21'h000023; 
        10'b0100000010: data <= 21'h1ff48c; 
        10'b0100000011: data <= 21'h1ff7c8; 
        10'b0100000100: data <= 21'h1ffaaa; 
        10'b0100000101: data <= 21'h1ffe3f; 
        10'b0100000110: data <= 21'h1ff9a5; 
        10'b0100000111: data <= 21'h1ff85b; 
        10'b0100001000: data <= 21'h1ff81f; 
        10'b0100001001: data <= 21'h1feb0b; 
        10'b0100001010: data <= 21'h1fb418; 
        10'b0100001011: data <= 21'h1fc736; 
        10'b0100001100: data <= 21'h1ff23a; 
        10'b0100001101: data <= 21'h1ff5d2; 
        10'b0100001110: data <= 21'h1ffcdb; 
        10'b0100001111: data <= 21'h0001af; 
        10'b0100010000: data <= 21'h1ff806; 
        10'b0100010001: data <= 21'h1ff835; 
        10'b0100010010: data <= 21'h0003ee; 
        10'b0100010011: data <= 21'h0000e5; 
        10'b0100010100: data <= 21'h1ff6f6; 
        10'b0100010101: data <= 21'h1ff699; 
        10'b0100010110: data <= 21'h1ffbec; 
        10'b0100010111: data <= 21'h000604; 
        10'b0100011000: data <= 21'h0004c0; 
        10'b0100011001: data <= 21'h00035d; 
        10'b0100011010: data <= 21'h000366; 
        10'b0100011011: data <= 21'h0000ee; 
        10'b0100011100: data <= 21'h000388; 
        10'b0100011101: data <= 21'h1ff5c8; 
        10'b0100011110: data <= 21'h1fef19; 
        10'b0100011111: data <= 21'h1ff7cb; 
        10'b0100100000: data <= 21'h000272; 
        10'b0100100001: data <= 21'h0015a1; 
        10'b0100100010: data <= 21'h000d18; 
        10'b0100100011: data <= 21'h0009ca; 
        10'b0100100100: data <= 21'h000bb8; 
        10'b0100100101: data <= 21'h1fe2f9; 
        10'b0100100110: data <= 21'h1fafd8; 
        10'b0100100111: data <= 21'h1fe791; 
        10'b0100101000: data <= 21'h0002cc; 
        10'b0100101001: data <= 21'h1ffc66; 
        10'b0100101010: data <= 21'h1ffd42; 
        10'b0100101011: data <= 21'h0002d6; 
        10'b0100101100: data <= 21'h1ff000; 
        10'b0100101101: data <= 21'h1ff56e; 
        10'b0100101110: data <= 21'h1ffe01; 
        10'b0100101111: data <= 21'h1fee95; 
        10'b0100110000: data <= 21'h1ff622; 
        10'b0100110001: data <= 21'h1ff9be; 
        10'b0100110010: data <= 21'h0004fd; 
        10'b0100110011: data <= 21'h00083e; 
        10'b0100110100: data <= 21'h00058c; 
        10'b0100110101: data <= 21'h0005c9; 
        10'b0100110110: data <= 21'h0004e2; 
        10'b0100110111: data <= 21'h1ffcf1; 
        10'b0100111000: data <= 21'h1ffedf; 
        10'b0100111001: data <= 21'h1ffa4a; 
        10'b0100111010: data <= 21'h1ff9f4; 
        10'b0100111011: data <= 21'h00051f; 
        10'b0100111100: data <= 21'h00105e; 
        10'b0100111101: data <= 21'h001b94; 
        10'b0100111110: data <= 21'h002603; 
        10'b0100111111: data <= 21'h00182e; 
        10'b0101000000: data <= 21'h001b4b; 
        10'b0101000001: data <= 21'h1fd389; 
        10'b0101000010: data <= 21'h1fc3a4; 
        10'b0101000011: data <= 21'h0007d6; 
        10'b0101000100: data <= 21'h001f37; 
        10'b0101000101: data <= 21'h000542; 
        10'b0101000110: data <= 21'h1ffe31; 
        10'b0101000111: data <= 21'h1ffafe; 
        10'b0101001000: data <= 21'h1feeed; 
        10'b0101001001: data <= 21'h1ff167; 
        10'b0101001010: data <= 21'h1ff88f; 
        10'b0101001011: data <= 21'h1ff27f; 
        10'b0101001100: data <= 21'h1ff0fe; 
        10'b0101001101: data <= 21'h1fff28; 
        10'b0101001110: data <= 21'h1fff7e; 
        10'b0101001111: data <= 21'h000211; 
        10'b0101010000: data <= 21'h000632; 
        10'b0101010001: data <= 21'h00056e; 
        10'b0101010010: data <= 21'h000294; 
        10'b0101010011: data <= 21'h0003b8; 
        10'b0101010100: data <= 21'h1fff9f; 
        10'b0101010101: data <= 21'h1ffa6b; 
        10'b0101010110: data <= 21'h00100e; 
        10'b0101010111: data <= 21'h001a76; 
        10'b0101011000: data <= 21'h0028fd; 
        10'b0101011001: data <= 21'h0023ea; 
        10'b0101011010: data <= 21'h003bbd; 
        10'b0101011011: data <= 21'h0043af; 
        10'b0101011100: data <= 21'h003ffa; 
        10'b0101011101: data <= 21'h1ffef0; 
        10'b0101011110: data <= 21'h1fe02d; 
        10'b0101011111: data <= 21'h00190a; 
        10'b0101100000: data <= 21'h0028a9; 
        10'b0101100001: data <= 21'h00049f; 
        10'b0101100010: data <= 21'h0001b6; 
        10'b0101100011: data <= 21'h00058e; 
        10'b0101100100: data <= 21'h1fff06; 
        10'b0101100101: data <= 21'h000133; 
        10'b0101100110: data <= 21'h1ffe2f; 
        10'b0101100111: data <= 21'h1ff709; 
        10'b0101101000: data <= 21'h1ff7fc; 
        10'b0101101001: data <= 21'h1ffdbe; 
        10'b0101101010: data <= 21'h0008d5; 
        10'b0101101011: data <= 21'h00051c; 
        10'b0101101100: data <= 21'h0000f7; 
        10'b0101101101: data <= 21'h0005d1; 
        10'b0101101110: data <= 21'h0000ce; 
        10'b0101101111: data <= 21'h000270; 
        10'b0101110000: data <= 21'h0006dd; 
        10'b0101110001: data <= 21'h00135e; 
        10'b0101110010: data <= 21'h002769; 
        10'b0101110011: data <= 21'h002dba; 
        10'b0101110100: data <= 21'h003492; 
        10'b0101110101: data <= 21'h002bec; 
        10'b0101110110: data <= 21'h003341; 
        10'b0101110111: data <= 21'h005386; 
        10'b0101111000: data <= 21'h003f51; 
        10'b0101111001: data <= 21'h0000f4; 
        10'b0101111010: data <= 21'h1ff703; 
        10'b0101111011: data <= 21'h001d56; 
        10'b0101111100: data <= 21'h001e22; 
        10'b0101111101: data <= 21'h002179; 
        10'b0101111110: data <= 21'h001715; 
        10'b0101111111: data <= 21'h000a63; 
        10'b0110000000: data <= 21'h00171e; 
        10'b0110000001: data <= 21'h001103; 
        10'b0110000010: data <= 21'h00081c; 
        10'b0110000011: data <= 21'h1ffb47; 
        10'b0110000100: data <= 21'h1ffbda; 
        10'b0110000101: data <= 21'h000078; 
        10'b0110000110: data <= 21'h000718; 
        10'b0110000111: data <= 21'h000514; 
        10'b0110001000: data <= 21'h0000e7; 
        10'b0110001001: data <= 21'h000741; 
        10'b0110001010: data <= 21'h000095; 
        10'b0110001011: data <= 21'h000888; 
        10'b0110001100: data <= 21'h001125; 
        10'b0110001101: data <= 21'h002284; 
        10'b0110001110: data <= 21'h002ffa; 
        10'b0110001111: data <= 21'h003482; 
        10'b0110010000: data <= 21'h00273a; 
        10'b0110010001: data <= 21'h00257e; 
        10'b0110010010: data <= 21'h002d2e; 
        10'b0110010011: data <= 21'h0036c1; 
        10'b0110010100: data <= 21'h0027dd; 
        10'b0110010101: data <= 21'h00034e; 
        10'b0110010110: data <= 21'h1ffa32; 
        10'b0110010111: data <= 21'h000a99; 
        10'b0110011000: data <= 21'h00218f; 
        10'b0110011001: data <= 21'h003727; 
        10'b0110011010: data <= 21'h002575; 
        10'b0110011011: data <= 21'h00226e; 
        10'b0110011100: data <= 21'h001338; 
        10'b0110011101: data <= 21'h000cec; 
        10'b0110011110: data <= 21'h000434; 
        10'b0110011111: data <= 21'h000260; 
        10'b0110100000: data <= 21'h1ffea3; 
        10'b0110100001: data <= 21'h00024d; 
        10'b0110100010: data <= 21'h000452; 
        10'b0110100011: data <= 21'h00020a; 
        10'b0110100100: data <= 21'h0005fc; 
        10'b0110100101: data <= 21'h000897; 
        10'b0110100110: data <= 21'h000584; 
        10'b0110100111: data <= 21'h00071a; 
        10'b0110101000: data <= 21'h000f80; 
        10'b0110101001: data <= 21'h001194; 
        10'b0110101010: data <= 21'h001b52; 
        10'b0110101011: data <= 21'h001929; 
        10'b0110101100: data <= 21'h00287b; 
        10'b0110101101: data <= 21'h0022c7; 
        10'b0110101110: data <= 21'h001834; 
        10'b0110101111: data <= 21'h001193; 
        10'b0110110000: data <= 21'h0014c3; 
        10'b0110110001: data <= 21'h00041a; 
        10'b0110110010: data <= 21'h0010a8; 
        10'b0110110011: data <= 21'h00174d; 
        10'b0110110100: data <= 21'h00305e; 
        10'b0110110101: data <= 21'h002af9; 
        10'b0110110110: data <= 21'h001eb8; 
        10'b0110110111: data <= 21'h001233; 
        10'b0110111000: data <= 21'h1ffb1a; 
        10'b0110111001: data <= 21'h0006c1; 
        10'b0110111010: data <= 21'h000c36; 
        10'b0110111011: data <= 21'h000149; 
        10'b0110111100: data <= 21'h1ff8a6; 
        10'b0110111101: data <= 21'h0003df; 
        10'b0110111110: data <= 21'h0000fd; 
        10'b0110111111: data <= 21'h000270; 
        10'b0111000000: data <= 21'h0002a8; 
        10'b0111000001: data <= 21'h00000d; 
        10'b0111000010: data <= 21'h000051; 
        10'b0111000011: data <= 21'h1ffef0; 
        10'b0111000100: data <= 21'h000436; 
        10'b0111000101: data <= 21'h000a60; 
        10'b0111000110: data <= 21'h0010e7; 
        10'b0111000111: data <= 21'h001d85; 
        10'b0111001000: data <= 21'h002af8; 
        10'b0111001001: data <= 21'h001e9d; 
        10'b0111001010: data <= 21'h000833; 
        10'b0111001011: data <= 21'h1ffee3; 
        10'b0111001100: data <= 21'h00086a; 
        10'b0111001101: data <= 21'h000a80; 
        10'b0111001110: data <= 21'h002770; 
        10'b0111001111: data <= 21'h003688; 
        10'b0111010000: data <= 21'h00382a; 
        10'b0111010001: data <= 21'h002ea9; 
        10'b0111010010: data <= 21'h001f95; 
        10'b0111010011: data <= 21'h0003f5; 
        10'b0111010100: data <= 21'h000d3f; 
        10'b0111010101: data <= 21'h0012d0; 
        10'b0111010110: data <= 21'h000466; 
        10'b0111010111: data <= 21'h1ffce6; 
        10'b0111011000: data <= 21'h1fff25; 
        10'b0111011001: data <= 21'h0001d5; 
        10'b0111011010: data <= 21'h000364; 
        10'b0111011011: data <= 21'h00038f; 
        10'b0111011100: data <= 21'h000328; 
        10'b0111011101: data <= 21'h000339; 
        10'b0111011110: data <= 21'h00066e; 
        10'b0111011111: data <= 21'h1fffe5; 
        10'b0111100000: data <= 21'h1ffb7d; 
        10'b0111100001: data <= 21'h1ff6b8; 
        10'b0111100010: data <= 21'h00057d; 
        10'b0111100011: data <= 21'h001769; 
        10'b0111100100: data <= 21'h002d26; 
        10'b0111100101: data <= 21'h002723; 
        10'b0111100110: data <= 21'h000e2d; 
        10'b0111100111: data <= 21'h000b28; 
        10'b0111101000: data <= 21'h001027; 
        10'b0111101001: data <= 21'h0026b9; 
        10'b0111101010: data <= 21'h003ffa; 
        10'b0111101011: data <= 21'h0032a1; 
        10'b0111101100: data <= 21'h002a5b; 
        10'b0111101101: data <= 21'h000d16; 
        10'b0111101110: data <= 21'h000206; 
        10'b0111101111: data <= 21'h1ff1d4; 
        10'b0111110000: data <= 21'h00043f; 
        10'b0111110001: data <= 21'h00018d; 
        10'b0111110010: data <= 21'h1ff756; 
        10'b0111110011: data <= 21'h1ffc45; 
        10'b0111110100: data <= 21'h1ffa5b; 
        10'b0111110101: data <= 21'h1ffcc5; 
        10'b0111110110: data <= 21'h0005b2; 
        10'b0111110111: data <= 21'h0006f7; 
        10'b0111111000: data <= 21'h00037d; 
        10'b0111111001: data <= 21'h000558; 
        10'b0111111010: data <= 21'h0004ad; 
        10'b0111111011: data <= 21'h0000b2; 
        10'b0111111100: data <= 21'h1ffa8c; 
        10'b0111111101: data <= 21'h1ff487; 
        10'b0111111110: data <= 21'h1ff2ae; 
        10'b0111111111: data <= 21'h1fffbe; 
        10'b1000000000: data <= 21'h000b8d; 
        10'b1000000001: data <= 21'h0002a4; 
        10'b1000000010: data <= 21'h1ff698; 
        10'b1000000011: data <= 21'h1ffa70; 
        10'b1000000100: data <= 21'h000ec4; 
        10'b1000000101: data <= 21'h0010a5; 
        10'b1000000110: data <= 21'h001c1e; 
        10'b1000000111: data <= 21'h00180e; 
        10'b1000001000: data <= 21'h000c91; 
        10'b1000001001: data <= 21'h1fec8b; 
        10'b1000001010: data <= 21'h1fed92; 
        10'b1000001011: data <= 21'h1fe4f8; 
        10'b1000001100: data <= 21'h1feff7; 
        10'b1000001101: data <= 21'h1fef5f; 
        10'b1000001110: data <= 21'h1fe9d9; 
        10'b1000001111: data <= 21'h1feed5; 
        10'b1000010000: data <= 21'h1ffb86; 
        10'b1000010001: data <= 21'h1ffda1; 
        10'b1000010010: data <= 21'h00020f; 
        10'b1000010011: data <= 21'h000049; 
        10'b1000010100: data <= 21'h000360; 
        10'b1000010101: data <= 21'h000640; 
        10'b1000010110: data <= 21'h000261; 
        10'b1000010111: data <= 21'h00016d; 
        10'b1000011000: data <= 21'h1ff3a0; 
        10'b1000011001: data <= 21'h1ff0a1; 
        10'b1000011010: data <= 21'h1febb0; 
        10'b1000011011: data <= 21'h1fe17c; 
        10'b1000011100: data <= 21'h1fdd95; 
        10'b1000011101: data <= 21'h1fdb52; 
        10'b1000011110: data <= 21'h1fd4b8; 
        10'b1000011111: data <= 21'h1fd69a; 
        10'b1000100000: data <= 21'h1fdb58; 
        10'b1000100001: data <= 21'h1fea84; 
        10'b1000100010: data <= 21'h1ff99e; 
        10'b1000100011: data <= 21'h000594; 
        10'b1000100100: data <= 21'h1fef55; 
        10'b1000100101: data <= 21'h1ff1a7; 
        10'b1000100110: data <= 21'h1fee54; 
        10'b1000100111: data <= 21'h1fe79e; 
        10'b1000101000: data <= 21'h1fe4be; 
        10'b1000101001: data <= 21'h1fe6e5; 
        10'b1000101010: data <= 21'h1fe67c; 
        10'b1000101011: data <= 21'h1feebf; 
        10'b1000101100: data <= 21'h1ffb73; 
        10'b1000101101: data <= 21'h00036b; 
        10'b1000101110: data <= 21'h00060b; 
        10'b1000101111: data <= 21'h000586; 
        10'b1000110000: data <= 21'h0008ff; 
        10'b1000110001: data <= 21'h000853; 
        10'b1000110010: data <= 21'h000268; 
        10'b1000110011: data <= 21'h00016e; 
        10'b1000110100: data <= 21'h1ff5f6; 
        10'b1000110101: data <= 21'h1feed3; 
        10'b1000110110: data <= 21'h1fe70b; 
        10'b1000110111: data <= 21'h1fd762; 
        10'b1000111000: data <= 21'h1fcfb9; 
        10'b1000111001: data <= 21'h1fccd8; 
        10'b1000111010: data <= 21'h1fcbe8; 
        10'b1000111011: data <= 21'h1fd9dc; 
        10'b1000111100: data <= 21'h1fe129; 
        10'b1000111101: data <= 21'h1fdd86; 
        10'b1000111110: data <= 21'h1fea56; 
        10'b1000111111: data <= 21'h1ff4b6; 
        10'b1001000000: data <= 21'h1ffc1a; 
        10'b1001000001: data <= 21'h1ffdd2; 
        10'b1001000010: data <= 21'h1ff70b; 
        10'b1001000011: data <= 21'h1fec97; 
        10'b1001000100: data <= 21'h1ff2f3; 
        10'b1001000101: data <= 21'h1ff13c; 
        10'b1001000110: data <= 21'h1fee2d; 
        10'b1001000111: data <= 21'h1ff6dc; 
        10'b1001001000: data <= 21'h1ff73a; 
        10'b1001001001: data <= 21'h0000a5; 
        10'b1001001010: data <= 21'h00021e; 
        10'b1001001011: data <= 21'h000604; 
        10'b1001001100: data <= 21'h0001a9; 
        10'b1001001101: data <= 21'h00029f; 
        10'b1001001110: data <= 21'h0000af; 
        10'b1001001111: data <= 21'h000132; 
        10'b1001010000: data <= 21'h1fffe6; 
        10'b1001010001: data <= 21'h1ff637; 
        10'b1001010010: data <= 21'h1fe769; 
        10'b1001010011: data <= 21'h1fdd8d; 
        10'b1001010100: data <= 21'h1fe0fd; 
        10'b1001010101: data <= 21'h1fdcbd; 
        10'b1001010110: data <= 21'h1fe14d; 
        10'b1001010111: data <= 21'h1fe934; 
        10'b1001011000: data <= 21'h1fed0a; 
        10'b1001011001: data <= 21'h1fee70; 
        10'b1001011010: data <= 21'h1febe2; 
        10'b1001011011: data <= 21'h1ff6b2; 
        10'b1001011100: data <= 21'h1ff397; 
        10'b1001011101: data <= 21'h00023c; 
        10'b1001011110: data <= 21'h1ffc4c; 
        10'b1001011111: data <= 21'h0000ac; 
        10'b1001100000: data <= 21'h1ffe63; 
        10'b1001100001: data <= 21'h1ff3ed; 
        10'b1001100010: data <= 21'h1ff5c5; 
        10'b1001100011: data <= 21'h1ffe1d; 
        10'b1001100100: data <= 21'h1fffac; 
        10'b1001100101: data <= 21'h0003b9; 
        10'b1001100110: data <= 21'h0004ff; 
        10'b1001100111: data <= 21'h0004d1; 
        10'b1001101000: data <= 21'h000455; 
        10'b1001101001: data <= 21'h000509; 
        10'b1001101010: data <= 21'h000201; 
        10'b1001101011: data <= 21'h000584; 
        10'b1001101100: data <= 21'h1ffeb3; 
        10'b1001101101: data <= 21'h1ffac8; 
        10'b1001101110: data <= 21'h1ff5da; 
        10'b1001101111: data <= 21'h1fef3f; 
        10'b1001110000: data <= 21'h1fe95d; 
        10'b1001110001: data <= 21'h1ff241; 
        10'b1001110010: data <= 21'h1ff1d5; 
        10'b1001110011: data <= 21'h1ff62c; 
        10'b1001110100: data <= 21'h1ff5a3; 
        10'b1001110101: data <= 21'h1ff71b; 
        10'b1001110110: data <= 21'h1ff4e4; 
        10'b1001110111: data <= 21'h1ff92c; 
        10'b1001111000: data <= 21'h1ff973; 
        10'b1001111001: data <= 21'h00025c; 
        10'b1001111010: data <= 21'h000a0a; 
        10'b1001111011: data <= 21'h001061; 
        10'b1001111100: data <= 21'h000c92; 
        10'b1001111101: data <= 21'h00083e; 
        10'b1001111110: data <= 21'h1ffa8c; 
        10'b1001111111: data <= 21'h1ffaa4; 
        10'b1010000000: data <= 21'h1fffcc; 
        10'b1010000001: data <= 21'h000398; 
        10'b1010000010: data <= 21'h000093; 
        10'b1010000011: data <= 21'h0002c2; 
        10'b1010000100: data <= 21'h0002cf; 
        10'b1010000101: data <= 21'h000031; 
        10'b1010000110: data <= 21'h00027c; 
        10'b1010000111: data <= 21'h0004e9; 
        10'b1010001000: data <= 21'h0002c6; 
        10'b1010001001: data <= 21'h000368; 
        10'b1010001010: data <= 21'h1ffa99; 
        10'b1010001011: data <= 21'h1ff9fd; 
        10'b1010001100: data <= 21'h1ff7de; 
        10'b1010001101: data <= 21'h0003ca; 
        10'b1010001110: data <= 21'h1ff740; 
        10'b1010001111: data <= 21'h00016a; 
        10'b1010010000: data <= 21'h1ff6f4; 
        10'b1010010001: data <= 21'h1ff8e4; 
        10'b1010010010: data <= 21'h1ff90e; 
        10'b1010010011: data <= 21'h1fff7d; 
        10'b1010010100: data <= 21'h000250; 
        10'b1010010101: data <= 21'h00061d; 
        10'b1010010110: data <= 21'h0012d8; 
        10'b1010010111: data <= 21'h001263; 
        10'b1010011000: data <= 21'h000fac; 
        10'b1010011001: data <= 21'h0006fb; 
        10'b1010011010: data <= 21'h1ffd69; 
        10'b1010011011: data <= 21'h00021f; 
        10'b1010011100: data <= 21'h000428; 
        10'b1010011101: data <= 21'h0005b0; 
        10'b1010011110: data <= 21'h0001db; 
        10'b1010011111: data <= 21'h000715; 
        10'b1010100000: data <= 21'h00055a; 
        10'b1010100001: data <= 21'h0007a6; 
        10'b1010100010: data <= 21'h00039f; 
        10'b1010100011: data <= 21'h000610; 
        10'b1010100100: data <= 21'h00016d; 
        10'b1010100101: data <= 21'h0004a4; 
        10'b1010100110: data <= 21'h0001c4; 
        10'b1010100111: data <= 21'h1ff763; 
        10'b1010101000: data <= 21'h1ff734; 
        10'b1010101001: data <= 21'h1ffd33; 
        10'b1010101010: data <= 21'h1ff6ac; 
        10'b1010101011: data <= 21'h1ffe7a; 
        10'b1010101100: data <= 21'h1ff94b; 
        10'b1010101101: data <= 21'h1ff9d2; 
        10'b1010101110: data <= 21'h1ff4a0; 
        10'b1010101111: data <= 21'h1ff33d; 
        10'b1010110000: data <= 21'h1ffa7e; 
        10'b1010110001: data <= 21'h1ffd24; 
        10'b1010110010: data <= 21'h000100; 
        10'b1010110011: data <= 21'h0009e8; 
        10'b1010110100: data <= 21'h00073c; 
        10'b1010110101: data <= 21'h1ffd0a; 
        10'b1010110110: data <= 21'h1fff26; 
        10'b1010110111: data <= 21'h0003d3; 
        10'b1010111000: data <= 21'h00064c; 
        10'b1010111001: data <= 21'h000101; 
        10'b1010111010: data <= 21'h0001a2; 
        10'b1010111011: data <= 21'h000574; 
        10'b1010111100: data <= 21'h000802; 
        10'b1010111101: data <= 21'h0007c4; 
        10'b1010111110: data <= 21'h000718; 
        10'b1010111111: data <= 21'h000197; 
        10'b1011000000: data <= 21'h000723; 
        10'b1011000001: data <= 21'h000057; 
        10'b1011000010: data <= 21'h1ffae6; 
        10'b1011000011: data <= 21'h1ff7b2; 
        10'b1011000100: data <= 21'h1ff381; 
        10'b1011000101: data <= 21'h1ff2db; 
        10'b1011000110: data <= 21'h1fea6b; 
        10'b1011000111: data <= 21'h1fe7a8; 
        10'b1011001000: data <= 21'h1fe903; 
        10'b1011001001: data <= 21'h1fe922; 
        10'b1011001010: data <= 21'h1fec91; 
        10'b1011001011: data <= 21'h1feb6e; 
        10'b1011001100: data <= 21'h1fe562; 
        10'b1011001101: data <= 21'h1fe1a9; 
        10'b1011001110: data <= 21'h1fe4c2; 
        10'b1011001111: data <= 21'h1ff111; 
        10'b1011010000: data <= 21'h1ff258; 
        10'b1011010001: data <= 21'h1ffb12; 
        10'b1011010010: data <= 21'h00004e; 
        10'b1011010011: data <= 21'h000539; 
        10'b1011010100: data <= 21'h000064; 
        10'b1011010101: data <= 21'h000742; 
        10'b1011010110: data <= 21'h0002e7; 
        10'b1011010111: data <= 21'h0002a3; 
        10'b1011011000: data <= 21'h0003bf; 
        10'b1011011001: data <= 21'h000566; 
        10'b1011011010: data <= 21'h000138; 
        10'b1011011011: data <= 21'h000399; 
        10'b1011011100: data <= 21'h1fffa3; 
        10'b1011011101: data <= 21'h1ffec3; 
        10'b1011011110: data <= 21'h00022b; 
        10'b1011011111: data <= 21'h000190; 
        10'b1011100000: data <= 21'h1ffe5b; 
        10'b1011100001: data <= 21'h1ff871; 
        10'b1011100010: data <= 21'h1fedc7; 
        10'b1011100011: data <= 21'h1ff01a; 
        10'b1011100100: data <= 21'h1fedd0; 
        10'b1011100101: data <= 21'h1fe74c; 
        10'b1011100110: data <= 21'h1fe503; 
        10'b1011100111: data <= 21'h1feafe; 
        10'b1011101000: data <= 21'h1fe813; 
        10'b1011101001: data <= 21'h1febaf; 
        10'b1011101010: data <= 21'h1fef53; 
        10'b1011101011: data <= 21'h1ff610; 
        10'b1011101100: data <= 21'h1ffc5d; 
        10'b1011101101: data <= 21'h000562; 
        10'b1011101110: data <= 21'h000555; 
        10'b1011101111: data <= 21'h0000ad; 
        10'b1011110000: data <= 21'h000380; 
        10'b1011110001: data <= 21'h000093; 
        10'b1011110010: data <= 21'h000896; 
        10'b1011110011: data <= 21'h0003c2; 
        10'b1011110100: data <= 21'h000535; 
        10'b1011110101: data <= 21'h0000c4; 
        10'b1011110110: data <= 21'h000128; 
        10'b1011110111: data <= 21'h000841; 
        10'b1011111000: data <= 21'h000318; 
        10'b1011111001: data <= 21'h0006df; 
        10'b1011111010: data <= 21'h00032b; 
        10'b1011111011: data <= 21'h00086a; 
        10'b1011111100: data <= 21'h1ffffc; 
        10'b1011111101: data <= 21'h0003a1; 
        10'b1011111110: data <= 21'h0001dc; 
        10'b1011111111: data <= 21'h1ffed4; 
        10'b1100000000: data <= 21'h1fff24; 
        10'b1100000001: data <= 21'h00004f; 
        10'b1100000010: data <= 21'h1ffc80; 
        10'b1100000011: data <= 21'h0006ad; 
        10'b1100000100: data <= 21'h1ffe4a; 
        10'b1100000101: data <= 21'h1ffe0b; 
        10'b1100000110: data <= 21'h1fff56; 
        10'b1100000111: data <= 21'h000384; 
        10'b1100001000: data <= 21'h0002b3; 
        10'b1100001001: data <= 21'h0002af; 
        10'b1100001010: data <= 21'h0002da; 
        10'b1100001011: data <= 21'h0004df; 
        10'b1100001100: data <= 21'h0004a9; 
        10'b1100001101: data <= 21'h000629; 
        10'b1100001110: data <= 21'h00046a; 
        10'b1100001111: data <= 21'h0002ee; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 16) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 22'h3ffffd; 
        10'b0000000001: data <= 22'h000240; 
        10'b0000000010: data <= 22'h000f1f; 
        10'b0000000011: data <= 22'h000f1a; 
        10'b0000000100: data <= 22'h000047; 
        10'b0000000101: data <= 22'h000049; 
        10'b0000000110: data <= 22'h000bd7; 
        10'b0000000111: data <= 22'h00033c; 
        10'b0000001000: data <= 22'h000100; 
        10'b0000001001: data <= 22'h00023c; 
        10'b0000001010: data <= 22'h000070; 
        10'b0000001011: data <= 22'h000adf; 
        10'b0000001100: data <= 22'h000e4e; 
        10'b0000001101: data <= 22'h000825; 
        10'b0000001110: data <= 22'h000a84; 
        10'b0000001111: data <= 22'h00012a; 
        10'b0000010000: data <= 22'h0009d9; 
        10'b0000010001: data <= 22'h000d81; 
        10'b0000010010: data <= 22'h0002d8; 
        10'b0000010011: data <= 22'h000ae6; 
        10'b0000010100: data <= 22'h0000d0; 
        10'b0000010101: data <= 22'h000679; 
        10'b0000010110: data <= 22'h000e90; 
        10'b0000010111: data <= 22'h000174; 
        10'b0000011000: data <= 22'h000e8e; 
        10'b0000011001: data <= 22'h00024f; 
        10'b0000011010: data <= 22'h000feb; 
        10'b0000011011: data <= 22'h00068e; 
        10'b0000011100: data <= 22'h00042a; 
        10'b0000011101: data <= 22'h000773; 
        10'b0000011110: data <= 22'h3fffe1; 
        10'b0000011111: data <= 22'h000140; 
        10'b0000100000: data <= 22'h000748; 
        10'b0000100001: data <= 22'h001190; 
        10'b0000100010: data <= 22'h0003a2; 
        10'b0000100011: data <= 22'h3ffd2f; 
        10'b0000100100: data <= 22'h0009c1; 
        10'b0000100101: data <= 22'h00005a; 
        10'b0000100110: data <= 22'h00068b; 
        10'b0000100111: data <= 22'h3ffae2; 
        10'b0000101000: data <= 22'h000481; 
        10'b0000101001: data <= 22'h3ff8f5; 
        10'b0000101010: data <= 22'h000060; 
        10'b0000101011: data <= 22'h0009a6; 
        10'b0000101100: data <= 22'h000b5f; 
        10'b0000101101: data <= 22'h000358; 
        10'b0000101110: data <= 22'h00002d; 
        10'b0000101111: data <= 22'h0002db; 
        10'b0000110000: data <= 22'h000c3b; 
        10'b0000110001: data <= 22'h3fffb6; 
        10'b0000110010: data <= 22'h3fff98; 
        10'b0000110011: data <= 22'h000101; 
        10'b0000110100: data <= 22'h000ad4; 
        10'b0000110101: data <= 22'h000b77; 
        10'b0000110110: data <= 22'h0002b7; 
        10'b0000110111: data <= 22'h000b6e; 
        10'b0000111000: data <= 22'h000d1c; 
        10'b0000111001: data <= 22'h000886; 
        10'b0000111010: data <= 22'h000cf0; 
        10'b0000111011: data <= 22'h000d45; 
        10'b0000111100: data <= 22'h000c92; 
        10'b0000111101: data <= 22'h000b35; 
        10'b0000111110: data <= 22'h000ee4; 
        10'b0000111111: data <= 22'h3ffb3d; 
        10'b0001000000: data <= 22'h3ffade; 
        10'b0001000001: data <= 22'h0002b6; 
        10'b0001000010: data <= 22'h3ffe40; 
        10'b0001000011: data <= 22'h3ff72b; 
        10'b0001000100: data <= 22'h3fddd8; 
        10'b0001000101: data <= 22'h3ff234; 
        10'b0001000110: data <= 22'h3fef78; 
        10'b0001000111: data <= 22'h3fe899; 
        10'b0001001000: data <= 22'h3feef5; 
        10'b0001001001: data <= 22'h3ffca6; 
        10'b0001001010: data <= 22'h000444; 
        10'b0001001011: data <= 22'h000c04; 
        10'b0001001100: data <= 22'h000f9b; 
        10'b0001001101: data <= 22'h0008ff; 
        10'b0001001110: data <= 22'h000eb4; 
        10'b0001001111: data <= 22'h0003f6; 
        10'b0001010000: data <= 22'h000592; 
        10'b0001010001: data <= 22'h0009f2; 
        10'b0001010010: data <= 22'h00009e; 
        10'b0001010011: data <= 22'h0006ed; 
        10'b0001010100: data <= 22'h000d39; 
        10'b0001010101: data <= 22'h000be3; 
        10'b0001010110: data <= 22'h000497; 
        10'b0001010111: data <= 22'h00077b; 
        10'b0001011000: data <= 22'h0007c1; 
        10'b0001011001: data <= 22'h00001b; 
        10'b0001011010: data <= 22'h0009ed; 
        10'b0001011011: data <= 22'h3ff734; 
        10'b0001011100: data <= 22'h3ff326; 
        10'b0001011101: data <= 22'h3ff8fe; 
        10'b0001011110: data <= 22'h3fe2a3; 
        10'b0001011111: data <= 22'h3fdd40; 
        10'b0001100000: data <= 22'h3fc88f; 
        10'b0001100001: data <= 22'h3fcb1b; 
        10'b0001100010: data <= 22'h3fcda1; 
        10'b0001100011: data <= 22'h3fc2e0; 
        10'b0001100100: data <= 22'h3fd731; 
        10'b0001100101: data <= 22'h3feb9e; 
        10'b0001100110: data <= 22'h0002ff; 
        10'b0001100111: data <= 22'h000689; 
        10'b0001101000: data <= 22'h000bd6; 
        10'b0001101001: data <= 22'h001171; 
        10'b0001101010: data <= 22'h000491; 
        10'b0001101011: data <= 22'h0004a8; 
        10'b0001101100: data <= 22'h0010f8; 
        10'b0001101101: data <= 22'h00104d; 
        10'b0001101110: data <= 22'h00050b; 
        10'b0001101111: data <= 22'h000991; 
        10'b0001110000: data <= 22'h00107c; 
        10'b0001110001: data <= 22'h000af0; 
        10'b0001110010: data <= 22'h000c52; 
        10'b0001110011: data <= 22'h000bf3; 
        10'b0001110100: data <= 22'h00071c; 
        10'b0001110101: data <= 22'h000d81; 
        10'b0001110110: data <= 22'h3ff5df; 
        10'b0001110111: data <= 22'h3ffdbe; 
        10'b0001111000: data <= 22'h3feb54; 
        10'b0001111001: data <= 22'h3fee84; 
        10'b0001111010: data <= 22'h3fce4a; 
        10'b0001111011: data <= 22'h3fd0b4; 
        10'b0001111100: data <= 22'h3fbf52; 
        10'b0001111101: data <= 22'h3fca49; 
        10'b0001111110: data <= 22'h3fbe0d; 
        10'b0001111111: data <= 22'h3fc78b; 
        10'b0010000000: data <= 22'h3fe492; 
        10'b0010000001: data <= 22'h3fe79e; 
        10'b0010000010: data <= 22'h3ff169; 
        10'b0010000011: data <= 22'h000e07; 
        10'b0010000100: data <= 22'h001353; 
        10'b0010000101: data <= 22'h001613; 
        10'b0010000110: data <= 22'h001505; 
        10'b0010000111: data <= 22'h001be1; 
        10'b0010001000: data <= 22'h0007ba; 
        10'b0010001001: data <= 22'h000faa; 
        10'b0010001010: data <= 22'h0003fc; 
        10'b0010001011: data <= 22'h000292; 
        10'b0010001100: data <= 22'h0010c5; 
        10'b0010001101: data <= 22'h0004b2; 
        10'b0010001110: data <= 22'h000bd7; 
        10'b0010001111: data <= 22'h0003e0; 
        10'b0010010000: data <= 22'h000ada; 
        10'b0010010001: data <= 22'h000230; 
        10'b0010010010: data <= 22'h0007ad; 
        10'b0010010011: data <= 22'h3ff6af; 
        10'b0010010100: data <= 22'h000280; 
        10'b0010010101: data <= 22'h3ff53b; 
        10'b0010010110: data <= 22'h3fdba3; 
        10'b0010010111: data <= 22'h3fe7eb; 
        10'b0010011000: data <= 22'h3fd6b0; 
        10'b0010011001: data <= 22'h3fccba; 
        10'b0010011010: data <= 22'h3fdc23; 
        10'b0010011011: data <= 22'h3fe267; 
        10'b0010011100: data <= 22'h3ffb0b; 
        10'b0010011101: data <= 22'h00048b; 
        10'b0010011110: data <= 22'h3ff8e8; 
        10'b0010011111: data <= 22'h000bf1; 
        10'b0010100000: data <= 22'h000ea6; 
        10'b0010100001: data <= 22'h0013ca; 
        10'b0010100010: data <= 22'h002e1e; 
        10'b0010100011: data <= 22'h003409; 
        10'b0010100100: data <= 22'h001c4e; 
        10'b0010100101: data <= 22'h3ffd3a; 
        10'b0010100110: data <= 22'h0004a6; 
        10'b0010100111: data <= 22'h0002cf; 
        10'b0010101000: data <= 22'h000f90; 
        10'b0010101001: data <= 22'h001136; 
        10'b0010101010: data <= 22'h000520; 
        10'b0010101011: data <= 22'h000d88; 
        10'b0010101100: data <= 22'h000eba; 
        10'b0010101101: data <= 22'h000c19; 
        10'b0010101110: data <= 22'h000bfe; 
        10'b0010101111: data <= 22'h3fff0d; 
        10'b0010110000: data <= 22'h3ffd49; 
        10'b0010110001: data <= 22'h3ff1b9; 
        10'b0010110010: data <= 22'h3fe328; 
        10'b0010110011: data <= 22'h3fcd41; 
        10'b0010110100: data <= 22'h3fb31c; 
        10'b0010110101: data <= 22'h3fa519; 
        10'b0010110110: data <= 22'h3fa112; 
        10'b0010110111: data <= 22'h3fad98; 
        10'b0010111000: data <= 22'h3fab90; 
        10'b0010111001: data <= 22'h3fce81; 
        10'b0010111010: data <= 22'h3fccd8; 
        10'b0010111011: data <= 22'h3fe8fd; 
        10'b0010111100: data <= 22'h3ff0dc; 
        10'b0010111101: data <= 22'h3ffed8; 
        10'b0010111110: data <= 22'h004203; 
        10'b0010111111: data <= 22'h004559; 
        10'b0011000000: data <= 22'h001aae; 
        10'b0011000001: data <= 22'h0014eb; 
        10'b0011000010: data <= 22'h000ef3; 
        10'b0011000011: data <= 22'h0000a4; 
        10'b0011000100: data <= 22'h00075b; 
        10'b0011000101: data <= 22'h0003da; 
        10'b0011000110: data <= 22'h00054c; 
        10'b0011000111: data <= 22'h00095e; 
        10'b0011001000: data <= 22'h00055f; 
        10'b0011001001: data <= 22'h000c88; 
        10'b0011001010: data <= 22'h3ff83f; 
        10'b0011001011: data <= 22'h3ffe96; 
        10'b0011001100: data <= 22'h3ff76a; 
        10'b0011001101: data <= 22'h3fec84; 
        10'b0011001110: data <= 22'h3fcec0; 
        10'b0011001111: data <= 22'h3fb333; 
        10'b0011010000: data <= 22'h3f9c3d; 
        10'b0011010001: data <= 22'h3fb97f; 
        10'b0011010010: data <= 22'h3fa7d6; 
        10'b0011010011: data <= 22'h3fa72e; 
        10'b0011010100: data <= 22'h3fa4a7; 
        10'b0011010101: data <= 22'h3fc5c3; 
        10'b0011010110: data <= 22'h3fc457; 
        10'b0011010111: data <= 22'h3fd677; 
        10'b0011011000: data <= 22'h3fcffe; 
        10'b0011011001: data <= 22'h3fea19; 
        10'b0011011010: data <= 22'h0028c6; 
        10'b0011011011: data <= 22'h00372c; 
        10'b0011011100: data <= 22'h001d6f; 
        10'b0011011101: data <= 22'h001095; 
        10'b0011011110: data <= 22'h000f8b; 
        10'b0011011111: data <= 22'h00093b; 
        10'b0011100000: data <= 22'h000efb; 
        10'b0011100001: data <= 22'h000c93; 
        10'b0011100010: data <= 22'h00108c; 
        10'b0011100011: data <= 22'h000333; 
        10'b0011100100: data <= 22'h0004fb; 
        10'b0011100101: data <= 22'h0006d2; 
        10'b0011100110: data <= 22'h000496; 
        10'b0011100111: data <= 22'h3ffc04; 
        10'b0011101000: data <= 22'h3fdadf; 
        10'b0011101001: data <= 22'h3fed1d; 
        10'b0011101010: data <= 22'h3fe754; 
        10'b0011101011: data <= 22'h3fce60; 
        10'b0011101100: data <= 22'h3fb752; 
        10'b0011101101: data <= 22'h3fd18a; 
        10'b0011101110: data <= 22'h3f96ae; 
        10'b0011101111: data <= 22'h3f93d0; 
        10'b0011110000: data <= 22'h3fabe7; 
        10'b0011110001: data <= 22'h3fcb55; 
        10'b0011110010: data <= 22'h3fd0ba; 
        10'b0011110011: data <= 22'h3ff11e; 
        10'b0011110100: data <= 22'h3fe327; 
        10'b0011110101: data <= 22'h3fe3a4; 
        10'b0011110110: data <= 22'h0012c9; 
        10'b0011110111: data <= 22'h001ce9; 
        10'b0011111000: data <= 22'h00160d; 
        10'b0011111001: data <= 22'h000462; 
        10'b0011111010: data <= 22'h0005f2; 
        10'b0011111011: data <= 22'h000ace; 
        10'b0011111100: data <= 22'h0011cf; 
        10'b0011111101: data <= 22'h000efb; 
        10'b0011111110: data <= 22'h000dfd; 
        10'b0011111111: data <= 22'h0002ef; 
        10'b0100000000: data <= 22'h3ff6b7; 
        10'b0100000001: data <= 22'h000046; 
        10'b0100000010: data <= 22'h3fe918; 
        10'b0100000011: data <= 22'h3fef90; 
        10'b0100000100: data <= 22'h3ff555; 
        10'b0100000101: data <= 22'h3ffc7e; 
        10'b0100000110: data <= 22'h3ff34a; 
        10'b0100000111: data <= 22'h3ff0b6; 
        10'b0100001000: data <= 22'h3ff03e; 
        10'b0100001001: data <= 22'h3fd616; 
        10'b0100001010: data <= 22'h3f6831; 
        10'b0100001011: data <= 22'h3f8e6d; 
        10'b0100001100: data <= 22'h3fe473; 
        10'b0100001101: data <= 22'h3feba3; 
        10'b0100001110: data <= 22'h3ff9b6; 
        10'b0100001111: data <= 22'h00035d; 
        10'b0100010000: data <= 22'h3ff00c; 
        10'b0100010001: data <= 22'h3ff06a; 
        10'b0100010010: data <= 22'h0007dc; 
        10'b0100010011: data <= 22'h0001c9; 
        10'b0100010100: data <= 22'h3feded; 
        10'b0100010101: data <= 22'h3fed31; 
        10'b0100010110: data <= 22'h3ff7d9; 
        10'b0100010111: data <= 22'h000c09; 
        10'b0100011000: data <= 22'h000981; 
        10'b0100011001: data <= 22'h0006b9; 
        10'b0100011010: data <= 22'h0006cc; 
        10'b0100011011: data <= 22'h0001dd; 
        10'b0100011100: data <= 22'h000710; 
        10'b0100011101: data <= 22'h3feb90; 
        10'b0100011110: data <= 22'h3fde32; 
        10'b0100011111: data <= 22'h3fef95; 
        10'b0100100000: data <= 22'h0004e3; 
        10'b0100100001: data <= 22'h002b43; 
        10'b0100100010: data <= 22'h001a2f; 
        10'b0100100011: data <= 22'h001393; 
        10'b0100100100: data <= 22'h001770; 
        10'b0100100101: data <= 22'h3fc5f1; 
        10'b0100100110: data <= 22'h3f5fb1; 
        10'b0100100111: data <= 22'h3fcf23; 
        10'b0100101000: data <= 22'h000598; 
        10'b0100101001: data <= 22'h3ff8cd; 
        10'b0100101010: data <= 22'h3ffa84; 
        10'b0100101011: data <= 22'h0005ac; 
        10'b0100101100: data <= 22'h3fe000; 
        10'b0100101101: data <= 22'h3feadd; 
        10'b0100101110: data <= 22'h3ffc03; 
        10'b0100101111: data <= 22'h3fdd2b; 
        10'b0100110000: data <= 22'h3fec43; 
        10'b0100110001: data <= 22'h3ff37b; 
        10'b0100110010: data <= 22'h0009fb; 
        10'b0100110011: data <= 22'h00107c; 
        10'b0100110100: data <= 22'h000b18; 
        10'b0100110101: data <= 22'h000b91; 
        10'b0100110110: data <= 22'h0009c4; 
        10'b0100110111: data <= 22'h3ff9e2; 
        10'b0100111000: data <= 22'h3ffdbd; 
        10'b0100111001: data <= 22'h3ff494; 
        10'b0100111010: data <= 22'h3ff3e8; 
        10'b0100111011: data <= 22'h000a3e; 
        10'b0100111100: data <= 22'h0020bc; 
        10'b0100111101: data <= 22'h003727; 
        10'b0100111110: data <= 22'h004c06; 
        10'b0100111111: data <= 22'h00305b; 
        10'b0101000000: data <= 22'h003695; 
        10'b0101000001: data <= 22'h3fa712; 
        10'b0101000010: data <= 22'h3f8747; 
        10'b0101000011: data <= 22'h000fac; 
        10'b0101000100: data <= 22'h003e6d; 
        10'b0101000101: data <= 22'h000a84; 
        10'b0101000110: data <= 22'h3ffc63; 
        10'b0101000111: data <= 22'h3ff5fd; 
        10'b0101001000: data <= 22'h3fddda; 
        10'b0101001001: data <= 22'h3fe2cf; 
        10'b0101001010: data <= 22'h3ff11d; 
        10'b0101001011: data <= 22'h3fe4fe; 
        10'b0101001100: data <= 22'h3fe1fd; 
        10'b0101001101: data <= 22'h3ffe4f; 
        10'b0101001110: data <= 22'h3ffefc; 
        10'b0101001111: data <= 22'h000423; 
        10'b0101010000: data <= 22'h000c65; 
        10'b0101010001: data <= 22'h000add; 
        10'b0101010010: data <= 22'h000527; 
        10'b0101010011: data <= 22'h000771; 
        10'b0101010100: data <= 22'h3fff3e; 
        10'b0101010101: data <= 22'h3ff4d6; 
        10'b0101010110: data <= 22'h00201c; 
        10'b0101010111: data <= 22'h0034ed; 
        10'b0101011000: data <= 22'h0051fa; 
        10'b0101011001: data <= 22'h0047d4; 
        10'b0101011010: data <= 22'h007779; 
        10'b0101011011: data <= 22'h00875e; 
        10'b0101011100: data <= 22'h007ff4; 
        10'b0101011101: data <= 22'h3ffde1; 
        10'b0101011110: data <= 22'h3fc059; 
        10'b0101011111: data <= 22'h003213; 
        10'b0101100000: data <= 22'h005152; 
        10'b0101100001: data <= 22'h00093d; 
        10'b0101100010: data <= 22'h00036c; 
        10'b0101100011: data <= 22'h000b1b; 
        10'b0101100100: data <= 22'h3ffe0b; 
        10'b0101100101: data <= 22'h000266; 
        10'b0101100110: data <= 22'h3ffc5f; 
        10'b0101100111: data <= 22'h3fee12; 
        10'b0101101000: data <= 22'h3feff9; 
        10'b0101101001: data <= 22'h3ffb7d; 
        10'b0101101010: data <= 22'h0011ab; 
        10'b0101101011: data <= 22'h000a38; 
        10'b0101101100: data <= 22'h0001ee; 
        10'b0101101101: data <= 22'h000ba2; 
        10'b0101101110: data <= 22'h00019c; 
        10'b0101101111: data <= 22'h0004df; 
        10'b0101110000: data <= 22'h000dbb; 
        10'b0101110001: data <= 22'h0026bb; 
        10'b0101110010: data <= 22'h004ed2; 
        10'b0101110011: data <= 22'h005b73; 
        10'b0101110100: data <= 22'h006923; 
        10'b0101110101: data <= 22'h0057d7; 
        10'b0101110110: data <= 22'h006682; 
        10'b0101110111: data <= 22'h00a70d; 
        10'b0101111000: data <= 22'h007ea2; 
        10'b0101111001: data <= 22'h0001e7; 
        10'b0101111010: data <= 22'h3fee06; 
        10'b0101111011: data <= 22'h003aad; 
        10'b0101111100: data <= 22'h003c45; 
        10'b0101111101: data <= 22'h0042f1; 
        10'b0101111110: data <= 22'h002e2a; 
        10'b0101111111: data <= 22'h0014c5; 
        10'b0110000000: data <= 22'h002e3b; 
        10'b0110000001: data <= 22'h002207; 
        10'b0110000010: data <= 22'h001037; 
        10'b0110000011: data <= 22'h3ff68e; 
        10'b0110000100: data <= 22'h3ff7b4; 
        10'b0110000101: data <= 22'h0000ef; 
        10'b0110000110: data <= 22'h000e30; 
        10'b0110000111: data <= 22'h000a28; 
        10'b0110001000: data <= 22'h0001ce; 
        10'b0110001001: data <= 22'h000e81; 
        10'b0110001010: data <= 22'h000129; 
        10'b0110001011: data <= 22'h001110; 
        10'b0110001100: data <= 22'h00224a; 
        10'b0110001101: data <= 22'h004507; 
        10'b0110001110: data <= 22'h005ff4; 
        10'b0110001111: data <= 22'h006904; 
        10'b0110010000: data <= 22'h004e74; 
        10'b0110010001: data <= 22'h004afd; 
        10'b0110010010: data <= 22'h005a5b; 
        10'b0110010011: data <= 22'h006d82; 
        10'b0110010100: data <= 22'h004fba; 
        10'b0110010101: data <= 22'h00069b; 
        10'b0110010110: data <= 22'h3ff464; 
        10'b0110010111: data <= 22'h001532; 
        10'b0110011000: data <= 22'h00431f; 
        10'b0110011001: data <= 22'h006e4d; 
        10'b0110011010: data <= 22'h004aea; 
        10'b0110011011: data <= 22'h0044dc; 
        10'b0110011100: data <= 22'h002670; 
        10'b0110011101: data <= 22'h0019d8; 
        10'b0110011110: data <= 22'h000868; 
        10'b0110011111: data <= 22'h0004c0; 
        10'b0110100000: data <= 22'h3ffd46; 
        10'b0110100001: data <= 22'h00049a; 
        10'b0110100010: data <= 22'h0008a3; 
        10'b0110100011: data <= 22'h000413; 
        10'b0110100100: data <= 22'h000bf8; 
        10'b0110100101: data <= 22'h00112e; 
        10'b0110100110: data <= 22'h000b08; 
        10'b0110100111: data <= 22'h000e33; 
        10'b0110101000: data <= 22'h001f00; 
        10'b0110101001: data <= 22'h002327; 
        10'b0110101010: data <= 22'h0036a4; 
        10'b0110101011: data <= 22'h003251; 
        10'b0110101100: data <= 22'h0050f7; 
        10'b0110101101: data <= 22'h00458e; 
        10'b0110101110: data <= 22'h003068; 
        10'b0110101111: data <= 22'h002326; 
        10'b0110110000: data <= 22'h002986; 
        10'b0110110001: data <= 22'h000833; 
        10'b0110110010: data <= 22'h002150; 
        10'b0110110011: data <= 22'h002e99; 
        10'b0110110100: data <= 22'h0060bc; 
        10'b0110110101: data <= 22'h0055f3; 
        10'b0110110110: data <= 22'h003d70; 
        10'b0110110111: data <= 22'h002465; 
        10'b0110111000: data <= 22'h3ff634; 
        10'b0110111001: data <= 22'h000d82; 
        10'b0110111010: data <= 22'h00186c; 
        10'b0110111011: data <= 22'h000292; 
        10'b0110111100: data <= 22'h3ff14c; 
        10'b0110111101: data <= 22'h0007bd; 
        10'b0110111110: data <= 22'h0001fa; 
        10'b0110111111: data <= 22'h0004e0; 
        10'b0111000000: data <= 22'h000550; 
        10'b0111000001: data <= 22'h00001a; 
        10'b0111000010: data <= 22'h0000a1; 
        10'b0111000011: data <= 22'h3ffde0; 
        10'b0111000100: data <= 22'h00086c; 
        10'b0111000101: data <= 22'h0014c0; 
        10'b0111000110: data <= 22'h0021cf; 
        10'b0111000111: data <= 22'h003b0a; 
        10'b0111001000: data <= 22'h0055f0; 
        10'b0111001001: data <= 22'h003d3a; 
        10'b0111001010: data <= 22'h001066; 
        10'b0111001011: data <= 22'h3ffdc5; 
        10'b0111001100: data <= 22'h0010d5; 
        10'b0111001101: data <= 22'h0014ff; 
        10'b0111001110: data <= 22'h004edf; 
        10'b0111001111: data <= 22'h006d11; 
        10'b0111010000: data <= 22'h007054; 
        10'b0111010001: data <= 22'h005d52; 
        10'b0111010010: data <= 22'h003f2a; 
        10'b0111010011: data <= 22'h0007ea; 
        10'b0111010100: data <= 22'h001a7f; 
        10'b0111010101: data <= 22'h0025a1; 
        10'b0111010110: data <= 22'h0008cb; 
        10'b0111010111: data <= 22'h3ff9cc; 
        10'b0111011000: data <= 22'h3ffe4b; 
        10'b0111011001: data <= 22'h0003aa; 
        10'b0111011010: data <= 22'h0006c8; 
        10'b0111011011: data <= 22'h00071f; 
        10'b0111011100: data <= 22'h000650; 
        10'b0111011101: data <= 22'h000672; 
        10'b0111011110: data <= 22'h000cdc; 
        10'b0111011111: data <= 22'h3fffcb; 
        10'b0111100000: data <= 22'h3ff6fa; 
        10'b0111100001: data <= 22'h3fed71; 
        10'b0111100010: data <= 22'h000afa; 
        10'b0111100011: data <= 22'h002ed2; 
        10'b0111100100: data <= 22'h005a4b; 
        10'b0111100101: data <= 22'h004e46; 
        10'b0111100110: data <= 22'h001c5a; 
        10'b0111100111: data <= 22'h00164f; 
        10'b0111101000: data <= 22'h00204d; 
        10'b0111101001: data <= 22'h004d73; 
        10'b0111101010: data <= 22'h007ff4; 
        10'b0111101011: data <= 22'h006543; 
        10'b0111101100: data <= 22'h0054b5; 
        10'b0111101101: data <= 22'h001a2b; 
        10'b0111101110: data <= 22'h00040b; 
        10'b0111101111: data <= 22'h3fe3a7; 
        10'b0111110000: data <= 22'h00087d; 
        10'b0111110001: data <= 22'h00031b; 
        10'b0111110010: data <= 22'h3feead; 
        10'b0111110011: data <= 22'h3ff88b; 
        10'b0111110100: data <= 22'h3ff4b7; 
        10'b0111110101: data <= 22'h3ff98b; 
        10'b0111110110: data <= 22'h000b64; 
        10'b0111110111: data <= 22'h000ded; 
        10'b0111111000: data <= 22'h0006fb; 
        10'b0111111001: data <= 22'h000aaf; 
        10'b0111111010: data <= 22'h00095a; 
        10'b0111111011: data <= 22'h000165; 
        10'b0111111100: data <= 22'h3ff519; 
        10'b0111111101: data <= 22'h3fe90f; 
        10'b0111111110: data <= 22'h3fe55c; 
        10'b0111111111: data <= 22'h3fff7c; 
        10'b1000000000: data <= 22'h00171a; 
        10'b1000000001: data <= 22'h000547; 
        10'b1000000010: data <= 22'h3fed30; 
        10'b1000000011: data <= 22'h3ff4e0; 
        10'b1000000100: data <= 22'h001d88; 
        10'b1000000101: data <= 22'h00214a; 
        10'b1000000110: data <= 22'h00383b; 
        10'b1000000111: data <= 22'h00301c; 
        10'b1000001000: data <= 22'h001921; 
        10'b1000001001: data <= 22'h3fd915; 
        10'b1000001010: data <= 22'h3fdb23; 
        10'b1000001011: data <= 22'h3fc9f1; 
        10'b1000001100: data <= 22'h3fdfef; 
        10'b1000001101: data <= 22'h3fdebd; 
        10'b1000001110: data <= 22'h3fd3b2; 
        10'b1000001111: data <= 22'h3fddab; 
        10'b1000010000: data <= 22'h3ff70d; 
        10'b1000010001: data <= 22'h3ffb41; 
        10'b1000010010: data <= 22'h00041d; 
        10'b1000010011: data <= 22'h000092; 
        10'b1000010100: data <= 22'h0006c0; 
        10'b1000010101: data <= 22'h000c81; 
        10'b1000010110: data <= 22'h0004c2; 
        10'b1000010111: data <= 22'h0002da; 
        10'b1000011000: data <= 22'h3fe741; 
        10'b1000011001: data <= 22'h3fe141; 
        10'b1000011010: data <= 22'h3fd761; 
        10'b1000011011: data <= 22'h3fc2f8; 
        10'b1000011100: data <= 22'h3fbb2a; 
        10'b1000011101: data <= 22'h3fb6a3; 
        10'b1000011110: data <= 22'h3fa971; 
        10'b1000011111: data <= 22'h3fad35; 
        10'b1000100000: data <= 22'h3fb6af; 
        10'b1000100001: data <= 22'h3fd508; 
        10'b1000100010: data <= 22'h3ff33d; 
        10'b1000100011: data <= 22'h000b29; 
        10'b1000100100: data <= 22'h3fdeaa; 
        10'b1000100101: data <= 22'h3fe34e; 
        10'b1000100110: data <= 22'h3fdca8; 
        10'b1000100111: data <= 22'h3fcf3c; 
        10'b1000101000: data <= 22'h3fc97c; 
        10'b1000101001: data <= 22'h3fcdc9; 
        10'b1000101010: data <= 22'h3fccf7; 
        10'b1000101011: data <= 22'h3fdd7d; 
        10'b1000101100: data <= 22'h3ff6e7; 
        10'b1000101101: data <= 22'h0006d6; 
        10'b1000101110: data <= 22'h000c16; 
        10'b1000101111: data <= 22'h000b0b; 
        10'b1000110000: data <= 22'h0011fd; 
        10'b1000110001: data <= 22'h0010a7; 
        10'b1000110010: data <= 22'h0004d0; 
        10'b1000110011: data <= 22'h0002dd; 
        10'b1000110100: data <= 22'h3febec; 
        10'b1000110101: data <= 22'h3fdda5; 
        10'b1000110110: data <= 22'h3fce17; 
        10'b1000110111: data <= 22'h3faec4; 
        10'b1000111000: data <= 22'h3f9f71; 
        10'b1000111001: data <= 22'h3f99b0; 
        10'b1000111010: data <= 22'h3f97d0; 
        10'b1000111011: data <= 22'h3fb3b9; 
        10'b1000111100: data <= 22'h3fc252; 
        10'b1000111101: data <= 22'h3fbb0b; 
        10'b1000111110: data <= 22'h3fd4ab; 
        10'b1000111111: data <= 22'h3fe96b; 
        10'b1001000000: data <= 22'h3ff833; 
        10'b1001000001: data <= 22'h3ffba5; 
        10'b1001000010: data <= 22'h3fee17; 
        10'b1001000011: data <= 22'h3fd92f; 
        10'b1001000100: data <= 22'h3fe5e7; 
        10'b1001000101: data <= 22'h3fe277; 
        10'b1001000110: data <= 22'h3fdc5a; 
        10'b1001000111: data <= 22'h3fedb9; 
        10'b1001001000: data <= 22'h3fee73; 
        10'b1001001001: data <= 22'h00014b; 
        10'b1001001010: data <= 22'h00043c; 
        10'b1001001011: data <= 22'h000c07; 
        10'b1001001100: data <= 22'h000353; 
        10'b1001001101: data <= 22'h00053d; 
        10'b1001001110: data <= 22'h00015f; 
        10'b1001001111: data <= 22'h000265; 
        10'b1001010000: data <= 22'h3fffcc; 
        10'b1001010001: data <= 22'h3fec6d; 
        10'b1001010010: data <= 22'h3fced2; 
        10'b1001010011: data <= 22'h3fbb19; 
        10'b1001010100: data <= 22'h3fc1fb; 
        10'b1001010101: data <= 22'h3fb97a; 
        10'b1001010110: data <= 22'h3fc29b; 
        10'b1001010111: data <= 22'h3fd267; 
        10'b1001011000: data <= 22'h3fda15; 
        10'b1001011001: data <= 22'h3fdce0; 
        10'b1001011010: data <= 22'h3fd7c4; 
        10'b1001011011: data <= 22'h3fed64; 
        10'b1001011100: data <= 22'h3fe72f; 
        10'b1001011101: data <= 22'h000479; 
        10'b1001011110: data <= 22'h3ff898; 
        10'b1001011111: data <= 22'h000157; 
        10'b1001100000: data <= 22'h3ffcc5; 
        10'b1001100001: data <= 22'h3fe7da; 
        10'b1001100010: data <= 22'h3feb8a; 
        10'b1001100011: data <= 22'h3ffc3b; 
        10'b1001100100: data <= 22'h3fff57; 
        10'b1001100101: data <= 22'h000772; 
        10'b1001100110: data <= 22'h0009fe; 
        10'b1001100111: data <= 22'h0009a2; 
        10'b1001101000: data <= 22'h0008ab; 
        10'b1001101001: data <= 22'h000a13; 
        10'b1001101010: data <= 22'h000403; 
        10'b1001101011: data <= 22'h000b08; 
        10'b1001101100: data <= 22'h3ffd67; 
        10'b1001101101: data <= 22'h3ff590; 
        10'b1001101110: data <= 22'h3febb4; 
        10'b1001101111: data <= 22'h3fde7f; 
        10'b1001110000: data <= 22'h3fd2bb; 
        10'b1001110001: data <= 22'h3fe482; 
        10'b1001110010: data <= 22'h3fe3ab; 
        10'b1001110011: data <= 22'h3fec59; 
        10'b1001110100: data <= 22'h3feb47; 
        10'b1001110101: data <= 22'h3fee36; 
        10'b1001110110: data <= 22'h3fe9c8; 
        10'b1001110111: data <= 22'h3ff259; 
        10'b1001111000: data <= 22'h3ff2e7; 
        10'b1001111001: data <= 22'h0004b8; 
        10'b1001111010: data <= 22'h001414; 
        10'b1001111011: data <= 22'h0020c3; 
        10'b1001111100: data <= 22'h001925; 
        10'b1001111101: data <= 22'h00107d; 
        10'b1001111110: data <= 22'h3ff518; 
        10'b1001111111: data <= 22'h3ff548; 
        10'b1010000000: data <= 22'h3fff99; 
        10'b1010000001: data <= 22'h000731; 
        10'b1010000010: data <= 22'h000126; 
        10'b1010000011: data <= 22'h000584; 
        10'b1010000100: data <= 22'h00059d; 
        10'b1010000101: data <= 22'h000063; 
        10'b1010000110: data <= 22'h0004f8; 
        10'b1010000111: data <= 22'h0009d2; 
        10'b1010001000: data <= 22'h00058d; 
        10'b1010001001: data <= 22'h0006d0; 
        10'b1010001010: data <= 22'h3ff531; 
        10'b1010001011: data <= 22'h3ff3fa; 
        10'b1010001100: data <= 22'h3fefbc; 
        10'b1010001101: data <= 22'h000794; 
        10'b1010001110: data <= 22'h3fee81; 
        10'b1010001111: data <= 22'h0002d4; 
        10'b1010010000: data <= 22'h3fede7; 
        10'b1010010001: data <= 22'h3ff1c8; 
        10'b1010010010: data <= 22'h3ff21c; 
        10'b1010010011: data <= 22'h3ffefa; 
        10'b1010010100: data <= 22'h0004a0; 
        10'b1010010101: data <= 22'h000c3a; 
        10'b1010010110: data <= 22'h0025b0; 
        10'b1010010111: data <= 22'h0024c6; 
        10'b1010011000: data <= 22'h001f59; 
        10'b1010011001: data <= 22'h000df7; 
        10'b1010011010: data <= 22'h3ffad3; 
        10'b1010011011: data <= 22'h00043f; 
        10'b1010011100: data <= 22'h000850; 
        10'b1010011101: data <= 22'h000b61; 
        10'b1010011110: data <= 22'h0003b7; 
        10'b1010011111: data <= 22'h000e29; 
        10'b1010100000: data <= 22'h000ab4; 
        10'b1010100001: data <= 22'h000f4b; 
        10'b1010100010: data <= 22'h00073d; 
        10'b1010100011: data <= 22'h000c20; 
        10'b1010100100: data <= 22'h0002d9; 
        10'b1010100101: data <= 22'h000948; 
        10'b1010100110: data <= 22'h000387; 
        10'b1010100111: data <= 22'h3feec6; 
        10'b1010101000: data <= 22'h3fee69; 
        10'b1010101001: data <= 22'h3ffa65; 
        10'b1010101010: data <= 22'h3fed58; 
        10'b1010101011: data <= 22'h3ffcf5; 
        10'b1010101100: data <= 22'h3ff296; 
        10'b1010101101: data <= 22'h3ff3a4; 
        10'b1010101110: data <= 22'h3fe93f; 
        10'b1010101111: data <= 22'h3fe67a; 
        10'b1010110000: data <= 22'h3ff4fd; 
        10'b1010110001: data <= 22'h3ffa47; 
        10'b1010110010: data <= 22'h000201; 
        10'b1010110011: data <= 22'h0013d1; 
        10'b1010110100: data <= 22'h000e78; 
        10'b1010110101: data <= 22'h3ffa14; 
        10'b1010110110: data <= 22'h3ffe4b; 
        10'b1010110111: data <= 22'h0007a7; 
        10'b1010111000: data <= 22'h000c99; 
        10'b1010111001: data <= 22'h000203; 
        10'b1010111010: data <= 22'h000344; 
        10'b1010111011: data <= 22'h000ae7; 
        10'b1010111100: data <= 22'h001004; 
        10'b1010111101: data <= 22'h000f88; 
        10'b1010111110: data <= 22'h000e30; 
        10'b1010111111: data <= 22'h00032d; 
        10'b1011000000: data <= 22'h000e47; 
        10'b1011000001: data <= 22'h0000ae; 
        10'b1011000010: data <= 22'h3ff5cb; 
        10'b1011000011: data <= 22'h3fef63; 
        10'b1011000100: data <= 22'h3fe703; 
        10'b1011000101: data <= 22'h3fe5b7; 
        10'b1011000110: data <= 22'h3fd4d6; 
        10'b1011000111: data <= 22'h3fcf50; 
        10'b1011001000: data <= 22'h3fd206; 
        10'b1011001001: data <= 22'h3fd243; 
        10'b1011001010: data <= 22'h3fd922; 
        10'b1011001011: data <= 22'h3fd6dc; 
        10'b1011001100: data <= 22'h3fcac4; 
        10'b1011001101: data <= 22'h3fc352; 
        10'b1011001110: data <= 22'h3fc983; 
        10'b1011001111: data <= 22'h3fe223; 
        10'b1011010000: data <= 22'h3fe4b1; 
        10'b1011010001: data <= 22'h3ff623; 
        10'b1011010010: data <= 22'h00009c; 
        10'b1011010011: data <= 22'h000a72; 
        10'b1011010100: data <= 22'h0000c8; 
        10'b1011010101: data <= 22'h000e84; 
        10'b1011010110: data <= 22'h0005ce; 
        10'b1011010111: data <= 22'h000545; 
        10'b1011011000: data <= 22'h00077d; 
        10'b1011011001: data <= 22'h000acc; 
        10'b1011011010: data <= 22'h000271; 
        10'b1011011011: data <= 22'h000732; 
        10'b1011011100: data <= 22'h3fff47; 
        10'b1011011101: data <= 22'h3ffd86; 
        10'b1011011110: data <= 22'h000456; 
        10'b1011011111: data <= 22'h000321; 
        10'b1011100000: data <= 22'h3ffcb5; 
        10'b1011100001: data <= 22'h3ff0e2; 
        10'b1011100010: data <= 22'h3fdb8e; 
        10'b1011100011: data <= 22'h3fe034; 
        10'b1011100100: data <= 22'h3fdb9f; 
        10'b1011100101: data <= 22'h3fce97; 
        10'b1011100110: data <= 22'h3fca05; 
        10'b1011100111: data <= 22'h3fd5fd; 
        10'b1011101000: data <= 22'h3fd027; 
        10'b1011101001: data <= 22'h3fd75f; 
        10'b1011101010: data <= 22'h3fdea5; 
        10'b1011101011: data <= 22'h3fec20; 
        10'b1011101100: data <= 22'h3ff8b9; 
        10'b1011101101: data <= 22'h000ac4; 
        10'b1011101110: data <= 22'h000aab; 
        10'b1011101111: data <= 22'h000159; 
        10'b1011110000: data <= 22'h000700; 
        10'b1011110001: data <= 22'h000125; 
        10'b1011110010: data <= 22'h00112b; 
        10'b1011110011: data <= 22'h000784; 
        10'b1011110100: data <= 22'h000a6b; 
        10'b1011110101: data <= 22'h000187; 
        10'b1011110110: data <= 22'h000251; 
        10'b1011110111: data <= 22'h001081; 
        10'b1011111000: data <= 22'h000631; 
        10'b1011111001: data <= 22'h000dbe; 
        10'b1011111010: data <= 22'h000656; 
        10'b1011111011: data <= 22'h0010d5; 
        10'b1011111100: data <= 22'h3ffff7; 
        10'b1011111101: data <= 22'h000742; 
        10'b1011111110: data <= 22'h0003b7; 
        10'b1011111111: data <= 22'h3ffda9; 
        10'b1100000000: data <= 22'h3ffe49; 
        10'b1100000001: data <= 22'h00009e; 
        10'b1100000010: data <= 22'h3ff901; 
        10'b1100000011: data <= 22'h000d5a; 
        10'b1100000100: data <= 22'h3ffc93; 
        10'b1100000101: data <= 22'h3ffc16; 
        10'b1100000110: data <= 22'h3ffead; 
        10'b1100000111: data <= 22'h000708; 
        10'b1100001000: data <= 22'h000567; 
        10'b1100001001: data <= 22'h00055e; 
        10'b1100001010: data <= 22'h0005b4; 
        10'b1100001011: data <= 22'h0009be; 
        10'b1100001100: data <= 22'h000952; 
        10'b1100001101: data <= 22'h000c51; 
        10'b1100001110: data <= 22'h0008d4; 
        10'b1100001111: data <= 22'h0005dc; 
      endcase 
    end 
  end 
endgenerate 
assign dout = data; 
endmodule
