`timescale 1ns / 1ps 
 
////////////////////////////////////////////////////////////////////////////////// 
// WEIGHT MEMORY (ROM) 
////////////////////////////////////////////////////////////////////////////////// 
module ROM_weights_5 #( 
    parameter int WGHT_INT = 6, // integer part 
    parameter int WGHT_FRC = 16 // fractional part 
)( 
    input logic clk, // clock 
    input logic [9:0] address,
    output [WGHT_INT + WGHT_FRC-1:0] dout 
); 

(* rom_style = "block" *) reg [WGHT_INT + WGHT_FRC-1:0] data;
generate 
  if (WGHT_FRC == 1) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 7'h00; 
        10'b0000000001: data <= 7'h00; 
        10'b0000000010: data <= 7'h00; 
        10'b0000000011: data <= 7'h00; 
        10'b0000000100: data <= 7'h00; 
        10'b0000000101: data <= 7'h00; 
        10'b0000000110: data <= 7'h00; 
        10'b0000000111: data <= 7'h00; 
        10'b0000001000: data <= 7'h00; 
        10'b0000001001: data <= 7'h00; 
        10'b0000001010: data <= 7'h00; 
        10'b0000001011: data <= 7'h00; 
        10'b0000001100: data <= 7'h00; 
        10'b0000001101: data <= 7'h00; 
        10'b0000001110: data <= 7'h00; 
        10'b0000001111: data <= 7'h00; 
        10'b0000010000: data <= 7'h00; 
        10'b0000010001: data <= 7'h00; 
        10'b0000010010: data <= 7'h00; 
        10'b0000010011: data <= 7'h00; 
        10'b0000010100: data <= 7'h00; 
        10'b0000010101: data <= 7'h00; 
        10'b0000010110: data <= 7'h00; 
        10'b0000010111: data <= 7'h00; 
        10'b0000011000: data <= 7'h00; 
        10'b0000011001: data <= 7'h00; 
        10'b0000011010: data <= 7'h00; 
        10'b0000011011: data <= 7'h00; 
        10'b0000011100: data <= 7'h00; 
        10'b0000011101: data <= 7'h00; 
        10'b0000011110: data <= 7'h00; 
        10'b0000011111: data <= 7'h00; 
        10'b0000100000: data <= 7'h00; 
        10'b0000100001: data <= 7'h00; 
        10'b0000100010: data <= 7'h00; 
        10'b0000100011: data <= 7'h00; 
        10'b0000100100: data <= 7'h00; 
        10'b0000100101: data <= 7'h00; 
        10'b0000100110: data <= 7'h00; 
        10'b0000100111: data <= 7'h00; 
        10'b0000101000: data <= 7'h00; 
        10'b0000101001: data <= 7'h00; 
        10'b0000101010: data <= 7'h00; 
        10'b0000101011: data <= 7'h00; 
        10'b0000101100: data <= 7'h00; 
        10'b0000101101: data <= 7'h00; 
        10'b0000101110: data <= 7'h00; 
        10'b0000101111: data <= 7'h00; 
        10'b0000110000: data <= 7'h00; 
        10'b0000110001: data <= 7'h00; 
        10'b0000110010: data <= 7'h00; 
        10'b0000110011: data <= 7'h00; 
        10'b0000110100: data <= 7'h00; 
        10'b0000110101: data <= 7'h00; 
        10'b0000110110: data <= 7'h00; 
        10'b0000110111: data <= 7'h00; 
        10'b0000111000: data <= 7'h00; 
        10'b0000111001: data <= 7'h00; 
        10'b0000111010: data <= 7'h00; 
        10'b0000111011: data <= 7'h00; 
        10'b0000111100: data <= 7'h00; 
        10'b0000111101: data <= 7'h00; 
        10'b0000111110: data <= 7'h00; 
        10'b0000111111: data <= 7'h00; 
        10'b0001000000: data <= 7'h00; 
        10'b0001000001: data <= 7'h00; 
        10'b0001000010: data <= 7'h00; 
        10'b0001000011: data <= 7'h00; 
        10'b0001000100: data <= 7'h00; 
        10'b0001000101: data <= 7'h00; 
        10'b0001000110: data <= 7'h00; 
        10'b0001000111: data <= 7'h00; 
        10'b0001001000: data <= 7'h00; 
        10'b0001001001: data <= 7'h00; 
        10'b0001001010: data <= 7'h00; 
        10'b0001001011: data <= 7'h00; 
        10'b0001001100: data <= 7'h00; 
        10'b0001001101: data <= 7'h00; 
        10'b0001001110: data <= 7'h00; 
        10'b0001001111: data <= 7'h00; 
        10'b0001010000: data <= 7'h00; 
        10'b0001010001: data <= 7'h00; 
        10'b0001010010: data <= 7'h00; 
        10'b0001010011: data <= 7'h00; 
        10'b0001010100: data <= 7'h00; 
        10'b0001010101: data <= 7'h00; 
        10'b0001010110: data <= 7'h00; 
        10'b0001010111: data <= 7'h00; 
        10'b0001011000: data <= 7'h00; 
        10'b0001011001: data <= 7'h00; 
        10'b0001011010: data <= 7'h00; 
        10'b0001011011: data <= 7'h00; 
        10'b0001011100: data <= 7'h00; 
        10'b0001011101: data <= 7'h00; 
        10'b0001011110: data <= 7'h00; 
        10'b0001011111: data <= 7'h00; 
        10'b0001100000: data <= 7'h00; 
        10'b0001100001: data <= 7'h00; 
        10'b0001100010: data <= 7'h00; 
        10'b0001100011: data <= 7'h00; 
        10'b0001100100: data <= 7'h00; 
        10'b0001100101: data <= 7'h00; 
        10'b0001100110: data <= 7'h00; 
        10'b0001100111: data <= 7'h00; 
        10'b0001101000: data <= 7'h00; 
        10'b0001101001: data <= 7'h00; 
        10'b0001101010: data <= 7'h00; 
        10'b0001101011: data <= 7'h00; 
        10'b0001101100: data <= 7'h00; 
        10'b0001101101: data <= 7'h00; 
        10'b0001101110: data <= 7'h00; 
        10'b0001101111: data <= 7'h00; 
        10'b0001110000: data <= 7'h00; 
        10'b0001110001: data <= 7'h00; 
        10'b0001110010: data <= 7'h00; 
        10'b0001110011: data <= 7'h00; 
        10'b0001110100: data <= 7'h00; 
        10'b0001110101: data <= 7'h00; 
        10'b0001110110: data <= 7'h00; 
        10'b0001110111: data <= 7'h00; 
        10'b0001111000: data <= 7'h00; 
        10'b0001111001: data <= 7'h00; 
        10'b0001111010: data <= 7'h7f; 
        10'b0001111011: data <= 7'h00; 
        10'b0001111100: data <= 7'h00; 
        10'b0001111101: data <= 7'h00; 
        10'b0001111110: data <= 7'h00; 
        10'b0001111111: data <= 7'h00; 
        10'b0010000000: data <= 7'h00; 
        10'b0010000001: data <= 7'h00; 
        10'b0010000010: data <= 7'h00; 
        10'b0010000011: data <= 7'h00; 
        10'b0010000100: data <= 7'h00; 
        10'b0010000101: data <= 7'h00; 
        10'b0010000110: data <= 7'h00; 
        10'b0010000111: data <= 7'h00; 
        10'b0010001000: data <= 7'h00; 
        10'b0010001001: data <= 7'h00; 
        10'b0010001010: data <= 7'h00; 
        10'b0010001011: data <= 7'h00; 
        10'b0010001100: data <= 7'h00; 
        10'b0010001101: data <= 7'h00; 
        10'b0010001110: data <= 7'h00; 
        10'b0010001111: data <= 7'h00; 
        10'b0010010000: data <= 7'h00; 
        10'b0010010001: data <= 7'h00; 
        10'b0010010010: data <= 7'h00; 
        10'b0010010011: data <= 7'h00; 
        10'b0010010100: data <= 7'h00; 
        10'b0010010101: data <= 7'h00; 
        10'b0010010110: data <= 7'h00; 
        10'b0010010111: data <= 7'h00; 
        10'b0010011000: data <= 7'h00; 
        10'b0010011001: data <= 7'h00; 
        10'b0010011010: data <= 7'h00; 
        10'b0010011011: data <= 7'h00; 
        10'b0010011100: data <= 7'h00; 
        10'b0010011101: data <= 7'h00; 
        10'b0010011110: data <= 7'h00; 
        10'b0010011111: data <= 7'h00; 
        10'b0010100000: data <= 7'h00; 
        10'b0010100001: data <= 7'h00; 
        10'b0010100010: data <= 7'h00; 
        10'b0010100011: data <= 7'h00; 
        10'b0010100100: data <= 7'h00; 
        10'b0010100101: data <= 7'h00; 
        10'b0010100110: data <= 7'h00; 
        10'b0010100111: data <= 7'h00; 
        10'b0010101000: data <= 7'h00; 
        10'b0010101001: data <= 7'h00; 
        10'b0010101010: data <= 7'h00; 
        10'b0010101011: data <= 7'h00; 
        10'b0010101100: data <= 7'h00; 
        10'b0010101101: data <= 7'h00; 
        10'b0010101110: data <= 7'h00; 
        10'b0010101111: data <= 7'h00; 
        10'b0010110000: data <= 7'h00; 
        10'b0010110001: data <= 7'h00; 
        10'b0010110010: data <= 7'h00; 
        10'b0010110011: data <= 7'h00; 
        10'b0010110100: data <= 7'h00; 
        10'b0010110101: data <= 7'h00; 
        10'b0010110110: data <= 7'h00; 
        10'b0010110111: data <= 7'h00; 
        10'b0010111000: data <= 7'h00; 
        10'b0010111001: data <= 7'h00; 
        10'b0010111010: data <= 7'h00; 
        10'b0010111011: data <= 7'h00; 
        10'b0010111100: data <= 7'h00; 
        10'b0010111101: data <= 7'h00; 
        10'b0010111110: data <= 7'h00; 
        10'b0010111111: data <= 7'h01; 
        10'b0011000000: data <= 7'h01; 
        10'b0011000001: data <= 7'h00; 
        10'b0011000010: data <= 7'h00; 
        10'b0011000011: data <= 7'h00; 
        10'b0011000100: data <= 7'h00; 
        10'b0011000101: data <= 7'h00; 
        10'b0011000110: data <= 7'h00; 
        10'b0011000111: data <= 7'h00; 
        10'b0011001000: data <= 7'h00; 
        10'b0011001001: data <= 7'h00; 
        10'b0011001010: data <= 7'h00; 
        10'b0011001011: data <= 7'h00; 
        10'b0011001100: data <= 7'h00; 
        10'b0011001101: data <= 7'h00; 
        10'b0011001110: data <= 7'h00; 
        10'b0011001111: data <= 7'h00; 
        10'b0011010000: data <= 7'h00; 
        10'b0011010001: data <= 7'h00; 
        10'b0011010010: data <= 7'h00; 
        10'b0011010011: data <= 7'h00; 
        10'b0011010100: data <= 7'h00; 
        10'b0011010101: data <= 7'h00; 
        10'b0011010110: data <= 7'h00; 
        10'b0011010111: data <= 7'h00; 
        10'b0011011000: data <= 7'h00; 
        10'b0011011001: data <= 7'h00; 
        10'b0011011010: data <= 7'h01; 
        10'b0011011011: data <= 7'h01; 
        10'b0011011100: data <= 7'h01; 
        10'b0011011101: data <= 7'h01; 
        10'b0011011110: data <= 7'h00; 
        10'b0011011111: data <= 7'h00; 
        10'b0011100000: data <= 7'h00; 
        10'b0011100001: data <= 7'h00; 
        10'b0011100010: data <= 7'h00; 
        10'b0011100011: data <= 7'h00; 
        10'b0011100100: data <= 7'h7f; 
        10'b0011100101: data <= 7'h00; 
        10'b0011100110: data <= 7'h00; 
        10'b0011100111: data <= 7'h00; 
        10'b0011101000: data <= 7'h00; 
        10'b0011101001: data <= 7'h00; 
        10'b0011101010: data <= 7'h00; 
        10'b0011101011: data <= 7'h00; 
        10'b0011101100: data <= 7'h00; 
        10'b0011101101: data <= 7'h00; 
        10'b0011101110: data <= 7'h00; 
        10'b0011101111: data <= 7'h00; 
        10'b0011110000: data <= 7'h00; 
        10'b0011110001: data <= 7'h00; 
        10'b0011110010: data <= 7'h00; 
        10'b0011110011: data <= 7'h00; 
        10'b0011110100: data <= 7'h00; 
        10'b0011110101: data <= 7'h00; 
        10'b0011110110: data <= 7'h01; 
        10'b0011110111: data <= 7'h01; 
        10'b0011111000: data <= 7'h01; 
        10'b0011111001: data <= 7'h01; 
        10'b0011111010: data <= 7'h00; 
        10'b0011111011: data <= 7'h00; 
        10'b0011111100: data <= 7'h00; 
        10'b0011111101: data <= 7'h00; 
        10'b0011111110: data <= 7'h00; 
        10'b0011111111: data <= 7'h00; 
        10'b0100000000: data <= 7'h00; 
        10'b0100000001: data <= 7'h00; 
        10'b0100000010: data <= 7'h00; 
        10'b0100000011: data <= 7'h00; 
        10'b0100000100: data <= 7'h00; 
        10'b0100000101: data <= 7'h00; 
        10'b0100000110: data <= 7'h00; 
        10'b0100000111: data <= 7'h01; 
        10'b0100001000: data <= 7'h00; 
        10'b0100001001: data <= 7'h00; 
        10'b0100001010: data <= 7'h00; 
        10'b0100001011: data <= 7'h7f; 
        10'b0100001100: data <= 7'h7f; 
        10'b0100001101: data <= 7'h00; 
        10'b0100001110: data <= 7'h00; 
        10'b0100001111: data <= 7'h00; 
        10'b0100010000: data <= 7'h00; 
        10'b0100010001: data <= 7'h01; 
        10'b0100010010: data <= 7'h01; 
        10'b0100010011: data <= 7'h01; 
        10'b0100010100: data <= 7'h02; 
        10'b0100010101: data <= 7'h01; 
        10'b0100010110: data <= 7'h00; 
        10'b0100010111: data <= 7'h00; 
        10'b0100011000: data <= 7'h00; 
        10'b0100011001: data <= 7'h00; 
        10'b0100011010: data <= 7'h00; 
        10'b0100011011: data <= 7'h00; 
        10'b0100011100: data <= 7'h00; 
        10'b0100011101: data <= 7'h00; 
        10'b0100011110: data <= 7'h00; 
        10'b0100011111: data <= 7'h00; 
        10'b0100100000: data <= 7'h00; 
        10'b0100100001: data <= 7'h01; 
        10'b0100100010: data <= 7'h01; 
        10'b0100100011: data <= 7'h01; 
        10'b0100100100: data <= 7'h01; 
        10'b0100100101: data <= 7'h00; 
        10'b0100100110: data <= 7'h00; 
        10'b0100100111: data <= 7'h00; 
        10'b0100101000: data <= 7'h7f; 
        10'b0100101001: data <= 7'h7f; 
        10'b0100101010: data <= 7'h7f; 
        10'b0100101011: data <= 7'h7f; 
        10'b0100101100: data <= 7'h00; 
        10'b0100101101: data <= 7'h00; 
        10'b0100101110: data <= 7'h00; 
        10'b0100101111: data <= 7'h00; 
        10'b0100110000: data <= 7'h01; 
        10'b0100110001: data <= 7'h01; 
        10'b0100110010: data <= 7'h00; 
        10'b0100110011: data <= 7'h00; 
        10'b0100110100: data <= 7'h00; 
        10'b0100110101: data <= 7'h00; 
        10'b0100110110: data <= 7'h00; 
        10'b0100110111: data <= 7'h00; 
        10'b0100111000: data <= 7'h00; 
        10'b0100111001: data <= 7'h00; 
        10'b0100111010: data <= 7'h00; 
        10'b0100111011: data <= 7'h00; 
        10'b0100111100: data <= 7'h00; 
        10'b0100111101: data <= 7'h00; 
        10'b0100111110: data <= 7'h00; 
        10'b0100111111: data <= 7'h00; 
        10'b0101000000: data <= 7'h01; 
        10'b0101000001: data <= 7'h01; 
        10'b0101000010: data <= 7'h00; 
        10'b0101000011: data <= 7'h00; 
        10'b0101000100: data <= 7'h00; 
        10'b0101000101: data <= 7'h00; 
        10'b0101000110: data <= 7'h7f; 
        10'b0101000111: data <= 7'h7f; 
        10'b0101001000: data <= 7'h7f; 
        10'b0101001001: data <= 7'h7f; 
        10'b0101001010: data <= 7'h7f; 
        10'b0101001011: data <= 7'h7f; 
        10'b0101001100: data <= 7'h00; 
        10'b0101001101: data <= 7'h00; 
        10'b0101001110: data <= 7'h00; 
        10'b0101001111: data <= 7'h00; 
        10'b0101010000: data <= 7'h00; 
        10'b0101010001: data <= 7'h00; 
        10'b0101010010: data <= 7'h00; 
        10'b0101010011: data <= 7'h00; 
        10'b0101010100: data <= 7'h00; 
        10'b0101010101: data <= 7'h00; 
        10'b0101010110: data <= 7'h00; 
        10'b0101010111: data <= 7'h00; 
        10'b0101011000: data <= 7'h00; 
        10'b0101011001: data <= 7'h00; 
        10'b0101011010: data <= 7'h00; 
        10'b0101011011: data <= 7'h01; 
        10'b0101011100: data <= 7'h01; 
        10'b0101011101: data <= 7'h01; 
        10'b0101011110: data <= 7'h00; 
        10'b0101011111: data <= 7'h00; 
        10'b0101100000: data <= 7'h7f; 
        10'b0101100001: data <= 7'h7f; 
        10'b0101100010: data <= 7'h00; 
        10'b0101100011: data <= 7'h7f; 
        10'b0101100100: data <= 7'h7f; 
        10'b0101100101: data <= 7'h7f; 
        10'b0101100110: data <= 7'h7f; 
        10'b0101100111: data <= 7'h7f; 
        10'b0101101000: data <= 7'h7f; 
        10'b0101101001: data <= 7'h00; 
        10'b0101101010: data <= 7'h00; 
        10'b0101101011: data <= 7'h00; 
        10'b0101101100: data <= 7'h00; 
        10'b0101101101: data <= 7'h00; 
        10'b0101101110: data <= 7'h00; 
        10'b0101101111: data <= 7'h00; 
        10'b0101110000: data <= 7'h00; 
        10'b0101110001: data <= 7'h00; 
        10'b0101110010: data <= 7'h00; 
        10'b0101110011: data <= 7'h00; 
        10'b0101110100: data <= 7'h00; 
        10'b0101110101: data <= 7'h00; 
        10'b0101110110: data <= 7'h00; 
        10'b0101110111: data <= 7'h01; 
        10'b0101111000: data <= 7'h00; 
        10'b0101111001: data <= 7'h00; 
        10'b0101111010: data <= 7'h00; 
        10'b0101111011: data <= 7'h00; 
        10'b0101111100: data <= 7'h7f; 
        10'b0101111101: data <= 7'h00; 
        10'b0101111110: data <= 7'h00; 
        10'b0101111111: data <= 7'h00; 
        10'b0110000000: data <= 7'h00; 
        10'b0110000001: data <= 7'h00; 
        10'b0110000010: data <= 7'h00; 
        10'b0110000011: data <= 7'h7f; 
        10'b0110000100: data <= 7'h7f; 
        10'b0110000101: data <= 7'h00; 
        10'b0110000110: data <= 7'h00; 
        10'b0110000111: data <= 7'h00; 
        10'b0110001000: data <= 7'h00; 
        10'b0110001001: data <= 7'h00; 
        10'b0110001010: data <= 7'h00; 
        10'b0110001011: data <= 7'h00; 
        10'b0110001100: data <= 7'h00; 
        10'b0110001101: data <= 7'h00; 
        10'b0110001110: data <= 7'h00; 
        10'b0110001111: data <= 7'h00; 
        10'b0110010000: data <= 7'h00; 
        10'b0110010001: data <= 7'h00; 
        10'b0110010010: data <= 7'h00; 
        10'b0110010011: data <= 7'h00; 
        10'b0110010100: data <= 7'h00; 
        10'b0110010101: data <= 7'h00; 
        10'b0110010110: data <= 7'h00; 
        10'b0110010111: data <= 7'h00; 
        10'b0110011000: data <= 7'h00; 
        10'b0110011001: data <= 7'h00; 
        10'b0110011010: data <= 7'h00; 
        10'b0110011011: data <= 7'h00; 
        10'b0110011100: data <= 7'h00; 
        10'b0110011101: data <= 7'h00; 
        10'b0110011110: data <= 7'h00; 
        10'b0110011111: data <= 7'h00; 
        10'b0110100000: data <= 7'h00; 
        10'b0110100001: data <= 7'h00; 
        10'b0110100010: data <= 7'h00; 
        10'b0110100011: data <= 7'h00; 
        10'b0110100100: data <= 7'h00; 
        10'b0110100101: data <= 7'h00; 
        10'b0110100110: data <= 7'h00; 
        10'b0110100111: data <= 7'h00; 
        10'b0110101000: data <= 7'h00; 
        10'b0110101001: data <= 7'h00; 
        10'b0110101010: data <= 7'h00; 
        10'b0110101011: data <= 7'h00; 
        10'b0110101100: data <= 7'h00; 
        10'b0110101101: data <= 7'h00; 
        10'b0110101110: data <= 7'h00; 
        10'b0110101111: data <= 7'h00; 
        10'b0110110000: data <= 7'h00; 
        10'b0110110001: data <= 7'h00; 
        10'b0110110010: data <= 7'h00; 
        10'b0110110011: data <= 7'h7f; 
        10'b0110110100: data <= 7'h00; 
        10'b0110110101: data <= 7'h00; 
        10'b0110110110: data <= 7'h00; 
        10'b0110110111: data <= 7'h00; 
        10'b0110111000: data <= 7'h00; 
        10'b0110111001: data <= 7'h00; 
        10'b0110111010: data <= 7'h00; 
        10'b0110111011: data <= 7'h00; 
        10'b0110111100: data <= 7'h00; 
        10'b0110111101: data <= 7'h00; 
        10'b0110111110: data <= 7'h00; 
        10'b0110111111: data <= 7'h00; 
        10'b0111000000: data <= 7'h00; 
        10'b0111000001: data <= 7'h00; 
        10'b0111000010: data <= 7'h00; 
        10'b0111000011: data <= 7'h00; 
        10'b0111000100: data <= 7'h00; 
        10'b0111000101: data <= 7'h00; 
        10'b0111000110: data <= 7'h7f; 
        10'b0111000111: data <= 7'h7f; 
        10'b0111001000: data <= 7'h00; 
        10'b0111001001: data <= 7'h00; 
        10'b0111001010: data <= 7'h00; 
        10'b0111001011: data <= 7'h00; 
        10'b0111001100: data <= 7'h00; 
        10'b0111001101: data <= 7'h00; 
        10'b0111001110: data <= 7'h7f; 
        10'b0111001111: data <= 7'h00; 
        10'b0111010000: data <= 7'h00; 
        10'b0111010001: data <= 7'h00; 
        10'b0111010010: data <= 7'h00; 
        10'b0111010011: data <= 7'h00; 
        10'b0111010100: data <= 7'h00; 
        10'b0111010101: data <= 7'h00; 
        10'b0111010110: data <= 7'h00; 
        10'b0111010111: data <= 7'h00; 
        10'b0111011000: data <= 7'h00; 
        10'b0111011001: data <= 7'h00; 
        10'b0111011010: data <= 7'h00; 
        10'b0111011011: data <= 7'h00; 
        10'b0111011100: data <= 7'h00; 
        10'b0111011101: data <= 7'h00; 
        10'b0111011110: data <= 7'h00; 
        10'b0111011111: data <= 7'h00; 
        10'b0111100000: data <= 7'h00; 
        10'b0111100001: data <= 7'h00; 
        10'b0111100010: data <= 7'h00; 
        10'b0111100011: data <= 7'h00; 
        10'b0111100100: data <= 7'h7f; 
        10'b0111100101: data <= 7'h7f; 
        10'b0111100110: data <= 7'h7f; 
        10'b0111100111: data <= 7'h00; 
        10'b0111101000: data <= 7'h7f; 
        10'b0111101001: data <= 7'h7f; 
        10'b0111101010: data <= 7'h7f; 
        10'b0111101011: data <= 7'h00; 
        10'b0111101100: data <= 7'h00; 
        10'b0111101101: data <= 7'h00; 
        10'b0111101110: data <= 7'h00; 
        10'b0111101111: data <= 7'h00; 
        10'b0111110000: data <= 7'h00; 
        10'b0111110001: data <= 7'h00; 
        10'b0111110010: data <= 7'h00; 
        10'b0111110011: data <= 7'h00; 
        10'b0111110100: data <= 7'h00; 
        10'b0111110101: data <= 7'h00; 
        10'b0111110110: data <= 7'h00; 
        10'b0111110111: data <= 7'h00; 
        10'b0111111000: data <= 7'h00; 
        10'b0111111001: data <= 7'h00; 
        10'b0111111010: data <= 7'h00; 
        10'b0111111011: data <= 7'h00; 
        10'b0111111100: data <= 7'h00; 
        10'b0111111101: data <= 7'h00; 
        10'b0111111110: data <= 7'h01; 
        10'b0111111111: data <= 7'h00; 
        10'b1000000000: data <= 7'h00; 
        10'b1000000001: data <= 7'h7f; 
        10'b1000000010: data <= 7'h7f; 
        10'b1000000011: data <= 7'h7f; 
        10'b1000000100: data <= 7'h7f; 
        10'b1000000101: data <= 7'h00; 
        10'b1000000110: data <= 7'h00; 
        10'b1000000111: data <= 7'h00; 
        10'b1000001000: data <= 7'h00; 
        10'b1000001001: data <= 7'h00; 
        10'b1000001010: data <= 7'h00; 
        10'b1000001011: data <= 7'h00; 
        10'b1000001100: data <= 7'h00; 
        10'b1000001101: data <= 7'h00; 
        10'b1000001110: data <= 7'h00; 
        10'b1000001111: data <= 7'h00; 
        10'b1000010000: data <= 7'h00; 
        10'b1000010001: data <= 7'h00; 
        10'b1000010010: data <= 7'h00; 
        10'b1000010011: data <= 7'h00; 
        10'b1000010100: data <= 7'h00; 
        10'b1000010101: data <= 7'h00; 
        10'b1000010110: data <= 7'h00; 
        10'b1000010111: data <= 7'h00; 
        10'b1000011000: data <= 7'h00; 
        10'b1000011001: data <= 7'h00; 
        10'b1000011010: data <= 7'h01; 
        10'b1000011011: data <= 7'h00; 
        10'b1000011100: data <= 7'h00; 
        10'b1000011101: data <= 7'h00; 
        10'b1000011110: data <= 7'h00; 
        10'b1000011111: data <= 7'h00; 
        10'b1000100000: data <= 7'h00; 
        10'b1000100001: data <= 7'h00; 
        10'b1000100010: data <= 7'h00; 
        10'b1000100011: data <= 7'h00; 
        10'b1000100100: data <= 7'h00; 
        10'b1000100101: data <= 7'h00; 
        10'b1000100110: data <= 7'h00; 
        10'b1000100111: data <= 7'h00; 
        10'b1000101000: data <= 7'h00; 
        10'b1000101001: data <= 7'h00; 
        10'b1000101010: data <= 7'h00; 
        10'b1000101011: data <= 7'h00; 
        10'b1000101100: data <= 7'h00; 
        10'b1000101101: data <= 7'h00; 
        10'b1000101110: data <= 7'h00; 
        10'b1000101111: data <= 7'h00; 
        10'b1000110000: data <= 7'h00; 
        10'b1000110001: data <= 7'h00; 
        10'b1000110010: data <= 7'h00; 
        10'b1000110011: data <= 7'h00; 
        10'b1000110100: data <= 7'h00; 
        10'b1000110101: data <= 7'h00; 
        10'b1000110110: data <= 7'h00; 
        10'b1000110111: data <= 7'h00; 
        10'b1000111000: data <= 7'h01; 
        10'b1000111001: data <= 7'h00; 
        10'b1000111010: data <= 7'h00; 
        10'b1000111011: data <= 7'h01; 
        10'b1000111100: data <= 7'h00; 
        10'b1000111101: data <= 7'h00; 
        10'b1000111110: data <= 7'h00; 
        10'b1000111111: data <= 7'h00; 
        10'b1001000000: data <= 7'h00; 
        10'b1001000001: data <= 7'h00; 
        10'b1001000010: data <= 7'h00; 
        10'b1001000011: data <= 7'h00; 
        10'b1001000100: data <= 7'h00; 
        10'b1001000101: data <= 7'h00; 
        10'b1001000110: data <= 7'h00; 
        10'b1001000111: data <= 7'h00; 
        10'b1001001000: data <= 7'h00; 
        10'b1001001001: data <= 7'h00; 
        10'b1001001010: data <= 7'h00; 
        10'b1001001011: data <= 7'h00; 
        10'b1001001100: data <= 7'h00; 
        10'b1001001101: data <= 7'h00; 
        10'b1001001110: data <= 7'h00; 
        10'b1001001111: data <= 7'h00; 
        10'b1001010000: data <= 7'h00; 
        10'b1001010001: data <= 7'h00; 
        10'b1001010010: data <= 7'h00; 
        10'b1001010011: data <= 7'h00; 
        10'b1001010100: data <= 7'h01; 
        10'b1001010101: data <= 7'h00; 
        10'b1001010110: data <= 7'h00; 
        10'b1001010111: data <= 7'h00; 
        10'b1001011000: data <= 7'h00; 
        10'b1001011001: data <= 7'h00; 
        10'b1001011010: data <= 7'h00; 
        10'b1001011011: data <= 7'h00; 
        10'b1001011100: data <= 7'h00; 
        10'b1001011101: data <= 7'h00; 
        10'b1001011110: data <= 7'h00; 
        10'b1001011111: data <= 7'h00; 
        10'b1001100000: data <= 7'h00; 
        10'b1001100001: data <= 7'h00; 
        10'b1001100010: data <= 7'h00; 
        10'b1001100011: data <= 7'h00; 
        10'b1001100100: data <= 7'h00; 
        10'b1001100101: data <= 7'h00; 
        10'b1001100110: data <= 7'h00; 
        10'b1001100111: data <= 7'h00; 
        10'b1001101000: data <= 7'h00; 
        10'b1001101001: data <= 7'h00; 
        10'b1001101010: data <= 7'h00; 
        10'b1001101011: data <= 7'h00; 
        10'b1001101100: data <= 7'h00; 
        10'b1001101101: data <= 7'h00; 
        10'b1001101110: data <= 7'h00; 
        10'b1001101111: data <= 7'h00; 
        10'b1001110000: data <= 7'h00; 
        10'b1001110001: data <= 7'h00; 
        10'b1001110010: data <= 7'h00; 
        10'b1001110011: data <= 7'h00; 
        10'b1001110100: data <= 7'h00; 
        10'b1001110101: data <= 7'h01; 
        10'b1001110110: data <= 7'h00; 
        10'b1001110111: data <= 7'h00; 
        10'b1001111000: data <= 7'h00; 
        10'b1001111001: data <= 7'h00; 
        10'b1001111010: data <= 7'h00; 
        10'b1001111011: data <= 7'h00; 
        10'b1001111100: data <= 7'h00; 
        10'b1001111101: data <= 7'h00; 
        10'b1001111110: data <= 7'h00; 
        10'b1001111111: data <= 7'h00; 
        10'b1010000000: data <= 7'h00; 
        10'b1010000001: data <= 7'h00; 
        10'b1010000010: data <= 7'h00; 
        10'b1010000011: data <= 7'h00; 
        10'b1010000100: data <= 7'h00; 
        10'b1010000101: data <= 7'h00; 
        10'b1010000110: data <= 7'h00; 
        10'b1010000111: data <= 7'h00; 
        10'b1010001000: data <= 7'h00; 
        10'b1010001001: data <= 7'h00; 
        10'b1010001010: data <= 7'h00; 
        10'b1010001011: data <= 7'h00; 
        10'b1010001100: data <= 7'h00; 
        10'b1010001101: data <= 7'h00; 
        10'b1010001110: data <= 7'h00; 
        10'b1010001111: data <= 7'h00; 
        10'b1010010000: data <= 7'h00; 
        10'b1010010001: data <= 7'h00; 
        10'b1010010010: data <= 7'h00; 
        10'b1010010011: data <= 7'h00; 
        10'b1010010100: data <= 7'h00; 
        10'b1010010101: data <= 7'h00; 
        10'b1010010110: data <= 7'h00; 
        10'b1010010111: data <= 7'h00; 
        10'b1010011000: data <= 7'h00; 
        10'b1010011001: data <= 7'h00; 
        10'b1010011010: data <= 7'h00; 
        10'b1010011011: data <= 7'h00; 
        10'b1010011100: data <= 7'h00; 
        10'b1010011101: data <= 7'h00; 
        10'b1010011110: data <= 7'h00; 
        10'b1010011111: data <= 7'h00; 
        10'b1010100000: data <= 7'h00; 
        10'b1010100001: data <= 7'h00; 
        10'b1010100010: data <= 7'h00; 
        10'b1010100011: data <= 7'h00; 
        10'b1010100100: data <= 7'h00; 
        10'b1010100101: data <= 7'h00; 
        10'b1010100110: data <= 7'h00; 
        10'b1010100111: data <= 7'h00; 
        10'b1010101000: data <= 7'h00; 
        10'b1010101001: data <= 7'h00; 
        10'b1010101010: data <= 7'h00; 
        10'b1010101011: data <= 7'h00; 
        10'b1010101100: data <= 7'h00; 
        10'b1010101101: data <= 7'h00; 
        10'b1010101110: data <= 7'h00; 
        10'b1010101111: data <= 7'h00; 
        10'b1010110000: data <= 7'h00; 
        10'b1010110001: data <= 7'h00; 
        10'b1010110010: data <= 7'h00; 
        10'b1010110011: data <= 7'h00; 
        10'b1010110100: data <= 7'h00; 
        10'b1010110101: data <= 7'h00; 
        10'b1010110110: data <= 7'h00; 
        10'b1010110111: data <= 7'h00; 
        10'b1010111000: data <= 7'h00; 
        10'b1010111001: data <= 7'h00; 
        10'b1010111010: data <= 7'h00; 
        10'b1010111011: data <= 7'h00; 
        10'b1010111100: data <= 7'h00; 
        10'b1010111101: data <= 7'h00; 
        10'b1010111110: data <= 7'h00; 
        10'b1010111111: data <= 7'h00; 
        10'b1011000000: data <= 7'h00; 
        10'b1011000001: data <= 7'h00; 
        10'b1011000010: data <= 7'h00; 
        10'b1011000011: data <= 7'h00; 
        10'b1011000100: data <= 7'h00; 
        10'b1011000101: data <= 7'h00; 
        10'b1011000110: data <= 7'h00; 
        10'b1011000111: data <= 7'h00; 
        10'b1011001000: data <= 7'h00; 
        10'b1011001001: data <= 7'h00; 
        10'b1011001010: data <= 7'h00; 
        10'b1011001011: data <= 7'h00; 
        10'b1011001100: data <= 7'h00; 
        10'b1011001101: data <= 7'h00; 
        10'b1011001110: data <= 7'h00; 
        10'b1011001111: data <= 7'h00; 
        10'b1011010000: data <= 7'h00; 
        10'b1011010001: data <= 7'h00; 
        10'b1011010010: data <= 7'h00; 
        10'b1011010011: data <= 7'h00; 
        10'b1011010100: data <= 7'h00; 
        10'b1011010101: data <= 7'h00; 
        10'b1011010110: data <= 7'h00; 
        10'b1011010111: data <= 7'h00; 
        10'b1011011000: data <= 7'h00; 
        10'b1011011001: data <= 7'h00; 
        10'b1011011010: data <= 7'h00; 
        10'b1011011011: data <= 7'h00; 
        10'b1011011100: data <= 7'h00; 
        10'b1011011101: data <= 7'h00; 
        10'b1011011110: data <= 7'h00; 
        10'b1011011111: data <= 7'h00; 
        10'b1011100000: data <= 7'h00; 
        10'b1011100001: data <= 7'h00; 
        10'b1011100010: data <= 7'h00; 
        10'b1011100011: data <= 7'h00; 
        10'b1011100100: data <= 7'h00; 
        10'b1011100101: data <= 7'h00; 
        10'b1011100110: data <= 7'h00; 
        10'b1011100111: data <= 7'h00; 
        10'b1011101000: data <= 7'h00; 
        10'b1011101001: data <= 7'h00; 
        10'b1011101010: data <= 7'h00; 
        10'b1011101011: data <= 7'h00; 
        10'b1011101100: data <= 7'h00; 
        10'b1011101101: data <= 7'h00; 
        10'b1011101110: data <= 7'h00; 
        10'b1011101111: data <= 7'h00; 
        10'b1011110000: data <= 7'h00; 
        10'b1011110001: data <= 7'h00; 
        10'b1011110010: data <= 7'h00; 
        10'b1011110011: data <= 7'h00; 
        10'b1011110100: data <= 7'h00; 
        10'b1011110101: data <= 7'h00; 
        10'b1011110110: data <= 7'h00; 
        10'b1011110111: data <= 7'h00; 
        10'b1011111000: data <= 7'h00; 
        10'b1011111001: data <= 7'h00; 
        10'b1011111010: data <= 7'h00; 
        10'b1011111011: data <= 7'h00; 
        10'b1011111100: data <= 7'h00; 
        10'b1011111101: data <= 7'h00; 
        10'b1011111110: data <= 7'h00; 
        10'b1011111111: data <= 7'h00; 
        10'b1100000000: data <= 7'h00; 
        10'b1100000001: data <= 7'h00; 
        10'b1100000010: data <= 7'h00; 
        10'b1100000011: data <= 7'h00; 
        10'b1100000100: data <= 7'h00; 
        10'b1100000101: data <= 7'h00; 
        10'b1100000110: data <= 7'h00; 
        10'b1100000111: data <= 7'h00; 
        10'b1100001000: data <= 7'h00; 
        10'b1100001001: data <= 7'h00; 
        10'b1100001010: data <= 7'h00; 
        10'b1100001011: data <= 7'h00; 
        10'b1100001100: data <= 7'h00; 
        10'b1100001101: data <= 7'h00; 
        10'b1100001110: data <= 7'h00; 
        10'b1100001111: data <= 7'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 2) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 8'h00; 
        10'b0000000001: data <= 8'h00; 
        10'b0000000010: data <= 8'h00; 
        10'b0000000011: data <= 8'h00; 
        10'b0000000100: data <= 8'h00; 
        10'b0000000101: data <= 8'h00; 
        10'b0000000110: data <= 8'h00; 
        10'b0000000111: data <= 8'h00; 
        10'b0000001000: data <= 8'h00; 
        10'b0000001001: data <= 8'h00; 
        10'b0000001010: data <= 8'h00; 
        10'b0000001011: data <= 8'h00; 
        10'b0000001100: data <= 8'h00; 
        10'b0000001101: data <= 8'h00; 
        10'b0000001110: data <= 8'h00; 
        10'b0000001111: data <= 8'h00; 
        10'b0000010000: data <= 8'h00; 
        10'b0000010001: data <= 8'h00; 
        10'b0000010010: data <= 8'h00; 
        10'b0000010011: data <= 8'h00; 
        10'b0000010100: data <= 8'h00; 
        10'b0000010101: data <= 8'h00; 
        10'b0000010110: data <= 8'h00; 
        10'b0000010111: data <= 8'h00; 
        10'b0000011000: data <= 8'h00; 
        10'b0000011001: data <= 8'h00; 
        10'b0000011010: data <= 8'h00; 
        10'b0000011011: data <= 8'h00; 
        10'b0000011100: data <= 8'h00; 
        10'b0000011101: data <= 8'h00; 
        10'b0000011110: data <= 8'h00; 
        10'b0000011111: data <= 8'h00; 
        10'b0000100000: data <= 8'h00; 
        10'b0000100001: data <= 8'h00; 
        10'b0000100010: data <= 8'h00; 
        10'b0000100011: data <= 8'h00; 
        10'b0000100100: data <= 8'h00; 
        10'b0000100101: data <= 8'h00; 
        10'b0000100110: data <= 8'h00; 
        10'b0000100111: data <= 8'h00; 
        10'b0000101000: data <= 8'h00; 
        10'b0000101001: data <= 8'h00; 
        10'b0000101010: data <= 8'h00; 
        10'b0000101011: data <= 8'h00; 
        10'b0000101100: data <= 8'h00; 
        10'b0000101101: data <= 8'h00; 
        10'b0000101110: data <= 8'h00; 
        10'b0000101111: data <= 8'h00; 
        10'b0000110000: data <= 8'h00; 
        10'b0000110001: data <= 8'h00; 
        10'b0000110010: data <= 8'h00; 
        10'b0000110011: data <= 8'h00; 
        10'b0000110100: data <= 8'h00; 
        10'b0000110101: data <= 8'h00; 
        10'b0000110110: data <= 8'h00; 
        10'b0000110111: data <= 8'h00; 
        10'b0000111000: data <= 8'h00; 
        10'b0000111001: data <= 8'h00; 
        10'b0000111010: data <= 8'h00; 
        10'b0000111011: data <= 8'h00; 
        10'b0000111100: data <= 8'h00; 
        10'b0000111101: data <= 8'h00; 
        10'b0000111110: data <= 8'h00; 
        10'b0000111111: data <= 8'h00; 
        10'b0001000000: data <= 8'h00; 
        10'b0001000001: data <= 8'h00; 
        10'b0001000010: data <= 8'h00; 
        10'b0001000011: data <= 8'h00; 
        10'b0001000100: data <= 8'h00; 
        10'b0001000101: data <= 8'h00; 
        10'b0001000110: data <= 8'h00; 
        10'b0001000111: data <= 8'h00; 
        10'b0001001000: data <= 8'h00; 
        10'b0001001001: data <= 8'h00; 
        10'b0001001010: data <= 8'h00; 
        10'b0001001011: data <= 8'h00; 
        10'b0001001100: data <= 8'h00; 
        10'b0001001101: data <= 8'h00; 
        10'b0001001110: data <= 8'h00; 
        10'b0001001111: data <= 8'h00; 
        10'b0001010000: data <= 8'h00; 
        10'b0001010001: data <= 8'h00; 
        10'b0001010010: data <= 8'h00; 
        10'b0001010011: data <= 8'h00; 
        10'b0001010100: data <= 8'h00; 
        10'b0001010101: data <= 8'h00; 
        10'b0001010110: data <= 8'h00; 
        10'b0001010111: data <= 8'h00; 
        10'b0001011000: data <= 8'h00; 
        10'b0001011001: data <= 8'h00; 
        10'b0001011010: data <= 8'h00; 
        10'b0001011011: data <= 8'h00; 
        10'b0001011100: data <= 8'h00; 
        10'b0001011101: data <= 8'h00; 
        10'b0001011110: data <= 8'h00; 
        10'b0001011111: data <= 8'h00; 
        10'b0001100000: data <= 8'h00; 
        10'b0001100001: data <= 8'h00; 
        10'b0001100010: data <= 8'h00; 
        10'b0001100011: data <= 8'h00; 
        10'b0001100100: data <= 8'h00; 
        10'b0001100101: data <= 8'h00; 
        10'b0001100110: data <= 8'h00; 
        10'b0001100111: data <= 8'h00; 
        10'b0001101000: data <= 8'h00; 
        10'b0001101001: data <= 8'h00; 
        10'b0001101010: data <= 8'h00; 
        10'b0001101011: data <= 8'h00; 
        10'b0001101100: data <= 8'h00; 
        10'b0001101101: data <= 8'h00; 
        10'b0001101110: data <= 8'h00; 
        10'b0001101111: data <= 8'h00; 
        10'b0001110000: data <= 8'h00; 
        10'b0001110001: data <= 8'h00; 
        10'b0001110010: data <= 8'h00; 
        10'b0001110011: data <= 8'h00; 
        10'b0001110100: data <= 8'h00; 
        10'b0001110101: data <= 8'h00; 
        10'b0001110110: data <= 8'h00; 
        10'b0001110111: data <= 8'h00; 
        10'b0001111000: data <= 8'hff; 
        10'b0001111001: data <= 8'hff; 
        10'b0001111010: data <= 8'hff; 
        10'b0001111011: data <= 8'hff; 
        10'b0001111100: data <= 8'hff; 
        10'b0001111101: data <= 8'hff; 
        10'b0001111110: data <= 8'hff; 
        10'b0001111111: data <= 8'h00; 
        10'b0010000000: data <= 8'h00; 
        10'b0010000001: data <= 8'h00; 
        10'b0010000010: data <= 8'h00; 
        10'b0010000011: data <= 8'h00; 
        10'b0010000100: data <= 8'h00; 
        10'b0010000101: data <= 8'h00; 
        10'b0010000110: data <= 8'h00; 
        10'b0010000111: data <= 8'h00; 
        10'b0010001000: data <= 8'h00; 
        10'b0010001001: data <= 8'h00; 
        10'b0010001010: data <= 8'h00; 
        10'b0010001011: data <= 8'h00; 
        10'b0010001100: data <= 8'h00; 
        10'b0010001101: data <= 8'h00; 
        10'b0010001110: data <= 8'h00; 
        10'b0010001111: data <= 8'h00; 
        10'b0010010000: data <= 8'h00; 
        10'b0010010001: data <= 8'h00; 
        10'b0010010010: data <= 8'hff; 
        10'b0010010011: data <= 8'hff; 
        10'b0010010100: data <= 8'h00; 
        10'b0010010101: data <= 8'h00; 
        10'b0010010110: data <= 8'h00; 
        10'b0010010111: data <= 8'h00; 
        10'b0010011000: data <= 8'h00; 
        10'b0010011001: data <= 8'h00; 
        10'b0010011010: data <= 8'h00; 
        10'b0010011011: data <= 8'h00; 
        10'b0010011100: data <= 8'h00; 
        10'b0010011101: data <= 8'h00; 
        10'b0010011110: data <= 8'h00; 
        10'b0010011111: data <= 8'h00; 
        10'b0010100000: data <= 8'h00; 
        10'b0010100001: data <= 8'h00; 
        10'b0010100010: data <= 8'h01; 
        10'b0010100011: data <= 8'h01; 
        10'b0010100100: data <= 8'h00; 
        10'b0010100101: data <= 8'h00; 
        10'b0010100110: data <= 8'h00; 
        10'b0010100111: data <= 8'h00; 
        10'b0010101000: data <= 8'h00; 
        10'b0010101001: data <= 8'h00; 
        10'b0010101010: data <= 8'h00; 
        10'b0010101011: data <= 8'h00; 
        10'b0010101100: data <= 8'h00; 
        10'b0010101101: data <= 8'hff; 
        10'b0010101110: data <= 8'h00; 
        10'b0010101111: data <= 8'h00; 
        10'b0010110000: data <= 8'h00; 
        10'b0010110001: data <= 8'h00; 
        10'b0010110010: data <= 8'h01; 
        10'b0010110011: data <= 8'h00; 
        10'b0010110100: data <= 8'h00; 
        10'b0010110101: data <= 8'h00; 
        10'b0010110110: data <= 8'h00; 
        10'b0010110111: data <= 8'h00; 
        10'b0010111000: data <= 8'h00; 
        10'b0010111001: data <= 8'h00; 
        10'b0010111010: data <= 8'h00; 
        10'b0010111011: data <= 8'h00; 
        10'b0010111100: data <= 8'h00; 
        10'b0010111101: data <= 8'h00; 
        10'b0010111110: data <= 8'h01; 
        10'b0010111111: data <= 8'h01; 
        10'b0011000000: data <= 8'h01; 
        10'b0011000001: data <= 8'h01; 
        10'b0011000010: data <= 8'h00; 
        10'b0011000011: data <= 8'h00; 
        10'b0011000100: data <= 8'h00; 
        10'b0011000101: data <= 8'h00; 
        10'b0011000110: data <= 8'h00; 
        10'b0011000111: data <= 8'h00; 
        10'b0011001000: data <= 8'hff; 
        10'b0011001001: data <= 8'hff; 
        10'b0011001010: data <= 8'hff; 
        10'b0011001011: data <= 8'h00; 
        10'b0011001100: data <= 8'h00; 
        10'b0011001101: data <= 8'h01; 
        10'b0011001110: data <= 8'h01; 
        10'b0011001111: data <= 8'h01; 
        10'b0011010000: data <= 8'h00; 
        10'b0011010001: data <= 8'h00; 
        10'b0011010010: data <= 8'h00; 
        10'b0011010011: data <= 8'h00; 
        10'b0011010100: data <= 8'h00; 
        10'b0011010101: data <= 8'h00; 
        10'b0011010110: data <= 8'h00; 
        10'b0011010111: data <= 8'h01; 
        10'b0011011000: data <= 8'h01; 
        10'b0011011001: data <= 8'h01; 
        10'b0011011010: data <= 8'h01; 
        10'b0011011011: data <= 8'h01; 
        10'b0011011100: data <= 8'h02; 
        10'b0011011101: data <= 8'h01; 
        10'b0011011110: data <= 8'h00; 
        10'b0011011111: data <= 8'h00; 
        10'b0011100000: data <= 8'h00; 
        10'b0011100001: data <= 8'h00; 
        10'b0011100010: data <= 8'h00; 
        10'b0011100011: data <= 8'h00; 
        10'b0011100100: data <= 8'hff; 
        10'b0011100101: data <= 8'hff; 
        10'b0011100110: data <= 8'hff; 
        10'b0011100111: data <= 8'h00; 
        10'b0011101000: data <= 8'h00; 
        10'b0011101001: data <= 8'h00; 
        10'b0011101010: data <= 8'h00; 
        10'b0011101011: data <= 8'h01; 
        10'b0011101100: data <= 8'h00; 
        10'b0011101101: data <= 8'h00; 
        10'b0011101110: data <= 8'hff; 
        10'b0011101111: data <= 8'h00; 
        10'b0011110000: data <= 8'h00; 
        10'b0011110001: data <= 8'h00; 
        10'b0011110010: data <= 8'h00; 
        10'b0011110011: data <= 8'h01; 
        10'b0011110100: data <= 8'h01; 
        10'b0011110101: data <= 8'h01; 
        10'b0011110110: data <= 8'h01; 
        10'b0011110111: data <= 8'h02; 
        10'b0011111000: data <= 8'h02; 
        10'b0011111001: data <= 8'h02; 
        10'b0011111010: data <= 8'h00; 
        10'b0011111011: data <= 8'h00; 
        10'b0011111100: data <= 8'h00; 
        10'b0011111101: data <= 8'h00; 
        10'b0011111110: data <= 8'h00; 
        10'b0011111111: data <= 8'h00; 
        10'b0100000000: data <= 8'hff; 
        10'b0100000001: data <= 8'hff; 
        10'b0100000010: data <= 8'h00; 
        10'b0100000011: data <= 8'h00; 
        10'b0100000100: data <= 8'h00; 
        10'b0100000101: data <= 8'h00; 
        10'b0100000110: data <= 8'h00; 
        10'b0100000111: data <= 8'h01; 
        10'b0100001000: data <= 8'h01; 
        10'b0100001001: data <= 8'h00; 
        10'b0100001010: data <= 8'hff; 
        10'b0100001011: data <= 8'hff; 
        10'b0100001100: data <= 8'hff; 
        10'b0100001101: data <= 8'hff; 
        10'b0100001110: data <= 8'h00; 
        10'b0100001111: data <= 8'h00; 
        10'b0100010000: data <= 8'h01; 
        10'b0100010001: data <= 8'h01; 
        10'b0100010010: data <= 8'h02; 
        10'b0100010011: data <= 8'h02; 
        10'b0100010100: data <= 8'h03; 
        10'b0100010101: data <= 8'h02; 
        10'b0100010110: data <= 8'h00; 
        10'b0100010111: data <= 8'h00; 
        10'b0100011000: data <= 8'h00; 
        10'b0100011001: data <= 8'h00; 
        10'b0100011010: data <= 8'h00; 
        10'b0100011011: data <= 8'h00; 
        10'b0100011100: data <= 8'h00; 
        10'b0100011101: data <= 8'h00; 
        10'b0100011110: data <= 8'h00; 
        10'b0100011111: data <= 8'h01; 
        10'b0100100000: data <= 8'h01; 
        10'b0100100001: data <= 8'h01; 
        10'b0100100010: data <= 8'h01; 
        10'b0100100011: data <= 8'h01; 
        10'b0100100100: data <= 8'h01; 
        10'b0100100101: data <= 8'h01; 
        10'b0100100110: data <= 8'h00; 
        10'b0100100111: data <= 8'hff; 
        10'b0100101000: data <= 8'hff; 
        10'b0100101001: data <= 8'hff; 
        10'b0100101010: data <= 8'hff; 
        10'b0100101011: data <= 8'hff; 
        10'b0100101100: data <= 8'hff; 
        10'b0100101101: data <= 8'h00; 
        10'b0100101110: data <= 8'h00; 
        10'b0100101111: data <= 8'h01; 
        10'b0100110000: data <= 8'h02; 
        10'b0100110001: data <= 8'h01; 
        10'b0100110010: data <= 8'h00; 
        10'b0100110011: data <= 8'h00; 
        10'b0100110100: data <= 8'h00; 
        10'b0100110101: data <= 8'h00; 
        10'b0100110110: data <= 8'h00; 
        10'b0100110111: data <= 8'h00; 
        10'b0100111000: data <= 8'h00; 
        10'b0100111001: data <= 8'h00; 
        10'b0100111010: data <= 8'h01; 
        10'b0100111011: data <= 8'h01; 
        10'b0100111100: data <= 8'h01; 
        10'b0100111101: data <= 8'h01; 
        10'b0100111110: data <= 8'h01; 
        10'b0100111111: data <= 8'h01; 
        10'b0101000000: data <= 8'h01; 
        10'b0101000001: data <= 8'h01; 
        10'b0101000010: data <= 8'h00; 
        10'b0101000011: data <= 8'hff; 
        10'b0101000100: data <= 8'hff; 
        10'b0101000101: data <= 8'hff; 
        10'b0101000110: data <= 8'hff; 
        10'b0101000111: data <= 8'hfe; 
        10'b0101001000: data <= 8'hfe; 
        10'b0101001001: data <= 8'hfe; 
        10'b0101001010: data <= 8'hfe; 
        10'b0101001011: data <= 8'hff; 
        10'b0101001100: data <= 8'h00; 
        10'b0101001101: data <= 8'h00; 
        10'b0101001110: data <= 8'h00; 
        10'b0101001111: data <= 8'h00; 
        10'b0101010000: data <= 8'h00; 
        10'b0101010001: data <= 8'h00; 
        10'b0101010010: data <= 8'h00; 
        10'b0101010011: data <= 8'h00; 
        10'b0101010100: data <= 8'h00; 
        10'b0101010101: data <= 8'h00; 
        10'b0101010110: data <= 8'h01; 
        10'b0101010111: data <= 8'h01; 
        10'b0101011000: data <= 8'h00; 
        10'b0101011001: data <= 8'h00; 
        10'b0101011010: data <= 8'h01; 
        10'b0101011011: data <= 8'h01; 
        10'b0101011100: data <= 8'h01; 
        10'b0101011101: data <= 8'h01; 
        10'b0101011110: data <= 8'h00; 
        10'b0101011111: data <= 8'hff; 
        10'b0101100000: data <= 8'hff; 
        10'b0101100001: data <= 8'hff; 
        10'b0101100010: data <= 8'hff; 
        10'b0101100011: data <= 8'hff; 
        10'b0101100100: data <= 8'hff; 
        10'b0101100101: data <= 8'hfe; 
        10'b0101100110: data <= 8'hfe; 
        10'b0101100111: data <= 8'hfe; 
        10'b0101101000: data <= 8'hff; 
        10'b0101101001: data <= 8'h00; 
        10'b0101101010: data <= 8'h00; 
        10'b0101101011: data <= 8'h00; 
        10'b0101101100: data <= 8'h00; 
        10'b0101101101: data <= 8'h00; 
        10'b0101101110: data <= 8'h00; 
        10'b0101101111: data <= 8'h00; 
        10'b0101110000: data <= 8'h00; 
        10'b0101110001: data <= 8'h00; 
        10'b0101110010: data <= 8'h00; 
        10'b0101110011: data <= 8'h00; 
        10'b0101110100: data <= 8'h00; 
        10'b0101110101: data <= 8'h00; 
        10'b0101110110: data <= 8'h01; 
        10'b0101110111: data <= 8'h01; 
        10'b0101111000: data <= 8'h01; 
        10'b0101111001: data <= 8'h01; 
        10'b0101111010: data <= 8'h00; 
        10'b0101111011: data <= 8'hff; 
        10'b0101111100: data <= 8'hff; 
        10'b0101111101: data <= 8'hff; 
        10'b0101111110: data <= 8'h00; 
        10'b0101111111: data <= 8'h00; 
        10'b0110000000: data <= 8'h00; 
        10'b0110000001: data <= 8'hff; 
        10'b0110000010: data <= 8'hff; 
        10'b0110000011: data <= 8'hff; 
        10'b0110000100: data <= 8'hff; 
        10'b0110000101: data <= 8'h00; 
        10'b0110000110: data <= 8'h00; 
        10'b0110000111: data <= 8'h00; 
        10'b0110001000: data <= 8'h00; 
        10'b0110001001: data <= 8'h00; 
        10'b0110001010: data <= 8'h00; 
        10'b0110001011: data <= 8'h00; 
        10'b0110001100: data <= 8'h00; 
        10'b0110001101: data <= 8'h00; 
        10'b0110001110: data <= 8'h00; 
        10'b0110001111: data <= 8'h00; 
        10'b0110010000: data <= 8'h00; 
        10'b0110010001: data <= 8'h01; 
        10'b0110010010: data <= 8'h01; 
        10'b0110010011: data <= 8'h00; 
        10'b0110010100: data <= 8'h00; 
        10'b0110010101: data <= 8'h00; 
        10'b0110010110: data <= 8'hff; 
        10'b0110010111: data <= 8'hff; 
        10'b0110011000: data <= 8'hff; 
        10'b0110011001: data <= 8'hff; 
        10'b0110011010: data <= 8'hff; 
        10'b0110011011: data <= 8'h00; 
        10'b0110011100: data <= 8'h00; 
        10'b0110011101: data <= 8'h00; 
        10'b0110011110: data <= 8'h00; 
        10'b0110011111: data <= 8'hff; 
        10'b0110100000: data <= 8'hff; 
        10'b0110100001: data <= 8'h00; 
        10'b0110100010: data <= 8'h00; 
        10'b0110100011: data <= 8'h00; 
        10'b0110100100: data <= 8'h00; 
        10'b0110100101: data <= 8'h00; 
        10'b0110100110: data <= 8'h00; 
        10'b0110100111: data <= 8'h00; 
        10'b0110101000: data <= 8'h00; 
        10'b0110101001: data <= 8'hff; 
        10'b0110101010: data <= 8'hff; 
        10'b0110101011: data <= 8'h00; 
        10'b0110101100: data <= 8'h00; 
        10'b0110101101: data <= 8'h01; 
        10'b0110101110: data <= 8'h00; 
        10'b0110101111: data <= 8'h00; 
        10'b0110110000: data <= 8'h00; 
        10'b0110110001: data <= 8'h00; 
        10'b0110110010: data <= 8'hff; 
        10'b0110110011: data <= 8'hff; 
        10'b0110110100: data <= 8'hff; 
        10'b0110110101: data <= 8'hff; 
        10'b0110110110: data <= 8'hff; 
        10'b0110110111: data <= 8'h00; 
        10'b0110111000: data <= 8'h00; 
        10'b0110111001: data <= 8'h00; 
        10'b0110111010: data <= 8'h00; 
        10'b0110111011: data <= 8'h00; 
        10'b0110111100: data <= 8'h00; 
        10'b0110111101: data <= 8'h00; 
        10'b0110111110: data <= 8'h00; 
        10'b0110111111: data <= 8'h00; 
        10'b0111000000: data <= 8'h00; 
        10'b0111000001: data <= 8'h00; 
        10'b0111000010: data <= 8'h00; 
        10'b0111000011: data <= 8'h00; 
        10'b0111000100: data <= 8'h00; 
        10'b0111000101: data <= 8'hff; 
        10'b0111000110: data <= 8'hff; 
        10'b0111000111: data <= 8'hff; 
        10'b0111001000: data <= 8'hff; 
        10'b0111001001: data <= 8'hff; 
        10'b0111001010: data <= 8'h00; 
        10'b0111001011: data <= 8'h00; 
        10'b0111001100: data <= 8'h00; 
        10'b0111001101: data <= 8'hff; 
        10'b0111001110: data <= 8'hff; 
        10'b0111001111: data <= 8'hff; 
        10'b0111010000: data <= 8'hff; 
        10'b0111010001: data <= 8'h00; 
        10'b0111010010: data <= 8'h00; 
        10'b0111010011: data <= 8'h00; 
        10'b0111010100: data <= 8'h00; 
        10'b0111010101: data <= 8'h00; 
        10'b0111010110: data <= 8'h00; 
        10'b0111010111: data <= 8'h00; 
        10'b0111011000: data <= 8'h00; 
        10'b0111011001: data <= 8'h00; 
        10'b0111011010: data <= 8'h00; 
        10'b0111011011: data <= 8'h00; 
        10'b0111011100: data <= 8'h00; 
        10'b0111011101: data <= 8'h00; 
        10'b0111011110: data <= 8'h00; 
        10'b0111011111: data <= 8'h00; 
        10'b0111100000: data <= 8'h00; 
        10'b0111100001: data <= 8'h00; 
        10'b0111100010: data <= 8'h00; 
        10'b0111100011: data <= 8'hff; 
        10'b0111100100: data <= 8'hfe; 
        10'b0111100101: data <= 8'hfe; 
        10'b0111100110: data <= 8'hff; 
        10'b0111100111: data <= 8'hff; 
        10'b0111101000: data <= 8'hff; 
        10'b0111101001: data <= 8'hff; 
        10'b0111101010: data <= 8'hff; 
        10'b0111101011: data <= 8'hff; 
        10'b0111101100: data <= 8'h00; 
        10'b0111101101: data <= 8'h00; 
        10'b0111101110: data <= 8'h01; 
        10'b0111101111: data <= 8'h00; 
        10'b0111110000: data <= 8'h00; 
        10'b0111110001: data <= 8'h00; 
        10'b0111110010: data <= 8'h00; 
        10'b0111110011: data <= 8'h00; 
        10'b0111110100: data <= 8'h00; 
        10'b0111110101: data <= 8'h00; 
        10'b0111110110: data <= 8'h00; 
        10'b0111110111: data <= 8'h00; 
        10'b0111111000: data <= 8'h00; 
        10'b0111111001: data <= 8'h00; 
        10'b0111111010: data <= 8'h00; 
        10'b0111111011: data <= 8'h00; 
        10'b0111111100: data <= 8'h00; 
        10'b0111111101: data <= 8'h00; 
        10'b0111111110: data <= 8'h01; 
        10'b0111111111: data <= 8'h00; 
        10'b1000000000: data <= 8'hff; 
        10'b1000000001: data <= 8'hff; 
        10'b1000000010: data <= 8'hfe; 
        10'b1000000011: data <= 8'hfe; 
        10'b1000000100: data <= 8'hff; 
        10'b1000000101: data <= 8'hff; 
        10'b1000000110: data <= 8'h00; 
        10'b1000000111: data <= 8'h00; 
        10'b1000001000: data <= 8'h00; 
        10'b1000001001: data <= 8'h00; 
        10'b1000001010: data <= 8'h00; 
        10'b1000001011: data <= 8'h00; 
        10'b1000001100: data <= 8'h00; 
        10'b1000001101: data <= 8'h00; 
        10'b1000001110: data <= 8'h00; 
        10'b1000001111: data <= 8'h00; 
        10'b1000010000: data <= 8'h00; 
        10'b1000010001: data <= 8'h00; 
        10'b1000010010: data <= 8'h00; 
        10'b1000010011: data <= 8'h00; 
        10'b1000010100: data <= 8'h00; 
        10'b1000010101: data <= 8'h00; 
        10'b1000010110: data <= 8'h00; 
        10'b1000010111: data <= 8'h00; 
        10'b1000011000: data <= 8'h00; 
        10'b1000011001: data <= 8'h01; 
        10'b1000011010: data <= 8'h01; 
        10'b1000011011: data <= 8'h01; 
        10'b1000011100: data <= 8'h00; 
        10'b1000011101: data <= 8'h00; 
        10'b1000011110: data <= 8'h00; 
        10'b1000011111: data <= 8'h00; 
        10'b1000100000: data <= 8'h00; 
        10'b1000100001: data <= 8'h00; 
        10'b1000100010: data <= 8'h00; 
        10'b1000100011: data <= 8'h00; 
        10'b1000100100: data <= 8'h00; 
        10'b1000100101: data <= 8'h00; 
        10'b1000100110: data <= 8'h00; 
        10'b1000100111: data <= 8'h00; 
        10'b1000101000: data <= 8'h00; 
        10'b1000101001: data <= 8'h00; 
        10'b1000101010: data <= 8'h01; 
        10'b1000101011: data <= 8'h00; 
        10'b1000101100: data <= 8'h00; 
        10'b1000101101: data <= 8'h00; 
        10'b1000101110: data <= 8'h00; 
        10'b1000101111: data <= 8'h00; 
        10'b1000110000: data <= 8'h00; 
        10'b1000110001: data <= 8'h00; 
        10'b1000110010: data <= 8'h00; 
        10'b1000110011: data <= 8'h00; 
        10'b1000110100: data <= 8'h00; 
        10'b1000110101: data <= 8'h01; 
        10'b1000110110: data <= 8'h01; 
        10'b1000110111: data <= 8'h01; 
        10'b1000111000: data <= 8'h01; 
        10'b1000111001: data <= 8'h01; 
        10'b1000111010: data <= 8'h01; 
        10'b1000111011: data <= 8'h01; 
        10'b1000111100: data <= 8'h01; 
        10'b1000111101: data <= 8'h01; 
        10'b1000111110: data <= 8'h00; 
        10'b1000111111: data <= 8'h00; 
        10'b1001000000: data <= 8'h00; 
        10'b1001000001: data <= 8'h00; 
        10'b1001000010: data <= 8'h00; 
        10'b1001000011: data <= 8'h00; 
        10'b1001000100: data <= 8'h00; 
        10'b1001000101: data <= 8'h00; 
        10'b1001000110: data <= 8'h01; 
        10'b1001000111: data <= 8'h01; 
        10'b1001001000: data <= 8'h00; 
        10'b1001001001: data <= 8'h00; 
        10'b1001001010: data <= 8'h00; 
        10'b1001001011: data <= 8'h00; 
        10'b1001001100: data <= 8'h00; 
        10'b1001001101: data <= 8'h00; 
        10'b1001001110: data <= 8'h00; 
        10'b1001001111: data <= 8'h00; 
        10'b1001010000: data <= 8'h00; 
        10'b1001010001: data <= 8'h00; 
        10'b1001010010: data <= 8'h00; 
        10'b1001010011: data <= 8'h01; 
        10'b1001010100: data <= 8'h01; 
        10'b1001010101: data <= 8'h01; 
        10'b1001010110: data <= 8'h01; 
        10'b1001010111: data <= 8'h00; 
        10'b1001011000: data <= 8'h00; 
        10'b1001011001: data <= 8'h00; 
        10'b1001011010: data <= 8'h00; 
        10'b1001011011: data <= 8'h00; 
        10'b1001011100: data <= 8'h00; 
        10'b1001011101: data <= 8'h00; 
        10'b1001011110: data <= 8'h00; 
        10'b1001011111: data <= 8'h00; 
        10'b1001100000: data <= 8'h00; 
        10'b1001100001: data <= 8'h01; 
        10'b1001100010: data <= 8'h01; 
        10'b1001100011: data <= 8'h00; 
        10'b1001100100: data <= 8'h00; 
        10'b1001100101: data <= 8'h00; 
        10'b1001100110: data <= 8'h00; 
        10'b1001100111: data <= 8'h00; 
        10'b1001101000: data <= 8'h00; 
        10'b1001101001: data <= 8'h00; 
        10'b1001101010: data <= 8'h00; 
        10'b1001101011: data <= 8'h00; 
        10'b1001101100: data <= 8'h00; 
        10'b1001101101: data <= 8'h00; 
        10'b1001101110: data <= 8'h00; 
        10'b1001101111: data <= 8'h00; 
        10'b1001110000: data <= 8'h00; 
        10'b1001110001: data <= 8'h01; 
        10'b1001110010: data <= 8'h00; 
        10'b1001110011: data <= 8'h01; 
        10'b1001110100: data <= 8'h01; 
        10'b1001110101: data <= 8'h01; 
        10'b1001110110: data <= 8'h01; 
        10'b1001110111: data <= 8'h00; 
        10'b1001111000: data <= 8'h00; 
        10'b1001111001: data <= 8'h00; 
        10'b1001111010: data <= 8'h00; 
        10'b1001111011: data <= 8'h00; 
        10'b1001111100: data <= 8'h00; 
        10'b1001111101: data <= 8'h00; 
        10'b1001111110: data <= 8'h00; 
        10'b1001111111: data <= 8'h00; 
        10'b1010000000: data <= 8'h00; 
        10'b1010000001: data <= 8'h00; 
        10'b1010000010: data <= 8'h00; 
        10'b1010000011: data <= 8'h00; 
        10'b1010000100: data <= 8'h00; 
        10'b1010000101: data <= 8'h00; 
        10'b1010000110: data <= 8'h00; 
        10'b1010000111: data <= 8'h00; 
        10'b1010001000: data <= 8'h00; 
        10'b1010001001: data <= 8'h00; 
        10'b1010001010: data <= 8'h00; 
        10'b1010001011: data <= 8'h00; 
        10'b1010001100: data <= 8'h00; 
        10'b1010001101: data <= 8'h00; 
        10'b1010001110: data <= 8'h00; 
        10'b1010001111: data <= 8'h01; 
        10'b1010010000: data <= 8'h01; 
        10'b1010010001: data <= 8'h00; 
        10'b1010010010: data <= 8'h00; 
        10'b1010010011: data <= 8'h00; 
        10'b1010010100: data <= 8'h00; 
        10'b1010010101: data <= 8'h00; 
        10'b1010010110: data <= 8'h00; 
        10'b1010010111: data <= 8'h00; 
        10'b1010011000: data <= 8'h00; 
        10'b1010011001: data <= 8'h00; 
        10'b1010011010: data <= 8'h00; 
        10'b1010011011: data <= 8'h00; 
        10'b1010011100: data <= 8'h00; 
        10'b1010011101: data <= 8'h00; 
        10'b1010011110: data <= 8'h00; 
        10'b1010011111: data <= 8'h00; 
        10'b1010100000: data <= 8'h00; 
        10'b1010100001: data <= 8'h00; 
        10'b1010100010: data <= 8'h00; 
        10'b1010100011: data <= 8'h00; 
        10'b1010100100: data <= 8'h00; 
        10'b1010100101: data <= 8'h00; 
        10'b1010100110: data <= 8'h00; 
        10'b1010100111: data <= 8'h00; 
        10'b1010101000: data <= 8'h00; 
        10'b1010101001: data <= 8'h00; 
        10'b1010101010: data <= 8'h01; 
        10'b1010101011: data <= 8'h00; 
        10'b1010101100: data <= 8'h00; 
        10'b1010101101: data <= 8'h00; 
        10'b1010101110: data <= 8'h01; 
        10'b1010101111: data <= 8'h01; 
        10'b1010110000: data <= 8'h00; 
        10'b1010110001: data <= 8'h00; 
        10'b1010110010: data <= 8'h00; 
        10'b1010110011: data <= 8'h00; 
        10'b1010110100: data <= 8'h00; 
        10'b1010110101: data <= 8'h00; 
        10'b1010110110: data <= 8'h00; 
        10'b1010110111: data <= 8'h00; 
        10'b1010111000: data <= 8'h00; 
        10'b1010111001: data <= 8'h00; 
        10'b1010111010: data <= 8'h00; 
        10'b1010111011: data <= 8'h00; 
        10'b1010111100: data <= 8'h00; 
        10'b1010111101: data <= 8'h00; 
        10'b1010111110: data <= 8'h00; 
        10'b1010111111: data <= 8'h00; 
        10'b1011000000: data <= 8'h00; 
        10'b1011000001: data <= 8'h00; 
        10'b1011000010: data <= 8'h00; 
        10'b1011000011: data <= 8'h00; 
        10'b1011000100: data <= 8'h00; 
        10'b1011000101: data <= 8'h00; 
        10'b1011000110: data <= 8'h00; 
        10'b1011000111: data <= 8'h00; 
        10'b1011001000: data <= 8'h00; 
        10'b1011001001: data <= 8'h00; 
        10'b1011001010: data <= 8'h00; 
        10'b1011001011: data <= 8'h00; 
        10'b1011001100: data <= 8'h00; 
        10'b1011001101: data <= 8'h00; 
        10'b1011001110: data <= 8'h00; 
        10'b1011001111: data <= 8'h00; 
        10'b1011010000: data <= 8'h00; 
        10'b1011010001: data <= 8'h00; 
        10'b1011010010: data <= 8'h00; 
        10'b1011010011: data <= 8'h00; 
        10'b1011010100: data <= 8'h00; 
        10'b1011010101: data <= 8'h00; 
        10'b1011010110: data <= 8'h00; 
        10'b1011010111: data <= 8'h00; 
        10'b1011011000: data <= 8'h00; 
        10'b1011011001: data <= 8'h00; 
        10'b1011011010: data <= 8'h00; 
        10'b1011011011: data <= 8'h00; 
        10'b1011011100: data <= 8'h00; 
        10'b1011011101: data <= 8'h00; 
        10'b1011011110: data <= 8'h00; 
        10'b1011011111: data <= 8'h00; 
        10'b1011100000: data <= 8'h00; 
        10'b1011100001: data <= 8'h00; 
        10'b1011100010: data <= 8'h00; 
        10'b1011100011: data <= 8'h00; 
        10'b1011100100: data <= 8'h00; 
        10'b1011100101: data <= 8'h00; 
        10'b1011100110: data <= 8'h00; 
        10'b1011100111: data <= 8'h00; 
        10'b1011101000: data <= 8'h00; 
        10'b1011101001: data <= 8'h00; 
        10'b1011101010: data <= 8'h00; 
        10'b1011101011: data <= 8'h00; 
        10'b1011101100: data <= 8'h00; 
        10'b1011101101: data <= 8'h00; 
        10'b1011101110: data <= 8'h00; 
        10'b1011101111: data <= 8'h00; 
        10'b1011110000: data <= 8'h00; 
        10'b1011110001: data <= 8'h00; 
        10'b1011110010: data <= 8'h00; 
        10'b1011110011: data <= 8'h00; 
        10'b1011110100: data <= 8'h00; 
        10'b1011110101: data <= 8'h00; 
        10'b1011110110: data <= 8'h00; 
        10'b1011110111: data <= 8'h00; 
        10'b1011111000: data <= 8'h00; 
        10'b1011111001: data <= 8'h00; 
        10'b1011111010: data <= 8'h00; 
        10'b1011111011: data <= 8'h00; 
        10'b1011111100: data <= 8'h00; 
        10'b1011111101: data <= 8'h00; 
        10'b1011111110: data <= 8'h00; 
        10'b1011111111: data <= 8'h00; 
        10'b1100000000: data <= 8'h00; 
        10'b1100000001: data <= 8'h00; 
        10'b1100000010: data <= 8'h00; 
        10'b1100000011: data <= 8'h00; 
        10'b1100000100: data <= 8'h00; 
        10'b1100000101: data <= 8'h00; 
        10'b1100000110: data <= 8'h00; 
        10'b1100000111: data <= 8'h00; 
        10'b1100001000: data <= 8'h00; 
        10'b1100001001: data <= 8'h00; 
        10'b1100001010: data <= 8'h00; 
        10'b1100001011: data <= 8'h00; 
        10'b1100001100: data <= 8'h00; 
        10'b1100001101: data <= 8'h00; 
        10'b1100001110: data <= 8'h00; 
        10'b1100001111: data <= 8'h00; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 3) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 9'h000; 
        10'b0000000001: data <= 9'h000; 
        10'b0000000010: data <= 9'h000; 
        10'b0000000011: data <= 9'h000; 
        10'b0000000100: data <= 9'h000; 
        10'b0000000101: data <= 9'h000; 
        10'b0000000110: data <= 9'h000; 
        10'b0000000111: data <= 9'h000; 
        10'b0000001000: data <= 9'h000; 
        10'b0000001001: data <= 9'h000; 
        10'b0000001010: data <= 9'h000; 
        10'b0000001011: data <= 9'h000; 
        10'b0000001100: data <= 9'h000; 
        10'b0000001101: data <= 9'h000; 
        10'b0000001110: data <= 9'h000; 
        10'b0000001111: data <= 9'h000; 
        10'b0000010000: data <= 9'h000; 
        10'b0000010001: data <= 9'h000; 
        10'b0000010010: data <= 9'h000; 
        10'b0000010011: data <= 9'h000; 
        10'b0000010100: data <= 9'h000; 
        10'b0000010101: data <= 9'h000; 
        10'b0000010110: data <= 9'h000; 
        10'b0000010111: data <= 9'h000; 
        10'b0000011000: data <= 9'h000; 
        10'b0000011001: data <= 9'h000; 
        10'b0000011010: data <= 9'h000; 
        10'b0000011011: data <= 9'h000; 
        10'b0000011100: data <= 9'h000; 
        10'b0000011101: data <= 9'h000; 
        10'b0000011110: data <= 9'h000; 
        10'b0000011111: data <= 9'h000; 
        10'b0000100000: data <= 9'h000; 
        10'b0000100001: data <= 9'h000; 
        10'b0000100010: data <= 9'h000; 
        10'b0000100011: data <= 9'h000; 
        10'b0000100100: data <= 9'h000; 
        10'b0000100101: data <= 9'h000; 
        10'b0000100110: data <= 9'h000; 
        10'b0000100111: data <= 9'h000; 
        10'b0000101000: data <= 9'h000; 
        10'b0000101001: data <= 9'h000; 
        10'b0000101010: data <= 9'h000; 
        10'b0000101011: data <= 9'h000; 
        10'b0000101100: data <= 9'h000; 
        10'b0000101101: data <= 9'h000; 
        10'b0000101110: data <= 9'h000; 
        10'b0000101111: data <= 9'h000; 
        10'b0000110000: data <= 9'h000; 
        10'b0000110001: data <= 9'h000; 
        10'b0000110010: data <= 9'h000; 
        10'b0000110011: data <= 9'h000; 
        10'b0000110100: data <= 9'h000; 
        10'b0000110101: data <= 9'h000; 
        10'b0000110110: data <= 9'h000; 
        10'b0000110111: data <= 9'h000; 
        10'b0000111000: data <= 9'h000; 
        10'b0000111001: data <= 9'h000; 
        10'b0000111010: data <= 9'h000; 
        10'b0000111011: data <= 9'h000; 
        10'b0000111100: data <= 9'h000; 
        10'b0000111101: data <= 9'h000; 
        10'b0000111110: data <= 9'h000; 
        10'b0000111111: data <= 9'h000; 
        10'b0001000000: data <= 9'h000; 
        10'b0001000001: data <= 9'h000; 
        10'b0001000010: data <= 9'h000; 
        10'b0001000011: data <= 9'h000; 
        10'b0001000100: data <= 9'h000; 
        10'b0001000101: data <= 9'h000; 
        10'b0001000110: data <= 9'h000; 
        10'b0001000111: data <= 9'h000; 
        10'b0001001000: data <= 9'h000; 
        10'b0001001001: data <= 9'h000; 
        10'b0001001010: data <= 9'h000; 
        10'b0001001011: data <= 9'h000; 
        10'b0001001100: data <= 9'h000; 
        10'b0001001101: data <= 9'h000; 
        10'b0001001110: data <= 9'h000; 
        10'b0001001111: data <= 9'h000; 
        10'b0001010000: data <= 9'h000; 
        10'b0001010001: data <= 9'h000; 
        10'b0001010010: data <= 9'h000; 
        10'b0001010011: data <= 9'h000; 
        10'b0001010100: data <= 9'h000; 
        10'b0001010101: data <= 9'h000; 
        10'b0001010110: data <= 9'h000; 
        10'b0001010111: data <= 9'h000; 
        10'b0001011000: data <= 9'h000; 
        10'b0001011001: data <= 9'h000; 
        10'b0001011010: data <= 9'h000; 
        10'b0001011011: data <= 9'h000; 
        10'b0001011100: data <= 9'h000; 
        10'b0001011101: data <= 9'h000; 
        10'b0001011110: data <= 9'h1ff; 
        10'b0001011111: data <= 9'h1ff; 
        10'b0001100000: data <= 9'h1ff; 
        10'b0001100001: data <= 9'h1ff; 
        10'b0001100010: data <= 9'h1ff; 
        10'b0001100011: data <= 9'h000; 
        10'b0001100100: data <= 9'h000; 
        10'b0001100101: data <= 9'h000; 
        10'b0001100110: data <= 9'h000; 
        10'b0001100111: data <= 9'h000; 
        10'b0001101000: data <= 9'h000; 
        10'b0001101001: data <= 9'h000; 
        10'b0001101010: data <= 9'h1ff; 
        10'b0001101011: data <= 9'h000; 
        10'b0001101100: data <= 9'h1ff; 
        10'b0001101101: data <= 9'h000; 
        10'b0001101110: data <= 9'h000; 
        10'b0001101111: data <= 9'h000; 
        10'b0001110000: data <= 9'h000; 
        10'b0001110001: data <= 9'h000; 
        10'b0001110010: data <= 9'h000; 
        10'b0001110011: data <= 9'h000; 
        10'b0001110100: data <= 9'h000; 
        10'b0001110101: data <= 9'h000; 
        10'b0001110110: data <= 9'h000; 
        10'b0001110111: data <= 9'h1ff; 
        10'b0001111000: data <= 9'h1ff; 
        10'b0001111001: data <= 9'h1fe; 
        10'b0001111010: data <= 9'h1fe; 
        10'b0001111011: data <= 9'h1ff; 
        10'b0001111100: data <= 9'h1ff; 
        10'b0001111101: data <= 9'h1fe; 
        10'b0001111110: data <= 9'h1ff; 
        10'b0001111111: data <= 9'h000; 
        10'b0010000000: data <= 9'h000; 
        10'b0010000001: data <= 9'h000; 
        10'b0010000010: data <= 9'h000; 
        10'b0010000011: data <= 9'h1ff; 
        10'b0010000100: data <= 9'h1ff; 
        10'b0010000101: data <= 9'h000; 
        10'b0010000110: data <= 9'h000; 
        10'b0010000111: data <= 9'h000; 
        10'b0010001000: data <= 9'h000; 
        10'b0010001001: data <= 9'h000; 
        10'b0010001010: data <= 9'h000; 
        10'b0010001011: data <= 9'h000; 
        10'b0010001100: data <= 9'h000; 
        10'b0010001101: data <= 9'h000; 
        10'b0010001110: data <= 9'h000; 
        10'b0010001111: data <= 9'h000; 
        10'b0010010000: data <= 9'h000; 
        10'b0010010001: data <= 9'h1ff; 
        10'b0010010010: data <= 9'h1ff; 
        10'b0010010011: data <= 9'h1ff; 
        10'b0010010100: data <= 9'h1ff; 
        10'b0010010101: data <= 9'h000; 
        10'b0010010110: data <= 9'h000; 
        10'b0010010111: data <= 9'h000; 
        10'b0010011000: data <= 9'h000; 
        10'b0010011001: data <= 9'h1ff; 
        10'b0010011010: data <= 9'h000; 
        10'b0010011011: data <= 9'h000; 
        10'b0010011100: data <= 9'h001; 
        10'b0010011101: data <= 9'h001; 
        10'b0010011110: data <= 9'h001; 
        10'b0010011111: data <= 9'h001; 
        10'b0010100000: data <= 9'h001; 
        10'b0010100001: data <= 9'h001; 
        10'b0010100010: data <= 9'h001; 
        10'b0010100011: data <= 9'h001; 
        10'b0010100100: data <= 9'h001; 
        10'b0010100101: data <= 9'h000; 
        10'b0010100110: data <= 9'h000; 
        10'b0010100111: data <= 9'h000; 
        10'b0010101000: data <= 9'h000; 
        10'b0010101001: data <= 9'h000; 
        10'b0010101010: data <= 9'h000; 
        10'b0010101011: data <= 9'h000; 
        10'b0010101100: data <= 9'h1ff; 
        10'b0010101101: data <= 9'h1ff; 
        10'b0010101110: data <= 9'h1ff; 
        10'b0010101111: data <= 9'h000; 
        10'b0010110000: data <= 9'h000; 
        10'b0010110001: data <= 9'h000; 
        10'b0010110010: data <= 9'h001; 
        10'b0010110011: data <= 9'h001; 
        10'b0010110100: data <= 9'h000; 
        10'b0010110101: data <= 9'h000; 
        10'b0010110110: data <= 9'h000; 
        10'b0010110111: data <= 9'h000; 
        10'b0010111000: data <= 9'h000; 
        10'b0010111001: data <= 9'h000; 
        10'b0010111010: data <= 9'h000; 
        10'b0010111011: data <= 9'h001; 
        10'b0010111100: data <= 9'h001; 
        10'b0010111101: data <= 9'h001; 
        10'b0010111110: data <= 9'h002; 
        10'b0010111111: data <= 9'h002; 
        10'b0011000000: data <= 9'h003; 
        10'b0011000001: data <= 9'h001; 
        10'b0011000010: data <= 9'h001; 
        10'b0011000011: data <= 9'h000; 
        10'b0011000100: data <= 9'h000; 
        10'b0011000101: data <= 9'h000; 
        10'b0011000110: data <= 9'h000; 
        10'b0011000111: data <= 9'h1ff; 
        10'b0011001000: data <= 9'h1ff; 
        10'b0011001001: data <= 9'h1fe; 
        10'b0011001010: data <= 9'h1ff; 
        10'b0011001011: data <= 9'h000; 
        10'b0011001100: data <= 9'h001; 
        10'b0011001101: data <= 9'h001; 
        10'b0011001110: data <= 9'h001; 
        10'b0011001111: data <= 9'h001; 
        10'b0011010000: data <= 9'h000; 
        10'b0011010001: data <= 9'h000; 
        10'b0011010010: data <= 9'h000; 
        10'b0011010011: data <= 9'h000; 
        10'b0011010100: data <= 9'h001; 
        10'b0011010101: data <= 9'h000; 
        10'b0011010110: data <= 9'h001; 
        10'b0011010111: data <= 9'h001; 
        10'b0011011000: data <= 9'h001; 
        10'b0011011001: data <= 9'h001; 
        10'b0011011010: data <= 9'h002; 
        10'b0011011011: data <= 9'h003; 
        10'b0011011100: data <= 9'h003; 
        10'b0011011101: data <= 9'h002; 
        10'b0011011110: data <= 9'h000; 
        10'b0011011111: data <= 9'h000; 
        10'b0011100000: data <= 9'h000; 
        10'b0011100001: data <= 9'h000; 
        10'b0011100010: data <= 9'h000; 
        10'b0011100011: data <= 9'h1ff; 
        10'b0011100100: data <= 9'h1fe; 
        10'b0011100101: data <= 9'h1fe; 
        10'b0011100110: data <= 9'h1ff; 
        10'b0011100111: data <= 9'h000; 
        10'b0011101000: data <= 9'h001; 
        10'b0011101001: data <= 9'h000; 
        10'b0011101010: data <= 9'h001; 
        10'b0011101011: data <= 9'h001; 
        10'b0011101100: data <= 9'h001; 
        10'b0011101101: data <= 9'h1ff; 
        10'b0011101110: data <= 9'h1fe; 
        10'b0011101111: data <= 9'h1ff; 
        10'b0011110000: data <= 9'h1ff; 
        10'b0011110001: data <= 9'h000; 
        10'b0011110010: data <= 9'h000; 
        10'b0011110011: data <= 9'h001; 
        10'b0011110100: data <= 9'h001; 
        10'b0011110101: data <= 9'h002; 
        10'b0011110110: data <= 9'h003; 
        10'b0011110111: data <= 9'h004; 
        10'b0011111000: data <= 9'h005; 
        10'b0011111001: data <= 9'h003; 
        10'b0011111010: data <= 9'h001; 
        10'b0011111011: data <= 9'h000; 
        10'b0011111100: data <= 9'h000; 
        10'b0011111101: data <= 9'h000; 
        10'b0011111110: data <= 9'h000; 
        10'b0011111111: data <= 9'h1ff; 
        10'b0100000000: data <= 9'h1ff; 
        10'b0100000001: data <= 9'h1ff; 
        10'b0100000010: data <= 9'h000; 
        10'b0100000011: data <= 9'h000; 
        10'b0100000100: data <= 9'h001; 
        10'b0100000101: data <= 9'h001; 
        10'b0100000110: data <= 9'h001; 
        10'b0100000111: data <= 9'h002; 
        10'b0100001000: data <= 9'h001; 
        10'b0100001001: data <= 9'h1ff; 
        10'b0100001010: data <= 9'h1fe; 
        10'b0100001011: data <= 9'h1fd; 
        10'b0100001100: data <= 9'h1fe; 
        10'b0100001101: data <= 9'h1ff; 
        10'b0100001110: data <= 9'h000; 
        10'b0100001111: data <= 9'h000; 
        10'b0100010000: data <= 9'h001; 
        10'b0100010001: data <= 9'h002; 
        10'b0100010010: data <= 9'h004; 
        10'b0100010011: data <= 9'h005; 
        10'b0100010100: data <= 9'h006; 
        10'b0100010101: data <= 9'h004; 
        10'b0100010110: data <= 9'h001; 
        10'b0100010111: data <= 9'h000; 
        10'b0100011000: data <= 9'h000; 
        10'b0100011001: data <= 9'h000; 
        10'b0100011010: data <= 9'h000; 
        10'b0100011011: data <= 9'h000; 
        10'b0100011100: data <= 9'h000; 
        10'b0100011101: data <= 9'h000; 
        10'b0100011110: data <= 9'h001; 
        10'b0100011111: data <= 9'h001; 
        10'b0100100000: data <= 9'h002; 
        10'b0100100001: data <= 9'h002; 
        10'b0100100010: data <= 9'h002; 
        10'b0100100011: data <= 9'h003; 
        10'b0100100100: data <= 9'h002; 
        10'b0100100101: data <= 9'h002; 
        10'b0100100110: data <= 9'h000; 
        10'b0100100111: data <= 9'h1ff; 
        10'b0100101000: data <= 9'h1fe; 
        10'b0100101001: data <= 9'h1fe; 
        10'b0100101010: data <= 9'h1fe; 
        10'b0100101011: data <= 9'h1fd; 
        10'b0100101100: data <= 9'h1fe; 
        10'b0100101101: data <= 9'h1ff; 
        10'b0100101110: data <= 9'h000; 
        10'b0100101111: data <= 9'h002; 
        10'b0100110000: data <= 9'h003; 
        10'b0100110001: data <= 9'h002; 
        10'b0100110010: data <= 9'h001; 
        10'b0100110011: data <= 9'h000; 
        10'b0100110100: data <= 9'h000; 
        10'b0100110101: data <= 9'h000; 
        10'b0100110110: data <= 9'h000; 
        10'b0100110111: data <= 9'h000; 
        10'b0100111000: data <= 9'h000; 
        10'b0100111001: data <= 9'h000; 
        10'b0100111010: data <= 9'h001; 
        10'b0100111011: data <= 9'h001; 
        10'b0100111100: data <= 9'h002; 
        10'b0100111101: data <= 9'h002; 
        10'b0100111110: data <= 9'h001; 
        10'b0100111111: data <= 9'h001; 
        10'b0101000000: data <= 9'h002; 
        10'b0101000001: data <= 9'h002; 
        10'b0101000010: data <= 9'h000; 
        10'b0101000011: data <= 9'h1ff; 
        10'b0101000100: data <= 9'h1fe; 
        10'b0101000101: data <= 9'h1fe; 
        10'b0101000110: data <= 9'h1fe; 
        10'b0101000111: data <= 9'h1fd; 
        10'b0101001000: data <= 9'h1fb; 
        10'b0101001001: data <= 9'h1fb; 
        10'b0101001010: data <= 9'h1fc; 
        10'b0101001011: data <= 9'h1fd; 
        10'b0101001100: data <= 9'h1ff; 
        10'b0101001101: data <= 9'h000; 
        10'b0101001110: data <= 9'h000; 
        10'b0101001111: data <= 9'h000; 
        10'b0101010000: data <= 9'h000; 
        10'b0101010001: data <= 9'h000; 
        10'b0101010010: data <= 9'h000; 
        10'b0101010011: data <= 9'h000; 
        10'b0101010100: data <= 9'h000; 
        10'b0101010101: data <= 9'h001; 
        10'b0101010110: data <= 9'h001; 
        10'b0101010111: data <= 9'h001; 
        10'b0101011000: data <= 9'h001; 
        10'b0101011001: data <= 9'h000; 
        10'b0101011010: data <= 9'h001; 
        10'b0101011011: data <= 9'h003; 
        10'b0101011100: data <= 9'h003; 
        10'b0101011101: data <= 9'h003; 
        10'b0101011110: data <= 9'h000; 
        10'b0101011111: data <= 9'h1ff; 
        10'b0101100000: data <= 9'h1fd; 
        10'b0101100001: data <= 9'h1fe; 
        10'b0101100010: data <= 9'h1ff; 
        10'b0101100011: data <= 9'h1fe; 
        10'b0101100100: data <= 9'h1fe; 
        10'b0101100101: data <= 9'h1fc; 
        10'b0101100110: data <= 9'h1fc; 
        10'b0101100111: data <= 9'h1fc; 
        10'b0101101000: data <= 9'h1fd; 
        10'b0101101001: data <= 9'h1ff; 
        10'b0101101010: data <= 9'h000; 
        10'b0101101011: data <= 9'h000; 
        10'b0101101100: data <= 9'h000; 
        10'b0101101101: data <= 9'h000; 
        10'b0101101110: data <= 9'h000; 
        10'b0101101111: data <= 9'h000; 
        10'b0101110000: data <= 9'h000; 
        10'b0101110001: data <= 9'h000; 
        10'b0101110010: data <= 9'h001; 
        10'b0101110011: data <= 9'h001; 
        10'b0101110100: data <= 9'h001; 
        10'b0101110101: data <= 9'h001; 
        10'b0101110110: data <= 9'h002; 
        10'b0101110111: data <= 9'h002; 
        10'b0101111000: data <= 9'h002; 
        10'b0101111001: data <= 9'h001; 
        10'b0101111010: data <= 9'h000; 
        10'b0101111011: data <= 9'h1fe; 
        10'b0101111100: data <= 9'h1fd; 
        10'b0101111101: data <= 9'h1ff; 
        10'b0101111110: data <= 9'h000; 
        10'b0101111111: data <= 9'h1ff; 
        10'b0110000000: data <= 9'h000; 
        10'b0110000001: data <= 9'h1ff; 
        10'b0110000010: data <= 9'h1fe; 
        10'b0110000011: data <= 9'h1fd; 
        10'b0110000100: data <= 9'h1fe; 
        10'b0110000101: data <= 9'h000; 
        10'b0110000110: data <= 9'h000; 
        10'b0110000111: data <= 9'h000; 
        10'b0110001000: data <= 9'h000; 
        10'b0110001001: data <= 9'h000; 
        10'b0110001010: data <= 9'h000; 
        10'b0110001011: data <= 9'h000; 
        10'b0110001100: data <= 9'h000; 
        10'b0110001101: data <= 9'h000; 
        10'b0110001110: data <= 9'h000; 
        10'b0110001111: data <= 9'h000; 
        10'b0110010000: data <= 9'h001; 
        10'b0110010001: data <= 9'h001; 
        10'b0110010010: data <= 9'h002; 
        10'b0110010011: data <= 9'h000; 
        10'b0110010100: data <= 9'h001; 
        10'b0110010101: data <= 9'h000; 
        10'b0110010110: data <= 9'h1ff; 
        10'b0110010111: data <= 9'h1ff; 
        10'b0110011000: data <= 9'h1fe; 
        10'b0110011001: data <= 9'h1fe; 
        10'b0110011010: data <= 9'h1fe; 
        10'b0110011011: data <= 9'h1ff; 
        10'b0110011100: data <= 9'h1ff; 
        10'b0110011101: data <= 9'h1ff; 
        10'b0110011110: data <= 9'h000; 
        10'b0110011111: data <= 9'h1fe; 
        10'b0110100000: data <= 9'h1ff; 
        10'b0110100001: data <= 9'h1ff; 
        10'b0110100010: data <= 9'h000; 
        10'b0110100011: data <= 9'h000; 
        10'b0110100100: data <= 9'h000; 
        10'b0110100101: data <= 9'h000; 
        10'b0110100110: data <= 9'h000; 
        10'b0110100111: data <= 9'h000; 
        10'b0110101000: data <= 9'h1ff; 
        10'b0110101001: data <= 9'h1ff; 
        10'b0110101010: data <= 9'h1ff; 
        10'b0110101011: data <= 9'h1ff; 
        10'b0110101100: data <= 9'h000; 
        10'b0110101101: data <= 9'h002; 
        10'b0110101110: data <= 9'h001; 
        10'b0110101111: data <= 9'h001; 
        10'b0110110000: data <= 9'h001; 
        10'b0110110001: data <= 9'h1ff; 
        10'b0110110010: data <= 9'h1fe; 
        10'b0110110011: data <= 9'h1fe; 
        10'b0110110100: data <= 9'h1fe; 
        10'b0110110101: data <= 9'h1fe; 
        10'b0110110110: data <= 9'h1ff; 
        10'b0110110111: data <= 9'h000; 
        10'b0110111000: data <= 9'h000; 
        10'b0110111001: data <= 9'h000; 
        10'b0110111010: data <= 9'h000; 
        10'b0110111011: data <= 9'h1ff; 
        10'b0110111100: data <= 9'h000; 
        10'b0110111101: data <= 9'h000; 
        10'b0110111110: data <= 9'h000; 
        10'b0110111111: data <= 9'h000; 
        10'b0111000000: data <= 9'h000; 
        10'b0111000001: data <= 9'h000; 
        10'b0111000010: data <= 9'h000; 
        10'b0111000011: data <= 9'h000; 
        10'b0111000100: data <= 9'h000; 
        10'b0111000101: data <= 9'h1ff; 
        10'b0111000110: data <= 9'h1fe; 
        10'b0111000111: data <= 9'h1fd; 
        10'b0111001000: data <= 9'h1fe; 
        10'b0111001001: data <= 9'h1ff; 
        10'b0111001010: data <= 9'h000; 
        10'b0111001011: data <= 9'h1ff; 
        10'b0111001100: data <= 9'h000; 
        10'b0111001101: data <= 9'h1ff; 
        10'b0111001110: data <= 9'h1fe; 
        10'b0111001111: data <= 9'h1fe; 
        10'b0111010000: data <= 9'h1ff; 
        10'b0111010001: data <= 9'h1ff; 
        10'b0111010010: data <= 9'h000; 
        10'b0111010011: data <= 9'h000; 
        10'b0111010100: data <= 9'h000; 
        10'b0111010101: data <= 9'h000; 
        10'b0111010110: data <= 9'h000; 
        10'b0111010111: data <= 9'h000; 
        10'b0111011000: data <= 9'h000; 
        10'b0111011001: data <= 9'h000; 
        10'b0111011010: data <= 9'h000; 
        10'b0111011011: data <= 9'h000; 
        10'b0111011100: data <= 9'h000; 
        10'b0111011101: data <= 9'h000; 
        10'b0111011110: data <= 9'h000; 
        10'b0111011111: data <= 9'h000; 
        10'b0111100000: data <= 9'h000; 
        10'b0111100001: data <= 9'h000; 
        10'b0111100010: data <= 9'h000; 
        10'b0111100011: data <= 9'h1fe; 
        10'b0111100100: data <= 9'h1fd; 
        10'b0111100101: data <= 9'h1fd; 
        10'b0111100110: data <= 9'h1fe; 
        10'b0111100111: data <= 9'h1ff; 
        10'b0111101000: data <= 9'h1fe; 
        10'b0111101001: data <= 9'h1fd; 
        10'b0111101010: data <= 9'h1fd; 
        10'b0111101011: data <= 9'h1ff; 
        10'b0111101100: data <= 9'h1ff; 
        10'b0111101101: data <= 9'h001; 
        10'b0111101110: data <= 9'h001; 
        10'b0111101111: data <= 9'h001; 
        10'b0111110000: data <= 9'h001; 
        10'b0111110001: data <= 9'h000; 
        10'b0111110010: data <= 9'h000; 
        10'b0111110011: data <= 9'h000; 
        10'b0111110100: data <= 9'h000; 
        10'b0111110101: data <= 9'h000; 
        10'b0111110110: data <= 9'h000; 
        10'b0111110111: data <= 9'h000; 
        10'b0111111000: data <= 9'h000; 
        10'b0111111001: data <= 9'h000; 
        10'b0111111010: data <= 9'h000; 
        10'b0111111011: data <= 9'h000; 
        10'b0111111100: data <= 9'h001; 
        10'b0111111101: data <= 9'h001; 
        10'b0111111110: data <= 9'h002; 
        10'b0111111111: data <= 9'h000; 
        10'b1000000000: data <= 9'h1fe; 
        10'b1000000001: data <= 9'h1fd; 
        10'b1000000010: data <= 9'h1fc; 
        10'b1000000011: data <= 9'h1fd; 
        10'b1000000100: data <= 9'h1fe; 
        10'b1000000101: data <= 9'h1ff; 
        10'b1000000110: data <= 9'h1ff; 
        10'b1000000111: data <= 9'h000; 
        10'b1000001000: data <= 9'h000; 
        10'b1000001001: data <= 9'h001; 
        10'b1000001010: data <= 9'h000; 
        10'b1000001011: data <= 9'h001; 
        10'b1000001100: data <= 9'h001; 
        10'b1000001101: data <= 9'h001; 
        10'b1000001110: data <= 9'h001; 
        10'b1000001111: data <= 9'h001; 
        10'b1000010000: data <= 9'h000; 
        10'b1000010001: data <= 9'h000; 
        10'b1000010010: data <= 9'h000; 
        10'b1000010011: data <= 9'h000; 
        10'b1000010100: data <= 9'h000; 
        10'b1000010101: data <= 9'h000; 
        10'b1000010110: data <= 9'h000; 
        10'b1000010111: data <= 9'h000; 
        10'b1000011000: data <= 9'h001; 
        10'b1000011001: data <= 9'h002; 
        10'b1000011010: data <= 9'h002; 
        10'b1000011011: data <= 9'h002; 
        10'b1000011100: data <= 9'h001; 
        10'b1000011101: data <= 9'h000; 
        10'b1000011110: data <= 9'h1ff; 
        10'b1000011111: data <= 9'h1ff; 
        10'b1000100000: data <= 9'h000; 
        10'b1000100001: data <= 9'h001; 
        10'b1000100010: data <= 9'h000; 
        10'b1000100011: data <= 9'h000; 
        10'b1000100100: data <= 9'h000; 
        10'b1000100101: data <= 9'h000; 
        10'b1000100110: data <= 9'h000; 
        10'b1000100111: data <= 9'h000; 
        10'b1000101000: data <= 9'h000; 
        10'b1000101001: data <= 9'h001; 
        10'b1000101010: data <= 9'h001; 
        10'b1000101011: data <= 9'h001; 
        10'b1000101100: data <= 9'h000; 
        10'b1000101101: data <= 9'h000; 
        10'b1000101110: data <= 9'h000; 
        10'b1000101111: data <= 9'h000; 
        10'b1000110000: data <= 9'h000; 
        10'b1000110001: data <= 9'h000; 
        10'b1000110010: data <= 9'h000; 
        10'b1000110011: data <= 9'h000; 
        10'b1000110100: data <= 9'h000; 
        10'b1000110101: data <= 9'h001; 
        10'b1000110110: data <= 9'h001; 
        10'b1000110111: data <= 9'h002; 
        10'b1000111000: data <= 9'h002; 
        10'b1000111001: data <= 9'h002; 
        10'b1000111010: data <= 9'h002; 
        10'b1000111011: data <= 9'h002; 
        10'b1000111100: data <= 9'h001; 
        10'b1000111101: data <= 9'h001; 
        10'b1000111110: data <= 9'h000; 
        10'b1000111111: data <= 9'h000; 
        10'b1001000000: data <= 9'h001; 
        10'b1001000001: data <= 9'h000; 
        10'b1001000010: data <= 9'h001; 
        10'b1001000011: data <= 9'h001; 
        10'b1001000100: data <= 9'h001; 
        10'b1001000101: data <= 9'h001; 
        10'b1001000110: data <= 9'h001; 
        10'b1001000111: data <= 9'h001; 
        10'b1001001000: data <= 9'h000; 
        10'b1001001001: data <= 9'h000; 
        10'b1001001010: data <= 9'h000; 
        10'b1001001011: data <= 9'h000; 
        10'b1001001100: data <= 9'h000; 
        10'b1001001101: data <= 9'h000; 
        10'b1001001110: data <= 9'h000; 
        10'b1001001111: data <= 9'h000; 
        10'b1001010000: data <= 9'h000; 
        10'b1001010001: data <= 9'h000; 
        10'b1001010010: data <= 9'h001; 
        10'b1001010011: data <= 9'h001; 
        10'b1001010100: data <= 9'h002; 
        10'b1001010101: data <= 9'h001; 
        10'b1001010110: data <= 9'h001; 
        10'b1001010111: data <= 9'h001; 
        10'b1001011000: data <= 9'h001; 
        10'b1001011001: data <= 9'h000; 
        10'b1001011010: data <= 9'h001; 
        10'b1001011011: data <= 9'h001; 
        10'b1001011100: data <= 9'h000; 
        10'b1001011101: data <= 9'h001; 
        10'b1001011110: data <= 9'h000; 
        10'b1001011111: data <= 9'h001; 
        10'b1001100000: data <= 9'h001; 
        10'b1001100001: data <= 9'h001; 
        10'b1001100010: data <= 9'h002; 
        10'b1001100011: data <= 9'h000; 
        10'b1001100100: data <= 9'h000; 
        10'b1001100101: data <= 9'h000; 
        10'b1001100110: data <= 9'h000; 
        10'b1001100111: data <= 9'h000; 
        10'b1001101000: data <= 9'h000; 
        10'b1001101001: data <= 9'h000; 
        10'b1001101010: data <= 9'h000; 
        10'b1001101011: data <= 9'h000; 
        10'b1001101100: data <= 9'h000; 
        10'b1001101101: data <= 9'h000; 
        10'b1001101110: data <= 9'h000; 
        10'b1001101111: data <= 9'h000; 
        10'b1001110000: data <= 9'h001; 
        10'b1001110001: data <= 9'h001; 
        10'b1001110010: data <= 9'h000; 
        10'b1001110011: data <= 9'h001; 
        10'b1001110100: data <= 9'h002; 
        10'b1001110101: data <= 9'h002; 
        10'b1001110110: data <= 9'h001; 
        10'b1001110111: data <= 9'h000; 
        10'b1001111000: data <= 9'h000; 
        10'b1001111001: data <= 9'h000; 
        10'b1001111010: data <= 9'h001; 
        10'b1001111011: data <= 9'h001; 
        10'b1001111100: data <= 9'h001; 
        10'b1001111101: data <= 9'h001; 
        10'b1001111110: data <= 9'h001; 
        10'b1001111111: data <= 9'h000; 
        10'b1010000000: data <= 9'h000; 
        10'b1010000001: data <= 9'h000; 
        10'b1010000010: data <= 9'h000; 
        10'b1010000011: data <= 9'h000; 
        10'b1010000100: data <= 9'h000; 
        10'b1010000101: data <= 9'h000; 
        10'b1010000110: data <= 9'h000; 
        10'b1010000111: data <= 9'h000; 
        10'b1010001000: data <= 9'h000; 
        10'b1010001001: data <= 9'h000; 
        10'b1010001010: data <= 9'h1ff; 
        10'b1010001011: data <= 9'h000; 
        10'b1010001100: data <= 9'h001; 
        10'b1010001101: data <= 9'h001; 
        10'b1010001110: data <= 9'h001; 
        10'b1010001111: data <= 9'h001; 
        10'b1010010000: data <= 9'h001; 
        10'b1010010001: data <= 9'h001; 
        10'b1010010010: data <= 9'h001; 
        10'b1010010011: data <= 9'h001; 
        10'b1010010100: data <= 9'h001; 
        10'b1010010101: data <= 9'h000; 
        10'b1010010110: data <= 9'h000; 
        10'b1010010111: data <= 9'h000; 
        10'b1010011000: data <= 9'h000; 
        10'b1010011001: data <= 9'h000; 
        10'b1010011010: data <= 9'h000; 
        10'b1010011011: data <= 9'h000; 
        10'b1010011100: data <= 9'h000; 
        10'b1010011101: data <= 9'h000; 
        10'b1010011110: data <= 9'h000; 
        10'b1010011111: data <= 9'h000; 
        10'b1010100000: data <= 9'h000; 
        10'b1010100001: data <= 9'h000; 
        10'b1010100010: data <= 9'h000; 
        10'b1010100011: data <= 9'h000; 
        10'b1010100100: data <= 9'h000; 
        10'b1010100101: data <= 9'h1ff; 
        10'b1010100110: data <= 9'h000; 
        10'b1010100111: data <= 9'h000; 
        10'b1010101000: data <= 9'h000; 
        10'b1010101001: data <= 9'h001; 
        10'b1010101010: data <= 9'h001; 
        10'b1010101011: data <= 9'h001; 
        10'b1010101100: data <= 9'h001; 
        10'b1010101101: data <= 9'h001; 
        10'b1010101110: data <= 9'h001; 
        10'b1010101111: data <= 9'h001; 
        10'b1010110000: data <= 9'h001; 
        10'b1010110001: data <= 9'h000; 
        10'b1010110010: data <= 9'h001; 
        10'b1010110011: data <= 9'h000; 
        10'b1010110100: data <= 9'h000; 
        10'b1010110101: data <= 9'h000; 
        10'b1010110110: data <= 9'h000; 
        10'b1010110111: data <= 9'h000; 
        10'b1010111000: data <= 9'h000; 
        10'b1010111001: data <= 9'h000; 
        10'b1010111010: data <= 9'h000; 
        10'b1010111011: data <= 9'h000; 
        10'b1010111100: data <= 9'h000; 
        10'b1010111101: data <= 9'h000; 
        10'b1010111110: data <= 9'h000; 
        10'b1010111111: data <= 9'h000; 
        10'b1011000000: data <= 9'h000; 
        10'b1011000001: data <= 9'h000; 
        10'b1011000010: data <= 9'h000; 
        10'b1011000011: data <= 9'h000; 
        10'b1011000100: data <= 9'h000; 
        10'b1011000101: data <= 9'h000; 
        10'b1011000110: data <= 9'h000; 
        10'b1011000111: data <= 9'h001; 
        10'b1011001000: data <= 9'h001; 
        10'b1011001001: data <= 9'h001; 
        10'b1011001010: data <= 9'h000; 
        10'b1011001011: data <= 9'h000; 
        10'b1011001100: data <= 9'h000; 
        10'b1011001101: data <= 9'h000; 
        10'b1011001110: data <= 9'h000; 
        10'b1011001111: data <= 9'h000; 
        10'b1011010000: data <= 9'h1ff; 
        10'b1011010001: data <= 9'h000; 
        10'b1011010010: data <= 9'h000; 
        10'b1011010011: data <= 9'h000; 
        10'b1011010100: data <= 9'h000; 
        10'b1011010101: data <= 9'h000; 
        10'b1011010110: data <= 9'h000; 
        10'b1011010111: data <= 9'h000; 
        10'b1011011000: data <= 9'h000; 
        10'b1011011001: data <= 9'h000; 
        10'b1011011010: data <= 9'h000; 
        10'b1011011011: data <= 9'h000; 
        10'b1011011100: data <= 9'h000; 
        10'b1011011101: data <= 9'h000; 
        10'b1011011110: data <= 9'h000; 
        10'b1011011111: data <= 9'h000; 
        10'b1011100000: data <= 9'h000; 
        10'b1011100001: data <= 9'h000; 
        10'b1011100010: data <= 9'h000; 
        10'b1011100011: data <= 9'h000; 
        10'b1011100100: data <= 9'h000; 
        10'b1011100101: data <= 9'h000; 
        10'b1011100110: data <= 9'h000; 
        10'b1011100111: data <= 9'h000; 
        10'b1011101000: data <= 9'h000; 
        10'b1011101001: data <= 9'h000; 
        10'b1011101010: data <= 9'h1ff; 
        10'b1011101011: data <= 9'h1ff; 
        10'b1011101100: data <= 9'h000; 
        10'b1011101101: data <= 9'h000; 
        10'b1011101110: data <= 9'h000; 
        10'b1011101111: data <= 9'h000; 
        10'b1011110000: data <= 9'h000; 
        10'b1011110001: data <= 9'h000; 
        10'b1011110010: data <= 9'h000; 
        10'b1011110011: data <= 9'h000; 
        10'b1011110100: data <= 9'h000; 
        10'b1011110101: data <= 9'h000; 
        10'b1011110110: data <= 9'h000; 
        10'b1011110111: data <= 9'h000; 
        10'b1011111000: data <= 9'h000; 
        10'b1011111001: data <= 9'h000; 
        10'b1011111010: data <= 9'h000; 
        10'b1011111011: data <= 9'h000; 
        10'b1011111100: data <= 9'h000; 
        10'b1011111101: data <= 9'h000; 
        10'b1011111110: data <= 9'h000; 
        10'b1011111111: data <= 9'h000; 
        10'b1100000000: data <= 9'h000; 
        10'b1100000001: data <= 9'h000; 
        10'b1100000010: data <= 9'h000; 
        10'b1100000011: data <= 9'h000; 
        10'b1100000100: data <= 9'h000; 
        10'b1100000101: data <= 9'h000; 
        10'b1100000110: data <= 9'h000; 
        10'b1100000111: data <= 9'h000; 
        10'b1100001000: data <= 9'h000; 
        10'b1100001001: data <= 9'h000; 
        10'b1100001010: data <= 9'h000; 
        10'b1100001011: data <= 9'h000; 
        10'b1100001100: data <= 9'h000; 
        10'b1100001101: data <= 9'h000; 
        10'b1100001110: data <= 9'h000; 
        10'b1100001111: data <= 9'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 4) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 10'h3ff; 
        10'b0000000001: data <= 10'h000; 
        10'b0000000010: data <= 10'h000; 
        10'b0000000011: data <= 10'h3ff; 
        10'b0000000100: data <= 10'h000; 
        10'b0000000101: data <= 10'h000; 
        10'b0000000110: data <= 10'h000; 
        10'b0000000111: data <= 10'h000; 
        10'b0000001000: data <= 10'h000; 
        10'b0000001001: data <= 10'h000; 
        10'b0000001010: data <= 10'h000; 
        10'b0000001011: data <= 10'h000; 
        10'b0000001100: data <= 10'h3ff; 
        10'b0000001101: data <= 10'h000; 
        10'b0000001110: data <= 10'h3ff; 
        10'b0000001111: data <= 10'h3ff; 
        10'b0000010000: data <= 10'h3ff; 
        10'b0000010001: data <= 10'h3ff; 
        10'b0000010010: data <= 10'h000; 
        10'b0000010011: data <= 10'h000; 
        10'b0000010100: data <= 10'h3ff; 
        10'b0000010101: data <= 10'h000; 
        10'b0000010110: data <= 10'h000; 
        10'b0000010111: data <= 10'h000; 
        10'b0000011000: data <= 10'h3ff; 
        10'b0000011001: data <= 10'h000; 
        10'b0000011010: data <= 10'h000; 
        10'b0000011011: data <= 10'h3ff; 
        10'b0000011100: data <= 10'h000; 
        10'b0000011101: data <= 10'h3ff; 
        10'b0000011110: data <= 10'h000; 
        10'b0000011111: data <= 10'h3ff; 
        10'b0000100000: data <= 10'h000; 
        10'b0000100001: data <= 10'h3ff; 
        10'b0000100010: data <= 10'h000; 
        10'b0000100011: data <= 10'h3ff; 
        10'b0000100100: data <= 10'h3ff; 
        10'b0000100101: data <= 10'h000; 
        10'b0000100110: data <= 10'h000; 
        10'b0000100111: data <= 10'h3ff; 
        10'b0000101000: data <= 10'h3ff; 
        10'b0000101001: data <= 10'h3ff; 
        10'b0000101010: data <= 10'h3ff; 
        10'b0000101011: data <= 10'h000; 
        10'b0000101100: data <= 10'h3ff; 
        10'b0000101101: data <= 10'h3ff; 
        10'b0000101110: data <= 10'h3ff; 
        10'b0000101111: data <= 10'h3ff; 
        10'b0000110000: data <= 10'h000; 
        10'b0000110001: data <= 10'h3ff; 
        10'b0000110010: data <= 10'h000; 
        10'b0000110011: data <= 10'h3ff; 
        10'b0000110100: data <= 10'h000; 
        10'b0000110101: data <= 10'h000; 
        10'b0000110110: data <= 10'h3ff; 
        10'b0000110111: data <= 10'h000; 
        10'b0000111000: data <= 10'h000; 
        10'b0000111001: data <= 10'h000; 
        10'b0000111010: data <= 10'h3ff; 
        10'b0000111011: data <= 10'h3ff; 
        10'b0000111100: data <= 10'h3ff; 
        10'b0000111101: data <= 10'h000; 
        10'b0000111110: data <= 10'h000; 
        10'b0000111111: data <= 10'h000; 
        10'b0001000000: data <= 10'h3ff; 
        10'b0001000001: data <= 10'h000; 
        10'b0001000010: data <= 10'h000; 
        10'b0001000011: data <= 10'h3ff; 
        10'b0001000100: data <= 10'h000; 
        10'b0001000101: data <= 10'h3ff; 
        10'b0001000110: data <= 10'h3ff; 
        10'b0001000111: data <= 10'h3ff; 
        10'b0001001000: data <= 10'h3ff; 
        10'b0001001001: data <= 10'h000; 
        10'b0001001010: data <= 10'h000; 
        10'b0001001011: data <= 10'h000; 
        10'b0001001100: data <= 10'h000; 
        10'b0001001101: data <= 10'h000; 
        10'b0001001110: data <= 10'h000; 
        10'b0001001111: data <= 10'h3ff; 
        10'b0001010000: data <= 10'h3ff; 
        10'b0001010001: data <= 10'h000; 
        10'b0001010010: data <= 10'h000; 
        10'b0001010011: data <= 10'h000; 
        10'b0001010100: data <= 10'h000; 
        10'b0001010101: data <= 10'h000; 
        10'b0001010110: data <= 10'h3ff; 
        10'b0001010111: data <= 10'h000; 
        10'b0001011000: data <= 10'h3ff; 
        10'b0001011001: data <= 10'h3ff; 
        10'b0001011010: data <= 10'h3ff; 
        10'b0001011011: data <= 10'h3ff; 
        10'b0001011100: data <= 10'h3ff; 
        10'b0001011101: data <= 10'h3ff; 
        10'b0001011110: data <= 10'h3ff; 
        10'b0001011111: data <= 10'h3fe; 
        10'b0001100000: data <= 10'h3ff; 
        10'b0001100001: data <= 10'h3ff; 
        10'b0001100010: data <= 10'h3ff; 
        10'b0001100011: data <= 10'h000; 
        10'b0001100100: data <= 10'h000; 
        10'b0001100101: data <= 10'h3ff; 
        10'b0001100110: data <= 10'h3ff; 
        10'b0001100111: data <= 10'h000; 
        10'b0001101000: data <= 10'h000; 
        10'b0001101001: data <= 10'h000; 
        10'b0001101010: data <= 10'h3ff; 
        10'b0001101011: data <= 10'h3ff; 
        10'b0001101100: data <= 10'h3ff; 
        10'b0001101101: data <= 10'h000; 
        10'b0001101110: data <= 10'h000; 
        10'b0001101111: data <= 10'h3ff; 
        10'b0001110000: data <= 10'h3ff; 
        10'b0001110001: data <= 10'h3ff; 
        10'b0001110010: data <= 10'h000; 
        10'b0001110011: data <= 10'h000; 
        10'b0001110100: data <= 10'h000; 
        10'b0001110101: data <= 10'h3ff; 
        10'b0001110110: data <= 10'h3ff; 
        10'b0001110111: data <= 10'h3ff; 
        10'b0001111000: data <= 10'h3fe; 
        10'b0001111001: data <= 10'h3fd; 
        10'b0001111010: data <= 10'h3fc; 
        10'b0001111011: data <= 10'h3fd; 
        10'b0001111100: data <= 10'h3fd; 
        10'b0001111101: data <= 10'h3fc; 
        10'b0001111110: data <= 10'h3fe; 
        10'b0001111111: data <= 10'h000; 
        10'b0010000000: data <= 10'h000; 
        10'b0010000001: data <= 10'h001; 
        10'b0010000010: data <= 10'h000; 
        10'b0010000011: data <= 10'h3ff; 
        10'b0010000100: data <= 10'h3ff; 
        10'b0010000101: data <= 10'h3ff; 
        10'b0010000110: data <= 10'h3ff; 
        10'b0010000111: data <= 10'h000; 
        10'b0010001000: data <= 10'h3ff; 
        10'b0010001001: data <= 10'h000; 
        10'b0010001010: data <= 10'h000; 
        10'b0010001011: data <= 10'h000; 
        10'b0010001100: data <= 10'h000; 
        10'b0010001101: data <= 10'h000; 
        10'b0010001110: data <= 10'h3ff; 
        10'b0010001111: data <= 10'h3ff; 
        10'b0010010000: data <= 10'h3ff; 
        10'b0010010001: data <= 10'h3ff; 
        10'b0010010010: data <= 10'h3fe; 
        10'b0010010011: data <= 10'h3fe; 
        10'b0010010100: data <= 10'h3ff; 
        10'b0010010101: data <= 10'h000; 
        10'b0010010110: data <= 10'h000; 
        10'b0010010111: data <= 10'h000; 
        10'b0010011000: data <= 10'h3ff; 
        10'b0010011001: data <= 10'h3ff; 
        10'b0010011010: data <= 10'h3ff; 
        10'b0010011011: data <= 10'h000; 
        10'b0010011100: data <= 10'h001; 
        10'b0010011101: data <= 10'h001; 
        10'b0010011110: data <= 10'h002; 
        10'b0010011111: data <= 10'h001; 
        10'b0010100000: data <= 10'h001; 
        10'b0010100001: data <= 10'h002; 
        10'b0010100010: data <= 10'h003; 
        10'b0010100011: data <= 10'h002; 
        10'b0010100100: data <= 10'h002; 
        10'b0010100101: data <= 10'h001; 
        10'b0010100110: data <= 10'h001; 
        10'b0010100111: data <= 10'h000; 
        10'b0010101000: data <= 10'h3ff; 
        10'b0010101001: data <= 10'h3ff; 
        10'b0010101010: data <= 10'h000; 
        10'b0010101011: data <= 10'h3ff; 
        10'b0010101100: data <= 10'h3ff; 
        10'b0010101101: data <= 10'h3fe; 
        10'b0010101110: data <= 10'h3ff; 
        10'b0010101111: data <= 10'h000; 
        10'b0010110000: data <= 10'h000; 
        10'b0010110001: data <= 10'h001; 
        10'b0010110010: data <= 10'h002; 
        10'b0010110011: data <= 10'h002; 
        10'b0010110100: data <= 10'h000; 
        10'b0010110101: data <= 10'h001; 
        10'b0010110110: data <= 10'h000; 
        10'b0010110111: data <= 10'h3ff; 
        10'b0010111000: data <= 10'h3ff; 
        10'b0010111001: data <= 10'h000; 
        10'b0010111010: data <= 10'h000; 
        10'b0010111011: data <= 10'h002; 
        10'b0010111100: data <= 10'h001; 
        10'b0010111101: data <= 10'h001; 
        10'b0010111110: data <= 10'h004; 
        10'b0010111111: data <= 10'h005; 
        10'b0011000000: data <= 10'h005; 
        10'b0011000001: data <= 10'h003; 
        10'b0011000010: data <= 10'h001; 
        10'b0011000011: data <= 10'h000; 
        10'b0011000100: data <= 10'h000; 
        10'b0011000101: data <= 10'h000; 
        10'b0011000110: data <= 10'h000; 
        10'b0011000111: data <= 10'h3ff; 
        10'b0011001000: data <= 10'h3fd; 
        10'b0011001001: data <= 10'h3fd; 
        10'b0011001010: data <= 10'h3fe; 
        10'b0011001011: data <= 10'h000; 
        10'b0011001100: data <= 10'h001; 
        10'b0011001101: data <= 10'h003; 
        10'b0011001110: data <= 10'h003; 
        10'b0011001111: data <= 10'h002; 
        10'b0011010000: data <= 10'h001; 
        10'b0011010001: data <= 10'h000; 
        10'b0011010010: data <= 10'h3ff; 
        10'b0011010011: data <= 10'h000; 
        10'b0011010100: data <= 10'h001; 
        10'b0011010101: data <= 10'h001; 
        10'b0011010110: data <= 10'h001; 
        10'b0011010111: data <= 10'h003; 
        10'b0011011000: data <= 10'h002; 
        10'b0011011001: data <= 10'h003; 
        10'b0011011010: data <= 10'h004; 
        10'b0011011011: data <= 10'h005; 
        10'b0011011100: data <= 10'h007; 
        10'b0011011101: data <= 10'h005; 
        10'b0011011110: data <= 10'h001; 
        10'b0011011111: data <= 10'h000; 
        10'b0011100000: data <= 10'h000; 
        10'b0011100001: data <= 10'h000; 
        10'b0011100010: data <= 10'h000; 
        10'b0011100011: data <= 10'h3ff; 
        10'b0011100100: data <= 10'h3fc; 
        10'b0011100101: data <= 10'h3fd; 
        10'b0011100110: data <= 10'h3fd; 
        10'b0011100111: data <= 10'h000; 
        10'b0011101000: data <= 10'h002; 
        10'b0011101001: data <= 10'h001; 
        10'b0011101010: data <= 10'h001; 
        10'b0011101011: data <= 10'h002; 
        10'b0011101100: data <= 10'h001; 
        10'b0011101101: data <= 10'h3ff; 
        10'b0011101110: data <= 10'h3fd; 
        10'b0011101111: data <= 10'h3fe; 
        10'b0011110000: data <= 10'h3ff; 
        10'b0011110001: data <= 10'h000; 
        10'b0011110010: data <= 10'h000; 
        10'b0011110011: data <= 10'h002; 
        10'b0011110100: data <= 10'h002; 
        10'b0011110101: data <= 10'h004; 
        10'b0011110110: data <= 10'h006; 
        10'b0011110111: data <= 10'h007; 
        10'b0011111000: data <= 10'h00a; 
        10'b0011111001: data <= 10'h006; 
        10'b0011111010: data <= 10'h001; 
        10'b0011111011: data <= 10'h000; 
        10'b0011111100: data <= 10'h3ff; 
        10'b0011111101: data <= 10'h000; 
        10'b0011111110: data <= 10'h3ff; 
        10'b0011111111: data <= 10'h3fe; 
        10'b0100000000: data <= 10'h3fe; 
        10'b0100000001: data <= 10'h3fe; 
        10'b0100000010: data <= 10'h000; 
        10'b0100000011: data <= 10'h000; 
        10'b0100000100: data <= 10'h002; 
        10'b0100000101: data <= 10'h001; 
        10'b0100000110: data <= 10'h002; 
        10'b0100000111: data <= 10'h004; 
        10'b0100001000: data <= 10'h003; 
        10'b0100001001: data <= 10'h3ff; 
        10'b0100001010: data <= 10'h3fc; 
        10'b0100001011: data <= 10'h3fb; 
        10'b0100001100: data <= 10'h3fb; 
        10'b0100001101: data <= 10'h3fd; 
        10'b0100001110: data <= 10'h3ff; 
        10'b0100001111: data <= 10'h000; 
        10'b0100010000: data <= 10'h002; 
        10'b0100010001: data <= 10'h005; 
        10'b0100010010: data <= 10'h007; 
        10'b0100010011: data <= 10'h00a; 
        10'b0100010100: data <= 10'h00c; 
        10'b0100010101: data <= 10'h008; 
        10'b0100010110: data <= 10'h001; 
        10'b0100010111: data <= 10'h3ff; 
        10'b0100011000: data <= 10'h000; 
        10'b0100011001: data <= 10'h3ff; 
        10'b0100011010: data <= 10'h3ff; 
        10'b0100011011: data <= 10'h3ff; 
        10'b0100011100: data <= 10'h3ff; 
        10'b0100011101: data <= 10'h000; 
        10'b0100011110: data <= 10'h001; 
        10'b0100011111: data <= 10'h003; 
        10'b0100100000: data <= 10'h004; 
        10'b0100100001: data <= 10'h004; 
        10'b0100100010: data <= 10'h004; 
        10'b0100100011: data <= 10'h005; 
        10'b0100100100: data <= 10'h004; 
        10'b0100100101: data <= 10'h003; 
        10'b0100100110: data <= 10'h3ff; 
        10'b0100100111: data <= 10'h3fd; 
        10'b0100101000: data <= 10'h3fc; 
        10'b0100101001: data <= 10'h3fc; 
        10'b0100101010: data <= 10'h3fc; 
        10'b0100101011: data <= 10'h3fb; 
        10'b0100101100: data <= 10'h3fd; 
        10'b0100101101: data <= 10'h3ff; 
        10'b0100101110: data <= 10'h001; 
        10'b0100101111: data <= 10'h003; 
        10'b0100110000: data <= 10'h006; 
        10'b0100110001: data <= 10'h005; 
        10'b0100110010: data <= 10'h002; 
        10'b0100110011: data <= 10'h3ff; 
        10'b0100110100: data <= 10'h3ff; 
        10'b0100110101: data <= 10'h000; 
        10'b0100110110: data <= 10'h3ff; 
        10'b0100110111: data <= 10'h000; 
        10'b0100111000: data <= 10'h3ff; 
        10'b0100111001: data <= 10'h000; 
        10'b0100111010: data <= 10'h002; 
        10'b0100111011: data <= 10'h003; 
        10'b0100111100: data <= 10'h004; 
        10'b0100111101: data <= 10'h004; 
        10'b0100111110: data <= 10'h003; 
        10'b0100111111: data <= 10'h003; 
        10'b0101000000: data <= 10'h005; 
        10'b0101000001: data <= 10'h004; 
        10'b0101000010: data <= 10'h000; 
        10'b0101000011: data <= 10'h3fd; 
        10'b0101000100: data <= 10'h3fd; 
        10'b0101000101: data <= 10'h3fc; 
        10'b0101000110: data <= 10'h3fb; 
        10'b0101000111: data <= 10'h3f9; 
        10'b0101001000: data <= 10'h3f6; 
        10'b0101001001: data <= 10'h3f7; 
        10'b0101001010: data <= 10'h3f9; 
        10'b0101001011: data <= 10'h3fb; 
        10'b0101001100: data <= 10'h3fe; 
        10'b0101001101: data <= 10'h000; 
        10'b0101001110: data <= 10'h001; 
        10'b0101001111: data <= 10'h000; 
        10'b0101010000: data <= 10'h000; 
        10'b0101010001: data <= 10'h000; 
        10'b0101010010: data <= 10'h000; 
        10'b0101010011: data <= 10'h3ff; 
        10'b0101010100: data <= 10'h000; 
        10'b0101010101: data <= 10'h001; 
        10'b0101010110: data <= 10'h002; 
        10'b0101010111: data <= 10'h002; 
        10'b0101011000: data <= 10'h002; 
        10'b0101011001: data <= 10'h001; 
        10'b0101011010: data <= 10'h003; 
        10'b0101011011: data <= 10'h006; 
        10'b0101011100: data <= 10'h005; 
        10'b0101011101: data <= 10'h005; 
        10'b0101011110: data <= 10'h001; 
        10'b0101011111: data <= 10'h3fd; 
        10'b0101100000: data <= 10'h3fb; 
        10'b0101100001: data <= 10'h3fc; 
        10'b0101100010: data <= 10'h3fd; 
        10'b0101100011: data <= 10'h3fc; 
        10'b0101100100: data <= 10'h3fb; 
        10'b0101100101: data <= 10'h3f8; 
        10'b0101100110: data <= 10'h3f7; 
        10'b0101100111: data <= 10'h3f8; 
        10'b0101101000: data <= 10'h3fb; 
        10'b0101101001: data <= 10'h3ff; 
        10'b0101101010: data <= 10'h000; 
        10'b0101101011: data <= 10'h000; 
        10'b0101101100: data <= 10'h000; 
        10'b0101101101: data <= 10'h3ff; 
        10'b0101101110: data <= 10'h3ff; 
        10'b0101101111: data <= 10'h3ff; 
        10'b0101110000: data <= 10'h000; 
        10'b0101110001: data <= 10'h001; 
        10'b0101110010: data <= 10'h002; 
        10'b0101110011: data <= 10'h001; 
        10'b0101110100: data <= 10'h001; 
        10'b0101110101: data <= 10'h001; 
        10'b0101110110: data <= 10'h004; 
        10'b0101110111: data <= 10'h004; 
        10'b0101111000: data <= 10'h003; 
        10'b0101111001: data <= 10'h003; 
        10'b0101111010: data <= 10'h3ff; 
        10'b0101111011: data <= 10'h3fd; 
        10'b0101111100: data <= 10'h3fb; 
        10'b0101111101: data <= 10'h3fd; 
        10'b0101111110: data <= 10'h3ff; 
        10'b0101111111: data <= 10'h3ff; 
        10'b0110000000: data <= 10'h3ff; 
        10'b0110000001: data <= 10'h3fe; 
        10'b0110000010: data <= 10'h3fc; 
        10'b0110000011: data <= 10'h3fa; 
        10'b0110000100: data <= 10'h3fc; 
        10'b0110000101: data <= 10'h3ff; 
        10'b0110000110: data <= 10'h3ff; 
        10'b0110000111: data <= 10'h000; 
        10'b0110001000: data <= 10'h000; 
        10'b0110001001: data <= 10'h3ff; 
        10'b0110001010: data <= 10'h000; 
        10'b0110001011: data <= 10'h3ff; 
        10'b0110001100: data <= 10'h000; 
        10'b0110001101: data <= 10'h000; 
        10'b0110001110: data <= 10'h000; 
        10'b0110001111: data <= 10'h000; 
        10'b0110010000: data <= 10'h002; 
        10'b0110010001: data <= 10'h003; 
        10'b0110010010: data <= 10'h003; 
        10'b0110010011: data <= 10'h001; 
        10'b0110010100: data <= 10'h001; 
        10'b0110010101: data <= 10'h000; 
        10'b0110010110: data <= 10'h3fe; 
        10'b0110010111: data <= 10'h3fd; 
        10'b0110011000: data <= 10'h3fc; 
        10'b0110011001: data <= 10'h3fd; 
        10'b0110011010: data <= 10'h3fd; 
        10'b0110011011: data <= 10'h3fe; 
        10'b0110011100: data <= 10'h3ff; 
        10'b0110011101: data <= 10'h3ff; 
        10'b0110011110: data <= 10'h3ff; 
        10'b0110011111: data <= 10'h3fd; 
        10'b0110100000: data <= 10'h3fe; 
        10'b0110100001: data <= 10'h3ff; 
        10'b0110100010: data <= 10'h000; 
        10'b0110100011: data <= 10'h3ff; 
        10'b0110100100: data <= 10'h3ff; 
        10'b0110100101: data <= 10'h000; 
        10'b0110100110: data <= 10'h3ff; 
        10'b0110100111: data <= 10'h000; 
        10'b0110101000: data <= 10'h3ff; 
        10'b0110101001: data <= 10'h3fe; 
        10'b0110101010: data <= 10'h3fd; 
        10'b0110101011: data <= 10'h3fe; 
        10'b0110101100: data <= 10'h001; 
        10'b0110101101: data <= 10'h003; 
        10'b0110101110: data <= 10'h001; 
        10'b0110101111: data <= 10'h001; 
        10'b0110110000: data <= 10'h001; 
        10'b0110110001: data <= 10'h3ff; 
        10'b0110110010: data <= 10'h3fc; 
        10'b0110110011: data <= 10'h3fc; 
        10'b0110110100: data <= 10'h3fc; 
        10'b0110110101: data <= 10'h3fc; 
        10'b0110110110: data <= 10'h3fd; 
        10'b0110110111: data <= 10'h000; 
        10'b0110111000: data <= 10'h3ff; 
        10'b0110111001: data <= 10'h3ff; 
        10'b0110111010: data <= 10'h3ff; 
        10'b0110111011: data <= 10'h3ff; 
        10'b0110111100: data <= 10'h3ff; 
        10'b0110111101: data <= 10'h000; 
        10'b0110111110: data <= 10'h000; 
        10'b0110111111: data <= 10'h3ff; 
        10'b0111000000: data <= 10'h3ff; 
        10'b0111000001: data <= 10'h000; 
        10'b0111000010: data <= 10'h000; 
        10'b0111000011: data <= 10'h3ff; 
        10'b0111000100: data <= 10'h3ff; 
        10'b0111000101: data <= 10'h3fe; 
        10'b0111000110: data <= 10'h3fb; 
        10'b0111000111: data <= 10'h3fb; 
        10'b0111001000: data <= 10'h3fc; 
        10'b0111001001: data <= 10'h3fe; 
        10'b0111001010: data <= 10'h3ff; 
        10'b0111001011: data <= 10'h3ff; 
        10'b0111001100: data <= 10'h3ff; 
        10'b0111001101: data <= 10'h3fd; 
        10'b0111001110: data <= 10'h3fb; 
        10'b0111001111: data <= 10'h3fc; 
        10'b0111010000: data <= 10'h3fd; 
        10'b0111010001: data <= 10'h3ff; 
        10'b0111010010: data <= 10'h3ff; 
        10'b0111010011: data <= 10'h000; 
        10'b0111010100: data <= 10'h001; 
        10'b0111010101: data <= 10'h000; 
        10'b0111010110: data <= 10'h001; 
        10'b0111010111: data <= 10'h000; 
        10'b0111011000: data <= 10'h000; 
        10'b0111011001: data <= 10'h000; 
        10'b0111011010: data <= 10'h3ff; 
        10'b0111011011: data <= 10'h000; 
        10'b0111011100: data <= 10'h3ff; 
        10'b0111011101: data <= 10'h000; 
        10'b0111011110: data <= 10'h000; 
        10'b0111011111: data <= 10'h000; 
        10'b0111100000: data <= 10'h3ff; 
        10'b0111100001: data <= 10'h000; 
        10'b0111100010: data <= 10'h000; 
        10'b0111100011: data <= 10'h3fc; 
        10'b0111100100: data <= 10'h3fa; 
        10'b0111100101: data <= 10'h3fa; 
        10'b0111100110: data <= 10'h3fc; 
        10'b0111100111: data <= 10'h3fd; 
        10'b0111101000: data <= 10'h3fc; 
        10'b0111101001: data <= 10'h3fb; 
        10'b0111101010: data <= 10'h3fb; 
        10'b0111101011: data <= 10'h3fe; 
        10'b0111101100: data <= 10'h3ff; 
        10'b0111101101: data <= 10'h002; 
        10'b0111101110: data <= 10'h002; 
        10'b0111101111: data <= 10'h002; 
        10'b0111110000: data <= 10'h002; 
        10'b0111110001: data <= 10'h000; 
        10'b0111110010: data <= 10'h000; 
        10'b0111110011: data <= 10'h001; 
        10'b0111110100: data <= 10'h001; 
        10'b0111110101: data <= 10'h3ff; 
        10'b0111110110: data <= 10'h000; 
        10'b0111110111: data <= 10'h000; 
        10'b0111111000: data <= 10'h000; 
        10'b0111111001: data <= 10'h3ff; 
        10'b0111111010: data <= 10'h000; 
        10'b0111111011: data <= 10'h3ff; 
        10'b0111111100: data <= 10'h001; 
        10'b0111111101: data <= 10'h002; 
        10'b0111111110: data <= 10'h004; 
        10'b0111111111: data <= 10'h001; 
        10'b1000000000: data <= 10'h3fc; 
        10'b1000000001: data <= 10'h3fa; 
        10'b1000000010: data <= 10'h3f9; 
        10'b1000000011: data <= 10'h3f9; 
        10'b1000000100: data <= 10'h3fb; 
        10'b1000000101: data <= 10'h3fd; 
        10'b1000000110: data <= 10'h3ff; 
        10'b1000000111: data <= 10'h3ff; 
        10'b1000001000: data <= 10'h000; 
        10'b1000001001: data <= 10'h002; 
        10'b1000001010: data <= 10'h001; 
        10'b1000001011: data <= 10'h002; 
        10'b1000001100: data <= 10'h001; 
        10'b1000001101: data <= 10'h002; 
        10'b1000001110: data <= 10'h001; 
        10'b1000001111: data <= 10'h002; 
        10'b1000010000: data <= 10'h001; 
        10'b1000010001: data <= 10'h000; 
        10'b1000010010: data <= 10'h3ff; 
        10'b1000010011: data <= 10'h000; 
        10'b1000010100: data <= 10'h000; 
        10'b1000010101: data <= 10'h3ff; 
        10'b1000010110: data <= 10'h000; 
        10'b1000010111: data <= 10'h000; 
        10'b1000011000: data <= 10'h002; 
        10'b1000011001: data <= 10'h003; 
        10'b1000011010: data <= 10'h004; 
        10'b1000011011: data <= 10'h003; 
        10'b1000011100: data <= 10'h002; 
        10'b1000011101: data <= 10'h001; 
        10'b1000011110: data <= 10'h3ff; 
        10'b1000011111: data <= 10'h3fe; 
        10'b1000100000: data <= 10'h000; 
        10'b1000100001: data <= 10'h002; 
        10'b1000100010: data <= 10'h001; 
        10'b1000100011: data <= 10'h001; 
        10'b1000100100: data <= 10'h001; 
        10'b1000100101: data <= 10'h000; 
        10'b1000100110: data <= 10'h001; 
        10'b1000100111: data <= 10'h001; 
        10'b1000101000: data <= 10'h000; 
        10'b1000101001: data <= 10'h001; 
        10'b1000101010: data <= 10'h002; 
        10'b1000101011: data <= 10'h001; 
        10'b1000101100: data <= 10'h000; 
        10'b1000101101: data <= 10'h000; 
        10'b1000101110: data <= 10'h000; 
        10'b1000101111: data <= 10'h3ff; 
        10'b1000110000: data <= 10'h000; 
        10'b1000110001: data <= 10'h3ff; 
        10'b1000110010: data <= 10'h000; 
        10'b1000110011: data <= 10'h3ff; 
        10'b1000110100: data <= 10'h000; 
        10'b1000110101: data <= 10'h002; 
        10'b1000110110: data <= 10'h003; 
        10'b1000110111: data <= 10'h003; 
        10'b1000111000: data <= 10'h004; 
        10'b1000111001: data <= 10'h004; 
        10'b1000111010: data <= 10'h003; 
        10'b1000111011: data <= 10'h005; 
        10'b1000111100: data <= 10'h003; 
        10'b1000111101: data <= 10'h002; 
        10'b1000111110: data <= 10'h3ff; 
        10'b1000111111: data <= 10'h3ff; 
        10'b1001000000: data <= 10'h002; 
        10'b1001000001: data <= 10'h001; 
        10'b1001000010: data <= 10'h001; 
        10'b1001000011: data <= 10'h002; 
        10'b1001000100: data <= 10'h002; 
        10'b1001000101: data <= 10'h001; 
        10'b1001000110: data <= 10'h003; 
        10'b1001000111: data <= 10'h002; 
        10'b1001001000: data <= 10'h000; 
        10'b1001001001: data <= 10'h3ff; 
        10'b1001001010: data <= 10'h000; 
        10'b1001001011: data <= 10'h3ff; 
        10'b1001001100: data <= 10'h3ff; 
        10'b1001001101: data <= 10'h000; 
        10'b1001001110: data <= 10'h3ff; 
        10'b1001001111: data <= 10'h000; 
        10'b1001010000: data <= 10'h001; 
        10'b1001010001: data <= 10'h000; 
        10'b1001010010: data <= 10'h001; 
        10'b1001010011: data <= 10'h003; 
        10'b1001010100: data <= 10'h004; 
        10'b1001010101: data <= 10'h003; 
        10'b1001010110: data <= 10'h002; 
        10'b1001010111: data <= 10'h001; 
        10'b1001011000: data <= 10'h002; 
        10'b1001011001: data <= 10'h001; 
        10'b1001011010: data <= 10'h001; 
        10'b1001011011: data <= 10'h001; 
        10'b1001011100: data <= 10'h000; 
        10'b1001011101: data <= 10'h001; 
        10'b1001011110: data <= 10'h001; 
        10'b1001011111: data <= 10'h002; 
        10'b1001100000: data <= 10'h002; 
        10'b1001100001: data <= 10'h003; 
        10'b1001100010: data <= 10'h003; 
        10'b1001100011: data <= 10'h001; 
        10'b1001100100: data <= 10'h000; 
        10'b1001100101: data <= 10'h3ff; 
        10'b1001100110: data <= 10'h3ff; 
        10'b1001100111: data <= 10'h3ff; 
        10'b1001101000: data <= 10'h000; 
        10'b1001101001: data <= 10'h3ff; 
        10'b1001101010: data <= 10'h000; 
        10'b1001101011: data <= 10'h3ff; 
        10'b1001101100: data <= 10'h000; 
        10'b1001101101: data <= 10'h000; 
        10'b1001101110: data <= 10'h3ff; 
        10'b1001101111: data <= 10'h000; 
        10'b1001110000: data <= 10'h002; 
        10'b1001110001: data <= 10'h002; 
        10'b1001110010: data <= 10'h000; 
        10'b1001110011: data <= 10'h002; 
        10'b1001110100: data <= 10'h003; 
        10'b1001110101: data <= 10'h004; 
        10'b1001110110: data <= 10'h002; 
        10'b1001110111: data <= 10'h000; 
        10'b1001111000: data <= 10'h000; 
        10'b1001111001: data <= 10'h001; 
        10'b1001111010: data <= 10'h001; 
        10'b1001111011: data <= 10'h001; 
        10'b1001111100: data <= 10'h002; 
        10'b1001111101: data <= 10'h002; 
        10'b1001111110: data <= 10'h002; 
        10'b1001111111: data <= 10'h001; 
        10'b1010000000: data <= 10'h000; 
        10'b1010000001: data <= 10'h000; 
        10'b1010000010: data <= 10'h000; 
        10'b1010000011: data <= 10'h000; 
        10'b1010000100: data <= 10'h3ff; 
        10'b1010000101: data <= 10'h000; 
        10'b1010000110: data <= 10'h000; 
        10'b1010000111: data <= 10'h000; 
        10'b1010001000: data <= 10'h3ff; 
        10'b1010001001: data <= 10'h000; 
        10'b1010001010: data <= 10'h3ff; 
        10'b1010001011: data <= 10'h3ff; 
        10'b1010001100: data <= 10'h001; 
        10'b1010001101: data <= 10'h001; 
        10'b1010001110: data <= 10'h001; 
        10'b1010001111: data <= 10'h002; 
        10'b1010010000: data <= 10'h002; 
        10'b1010010001: data <= 10'h001; 
        10'b1010010010: data <= 10'h002; 
        10'b1010010011: data <= 10'h002; 
        10'b1010010100: data <= 10'h001; 
        10'b1010010101: data <= 10'h001; 
        10'b1010010110: data <= 10'h3ff; 
        10'b1010010111: data <= 10'h000; 
        10'b1010011000: data <= 10'h001; 
        10'b1010011001: data <= 10'h000; 
        10'b1010011010: data <= 10'h001; 
        10'b1010011011: data <= 10'h3ff; 
        10'b1010011100: data <= 10'h000; 
        10'b1010011101: data <= 10'h000; 
        10'b1010011110: data <= 10'h3ff; 
        10'b1010011111: data <= 10'h000; 
        10'b1010100000: data <= 10'h000; 
        10'b1010100001: data <= 10'h000; 
        10'b1010100010: data <= 10'h3ff; 
        10'b1010100011: data <= 10'h000; 
        10'b1010100100: data <= 10'h3ff; 
        10'b1010100101: data <= 10'h3ff; 
        10'b1010100110: data <= 10'h000; 
        10'b1010100111: data <= 10'h000; 
        10'b1010101000: data <= 10'h000; 
        10'b1010101001: data <= 10'h002; 
        10'b1010101010: data <= 10'h002; 
        10'b1010101011: data <= 10'h002; 
        10'b1010101100: data <= 10'h001; 
        10'b1010101101: data <= 10'h001; 
        10'b1010101110: data <= 10'h003; 
        10'b1010101111: data <= 10'h002; 
        10'b1010110000: data <= 10'h001; 
        10'b1010110001: data <= 10'h001; 
        10'b1010110010: data <= 10'h001; 
        10'b1010110011: data <= 10'h001; 
        10'b1010110100: data <= 10'h000; 
        10'b1010110101: data <= 10'h000; 
        10'b1010110110: data <= 10'h000; 
        10'b1010110111: data <= 10'h000; 
        10'b1010111000: data <= 10'h3ff; 
        10'b1010111001: data <= 10'h000; 
        10'b1010111010: data <= 10'h000; 
        10'b1010111011: data <= 10'h3ff; 
        10'b1010111100: data <= 10'h000; 
        10'b1010111101: data <= 10'h000; 
        10'b1010111110: data <= 10'h000; 
        10'b1010111111: data <= 10'h3ff; 
        10'b1011000000: data <= 10'h000; 
        10'b1011000001: data <= 10'h000; 
        10'b1011000010: data <= 10'h3ff; 
        10'b1011000011: data <= 10'h000; 
        10'b1011000100: data <= 10'h3ff; 
        10'b1011000101: data <= 10'h001; 
        10'b1011000110: data <= 10'h000; 
        10'b1011000111: data <= 10'h001; 
        10'b1011001000: data <= 10'h001; 
        10'b1011001001: data <= 10'h002; 
        10'b1011001010: data <= 10'h000; 
        10'b1011001011: data <= 10'h001; 
        10'b1011001100: data <= 10'h000; 
        10'b1011001101: data <= 10'h001; 
        10'b1011001110: data <= 10'h3ff; 
        10'b1011001111: data <= 10'h000; 
        10'b1011010000: data <= 10'h3ff; 
        10'b1011010001: data <= 10'h000; 
        10'b1011010010: data <= 10'h000; 
        10'b1011010011: data <= 10'h3ff; 
        10'b1011010100: data <= 10'h000; 
        10'b1011010101: data <= 10'h000; 
        10'b1011010110: data <= 10'h3ff; 
        10'b1011010111: data <= 10'h000; 
        10'b1011011000: data <= 10'h000; 
        10'b1011011001: data <= 10'h000; 
        10'b1011011010: data <= 10'h3ff; 
        10'b1011011011: data <= 10'h000; 
        10'b1011011100: data <= 10'h3ff; 
        10'b1011011101: data <= 10'h000; 
        10'b1011011110: data <= 10'h000; 
        10'b1011011111: data <= 10'h3ff; 
        10'b1011100000: data <= 10'h3ff; 
        10'b1011100001: data <= 10'h000; 
        10'b1011100010: data <= 10'h3ff; 
        10'b1011100011: data <= 10'h000; 
        10'b1011100100: data <= 10'h000; 
        10'b1011100101: data <= 10'h000; 
        10'b1011100110: data <= 10'h3ff; 
        10'b1011100111: data <= 10'h000; 
        10'b1011101000: data <= 10'h000; 
        10'b1011101001: data <= 10'h3ff; 
        10'b1011101010: data <= 10'h3ff; 
        10'b1011101011: data <= 10'h3ff; 
        10'b1011101100: data <= 10'h000; 
        10'b1011101101: data <= 10'h000; 
        10'b1011101110: data <= 10'h3ff; 
        10'b1011101111: data <= 10'h000; 
        10'b1011110000: data <= 10'h000; 
        10'b1011110001: data <= 10'h000; 
        10'b1011110010: data <= 10'h3ff; 
        10'b1011110011: data <= 10'h3ff; 
        10'b1011110100: data <= 10'h000; 
        10'b1011110101: data <= 10'h000; 
        10'b1011110110: data <= 10'h000; 
        10'b1011110111: data <= 10'h000; 
        10'b1011111000: data <= 10'h3ff; 
        10'b1011111001: data <= 10'h000; 
        10'b1011111010: data <= 10'h3ff; 
        10'b1011111011: data <= 10'h3ff; 
        10'b1011111100: data <= 10'h000; 
        10'b1011111101: data <= 10'h3ff; 
        10'b1011111110: data <= 10'h3ff; 
        10'b1011111111: data <= 10'h000; 
        10'b1100000000: data <= 10'h000; 
        10'b1100000001: data <= 10'h3ff; 
        10'b1100000010: data <= 10'h000; 
        10'b1100000011: data <= 10'h000; 
        10'b1100000100: data <= 10'h3ff; 
        10'b1100000101: data <= 10'h3ff; 
        10'b1100000110: data <= 10'h3ff; 
        10'b1100000111: data <= 10'h3ff; 
        10'b1100001000: data <= 10'h000; 
        10'b1100001001: data <= 10'h3ff; 
        10'b1100001010: data <= 10'h000; 
        10'b1100001011: data <= 10'h3ff; 
        10'b1100001100: data <= 10'h000; 
        10'b1100001101: data <= 10'h000; 
        10'b1100001110: data <= 10'h3ff; 
        10'b1100001111: data <= 10'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 5) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 11'h7ff; 
        10'b0000000001: data <= 11'h000; 
        10'b0000000010: data <= 11'h000; 
        10'b0000000011: data <= 11'h7ff; 
        10'b0000000100: data <= 11'h7ff; 
        10'b0000000101: data <= 11'h7ff; 
        10'b0000000110: data <= 11'h000; 
        10'b0000000111: data <= 11'h7ff; 
        10'b0000001000: data <= 11'h000; 
        10'b0000001001: data <= 11'h000; 
        10'b0000001010: data <= 11'h000; 
        10'b0000001011: data <= 11'h000; 
        10'b0000001100: data <= 11'h7ff; 
        10'b0000001101: data <= 11'h000; 
        10'b0000001110: data <= 11'h7fe; 
        10'b0000001111: data <= 11'h7ff; 
        10'b0000010000: data <= 11'h7fe; 
        10'b0000010001: data <= 11'h7ff; 
        10'b0000010010: data <= 11'h000; 
        10'b0000010011: data <= 11'h000; 
        10'b0000010100: data <= 11'h7fe; 
        10'b0000010101: data <= 11'h7ff; 
        10'b0000010110: data <= 11'h000; 
        10'b0000010111: data <= 11'h7ff; 
        10'b0000011000: data <= 11'h7fe; 
        10'b0000011001: data <= 11'h7ff; 
        10'b0000011010: data <= 11'h000; 
        10'b0000011011: data <= 11'h7ff; 
        10'b0000011100: data <= 11'h000; 
        10'b0000011101: data <= 11'h7fe; 
        10'b0000011110: data <= 11'h000; 
        10'b0000011111: data <= 11'h7fe; 
        10'b0000100000: data <= 11'h000; 
        10'b0000100001: data <= 11'h7ff; 
        10'b0000100010: data <= 11'h7ff; 
        10'b0000100011: data <= 11'h7ff; 
        10'b0000100100: data <= 11'h7ff; 
        10'b0000100101: data <= 11'h000; 
        10'b0000100110: data <= 11'h000; 
        10'b0000100111: data <= 11'h7fe; 
        10'b0000101000: data <= 11'h7ff; 
        10'b0000101001: data <= 11'h7ff; 
        10'b0000101010: data <= 11'h7fe; 
        10'b0000101011: data <= 11'h000; 
        10'b0000101100: data <= 11'h7ff; 
        10'b0000101101: data <= 11'h7ff; 
        10'b0000101110: data <= 11'h7ff; 
        10'b0000101111: data <= 11'h7ff; 
        10'b0000110000: data <= 11'h000; 
        10'b0000110001: data <= 11'h7fe; 
        10'b0000110010: data <= 11'h000; 
        10'b0000110011: data <= 11'h7ff; 
        10'b0000110100: data <= 11'h000; 
        10'b0000110101: data <= 11'h000; 
        10'b0000110110: data <= 11'h7ff; 
        10'b0000110111: data <= 11'h7ff; 
        10'b0000111000: data <= 11'h7ff; 
        10'b0000111001: data <= 11'h000; 
        10'b0000111010: data <= 11'h7ff; 
        10'b0000111011: data <= 11'h7fe; 
        10'b0000111100: data <= 11'h7ff; 
        10'b0000111101: data <= 11'h7ff; 
        10'b0000111110: data <= 11'h000; 
        10'b0000111111: data <= 11'h000; 
        10'b0001000000: data <= 11'h7ff; 
        10'b0001000001: data <= 11'h7ff; 
        10'b0001000010: data <= 11'h000; 
        10'b0001000011: data <= 11'h7fe; 
        10'b0001000100: data <= 11'h000; 
        10'b0001000101: data <= 11'h7ff; 
        10'b0001000110: data <= 11'h7fe; 
        10'b0001000111: data <= 11'h7ff; 
        10'b0001001000: data <= 11'h7ff; 
        10'b0001001001: data <= 11'h7ff; 
        10'b0001001010: data <= 11'h7ff; 
        10'b0001001011: data <= 11'h7ff; 
        10'b0001001100: data <= 11'h000; 
        10'b0001001101: data <= 11'h000; 
        10'b0001001110: data <= 11'h000; 
        10'b0001001111: data <= 11'h7ff; 
        10'b0001010000: data <= 11'h7fe; 
        10'b0001010001: data <= 11'h7ff; 
        10'b0001010010: data <= 11'h000; 
        10'b0001010011: data <= 11'h000; 
        10'b0001010100: data <= 11'h000; 
        10'b0001010101: data <= 11'h7ff; 
        10'b0001010110: data <= 11'h7ff; 
        10'b0001010111: data <= 11'h000; 
        10'b0001011000: data <= 11'h7fe; 
        10'b0001011001: data <= 11'h7ff; 
        10'b0001011010: data <= 11'h7fe; 
        10'b0001011011: data <= 11'h7ff; 
        10'b0001011100: data <= 11'h7fe; 
        10'b0001011101: data <= 11'h7ff; 
        10'b0001011110: data <= 11'h7fd; 
        10'b0001011111: data <= 11'h7fc; 
        10'b0001100000: data <= 11'h7fe; 
        10'b0001100001: data <= 11'h7fe; 
        10'b0001100010: data <= 11'h7fd; 
        10'b0001100011: data <= 11'h7ff; 
        10'b0001100100: data <= 11'h000; 
        10'b0001100101: data <= 11'h7fe; 
        10'b0001100110: data <= 11'h7ff; 
        10'b0001100111: data <= 11'h000; 
        10'b0001101000: data <= 11'h000; 
        10'b0001101001: data <= 11'h7ff; 
        10'b0001101010: data <= 11'h7fe; 
        10'b0001101011: data <= 11'h7ff; 
        10'b0001101100: data <= 11'h7fe; 
        10'b0001101101: data <= 11'h000; 
        10'b0001101110: data <= 11'h000; 
        10'b0001101111: data <= 11'h7fe; 
        10'b0001110000: data <= 11'h7fe; 
        10'b0001110001: data <= 11'h7ff; 
        10'b0001110010: data <= 11'h000; 
        10'b0001110011: data <= 11'h000; 
        10'b0001110100: data <= 11'h000; 
        10'b0001110101: data <= 11'h7ff; 
        10'b0001110110: data <= 11'h7ff; 
        10'b0001110111: data <= 11'h7fd; 
        10'b0001111000: data <= 11'h7fb; 
        10'b0001111001: data <= 11'h7fa; 
        10'b0001111010: data <= 11'h7f7; 
        10'b0001111011: data <= 11'h7fa; 
        10'b0001111100: data <= 11'h7fa; 
        10'b0001111101: data <= 11'h7f8; 
        10'b0001111110: data <= 11'h7fc; 
        10'b0001111111: data <= 11'h000; 
        10'b0010000000: data <= 11'h000; 
        10'b0010000001: data <= 11'h001; 
        10'b0010000010: data <= 11'h000; 
        10'b0010000011: data <= 11'h7fe; 
        10'b0010000100: data <= 11'h7fd; 
        10'b0010000101: data <= 11'h7ff; 
        10'b0010000110: data <= 11'h7ff; 
        10'b0010000111: data <= 11'h7ff; 
        10'b0010001000: data <= 11'h7ff; 
        10'b0010001001: data <= 11'h000; 
        10'b0010001010: data <= 11'h000; 
        10'b0010001011: data <= 11'h7ff; 
        10'b0010001100: data <= 11'h7ff; 
        10'b0010001101: data <= 11'h000; 
        10'b0010001110: data <= 11'h7ff; 
        10'b0010001111: data <= 11'h7fe; 
        10'b0010010000: data <= 11'h7ff; 
        10'b0010010001: data <= 11'h7fd; 
        10'b0010010010: data <= 11'h7fc; 
        10'b0010010011: data <= 11'h7fc; 
        10'b0010010100: data <= 11'h7fd; 
        10'b0010010101: data <= 11'h000; 
        10'b0010010110: data <= 11'h001; 
        10'b0010010111: data <= 11'h001; 
        10'b0010011000: data <= 11'h7ff; 
        10'b0010011001: data <= 11'h7fe; 
        10'b0010011010: data <= 11'h7ff; 
        10'b0010011011: data <= 11'h7ff; 
        10'b0010011100: data <= 11'h002; 
        10'b0010011101: data <= 11'h002; 
        10'b0010011110: data <= 11'h004; 
        10'b0010011111: data <= 11'h002; 
        10'b0010100000: data <= 11'h002; 
        10'b0010100001: data <= 11'h003; 
        10'b0010100010: data <= 11'h006; 
        10'b0010100011: data <= 11'h005; 
        10'b0010100100: data <= 11'h003; 
        10'b0010100101: data <= 11'h002; 
        10'b0010100110: data <= 11'h001; 
        10'b0010100111: data <= 11'h000; 
        10'b0010101000: data <= 11'h7fe; 
        10'b0010101001: data <= 11'h7fe; 
        10'b0010101010: data <= 11'h000; 
        10'b0010101011: data <= 11'h7fe; 
        10'b0010101100: data <= 11'h7fe; 
        10'b0010101101: data <= 11'h7fb; 
        10'b0010101110: data <= 11'h7fe; 
        10'b0010101111: data <= 11'h000; 
        10'b0010110000: data <= 11'h000; 
        10'b0010110001: data <= 11'h002; 
        10'b0010110010: data <= 11'h004; 
        10'b0010110011: data <= 11'h003; 
        10'b0010110100: data <= 11'h001; 
        10'b0010110101: data <= 11'h001; 
        10'b0010110110: data <= 11'h7ff; 
        10'b0010110111: data <= 11'h7fe; 
        10'b0010111000: data <= 11'h7ff; 
        10'b0010111001: data <= 11'h7ff; 
        10'b0010111010: data <= 11'h000; 
        10'b0010111011: data <= 11'h004; 
        10'b0010111100: data <= 11'h002; 
        10'b0010111101: data <= 11'h003; 
        10'b0010111110: data <= 11'h008; 
        10'b0010111111: data <= 11'h009; 
        10'b0011000000: data <= 11'h00a; 
        10'b0011000001: data <= 11'h006; 
        10'b0011000010: data <= 11'h003; 
        10'b0011000011: data <= 11'h001; 
        10'b0011000100: data <= 11'h7ff; 
        10'b0011000101: data <= 11'h000; 
        10'b0011000110: data <= 11'h7ff; 
        10'b0011000111: data <= 11'h7fe; 
        10'b0011001000: data <= 11'h7fa; 
        10'b0011001001: data <= 11'h7f9; 
        10'b0011001010: data <= 11'h7fc; 
        10'b0011001011: data <= 11'h001; 
        10'b0011001100: data <= 11'h003; 
        10'b0011001101: data <= 11'h005; 
        10'b0011001110: data <= 11'h005; 
        10'b0011001111: data <= 11'h004; 
        10'b0011010000: data <= 11'h001; 
        10'b0011010001: data <= 11'h000; 
        10'b0011010010: data <= 11'h7ff; 
        10'b0011010011: data <= 11'h000; 
        10'b0011010100: data <= 11'h002; 
        10'b0011010101: data <= 11'h002; 
        10'b0011010110: data <= 11'h003; 
        10'b0011010111: data <= 11'h006; 
        10'b0011011000: data <= 11'h005; 
        10'b0011011001: data <= 11'h006; 
        10'b0011011010: data <= 11'h008; 
        10'b0011011011: data <= 11'h00b; 
        10'b0011011100: data <= 11'h00d; 
        10'b0011011101: data <= 11'h00a; 
        10'b0011011110: data <= 11'h001; 
        10'b0011011111: data <= 11'h000; 
        10'b0011100000: data <= 11'h000; 
        10'b0011100001: data <= 11'h000; 
        10'b0011100010: data <= 11'h000; 
        10'b0011100011: data <= 11'h7fd; 
        10'b0011100100: data <= 11'h7f8; 
        10'b0011100101: data <= 11'h7f9; 
        10'b0011100110: data <= 11'h7fb; 
        10'b0011100111: data <= 11'h000; 
        10'b0011101000: data <= 11'h004; 
        10'b0011101001: data <= 11'h001; 
        10'b0011101010: data <= 11'h002; 
        10'b0011101011: data <= 11'h004; 
        10'b0011101100: data <= 11'h003; 
        10'b0011101101: data <= 11'h7fd; 
        10'b0011101110: data <= 11'h7fa; 
        10'b0011101111: data <= 11'h7fc; 
        10'b0011110000: data <= 11'h7fe; 
        10'b0011110001: data <= 11'h000; 
        10'b0011110010: data <= 11'h001; 
        10'b0011110011: data <= 11'h005; 
        10'b0011110100: data <= 11'h005; 
        10'b0011110101: data <= 11'h007; 
        10'b0011110110: data <= 11'h00b; 
        10'b0011110111: data <= 11'h00f; 
        10'b0011111000: data <= 11'h013; 
        10'b0011111001: data <= 11'h00d; 
        10'b0011111010: data <= 11'h002; 
        10'b0011111011: data <= 11'h000; 
        10'b0011111100: data <= 11'h7fe; 
        10'b0011111101: data <= 11'h7ff; 
        10'b0011111110: data <= 11'h7fe; 
        10'b0011111111: data <= 11'h7fc; 
        10'b0100000000: data <= 11'h7fc; 
        10'b0100000001: data <= 11'h7fc; 
        10'b0100000010: data <= 11'h000; 
        10'b0100000011: data <= 11'h000; 
        10'b0100000100: data <= 11'h003; 
        10'b0100000101: data <= 11'h003; 
        10'b0100000110: data <= 11'h003; 
        10'b0100000111: data <= 11'h008; 
        10'b0100001000: data <= 11'h005; 
        10'b0100001001: data <= 11'h7fe; 
        10'b0100001010: data <= 11'h7f9; 
        10'b0100001011: data <= 11'h7f5; 
        10'b0100001100: data <= 11'h7f6; 
        10'b0100001101: data <= 11'h7fa; 
        10'b0100001110: data <= 11'h7ff; 
        10'b0100001111: data <= 11'h000; 
        10'b0100010000: data <= 11'h005; 
        10'b0100010001: data <= 11'h00a; 
        10'b0100010010: data <= 11'h00e; 
        10'b0100010011: data <= 11'h013; 
        10'b0100010100: data <= 11'h018; 
        10'b0100010101: data <= 11'h010; 
        10'b0100010110: data <= 11'h003; 
        10'b0100010111: data <= 11'h7ff; 
        10'b0100011000: data <= 11'h000; 
        10'b0100011001: data <= 11'h7ff; 
        10'b0100011010: data <= 11'h7ff; 
        10'b0100011011: data <= 11'h7ff; 
        10'b0100011100: data <= 11'h7ff; 
        10'b0100011101: data <= 11'h7ff; 
        10'b0100011110: data <= 11'h003; 
        10'b0100011111: data <= 11'h005; 
        10'b0100100000: data <= 11'h008; 
        10'b0100100001: data <= 11'h009; 
        10'b0100100010: data <= 11'h008; 
        10'b0100100011: data <= 11'h00a; 
        10'b0100100100: data <= 11'h008; 
        10'b0100100101: data <= 11'h006; 
        10'b0100100110: data <= 11'h7ff; 
        10'b0100100111: data <= 11'h7fb; 
        10'b0100101000: data <= 11'h7f7; 
        10'b0100101001: data <= 11'h7f7; 
        10'b0100101010: data <= 11'h7f7; 
        10'b0100101011: data <= 11'h7f6; 
        10'b0100101100: data <= 11'h7f9; 
        10'b0100101101: data <= 11'h7fe; 
        10'b0100101110: data <= 11'h001; 
        10'b0100101111: data <= 11'h006; 
        10'b0100110000: data <= 11'h00d; 
        10'b0100110001: data <= 11'h00a; 
        10'b0100110010: data <= 11'h003; 
        10'b0100110011: data <= 11'h7ff; 
        10'b0100110100: data <= 11'h7fe; 
        10'b0100110101: data <= 11'h000; 
        10'b0100110110: data <= 11'h7ff; 
        10'b0100110111: data <= 11'h7ff; 
        10'b0100111000: data <= 11'h7ff; 
        10'b0100111001: data <= 11'h000; 
        10'b0100111010: data <= 11'h004; 
        10'b0100111011: data <= 11'h005; 
        10'b0100111100: data <= 11'h008; 
        10'b0100111101: data <= 11'h007; 
        10'b0100111110: data <= 11'h005; 
        10'b0100111111: data <= 11'h006; 
        10'b0101000000: data <= 11'h009; 
        10'b0101000001: data <= 11'h009; 
        10'b0101000010: data <= 11'h000; 
        10'b0101000011: data <= 11'h7fb; 
        10'b0101000100: data <= 11'h7f9; 
        10'b0101000101: data <= 11'h7f9; 
        10'b0101000110: data <= 11'h7f6; 
        10'b0101000111: data <= 11'h7f2; 
        10'b0101001000: data <= 11'h7ec; 
        10'b0101001001: data <= 11'h7ee; 
        10'b0101001010: data <= 11'h7f1; 
        10'b0101001011: data <= 11'h7f5; 
        10'b0101001100: data <= 11'h7fc; 
        10'b0101001101: data <= 11'h000; 
        10'b0101001110: data <= 11'h001; 
        10'b0101001111: data <= 11'h7ff; 
        10'b0101010000: data <= 11'h7ff; 
        10'b0101010001: data <= 11'h7ff; 
        10'b0101010010: data <= 11'h7ff; 
        10'b0101010011: data <= 11'h7ff; 
        10'b0101010100: data <= 11'h7ff; 
        10'b0101010101: data <= 11'h002; 
        10'b0101010110: data <= 11'h005; 
        10'b0101010111: data <= 11'h004; 
        10'b0101011000: data <= 11'h003; 
        10'b0101011001: data <= 11'h002; 
        10'b0101011010: data <= 11'h005; 
        10'b0101011011: data <= 11'h00b; 
        10'b0101011100: data <= 11'h00b; 
        10'b0101011101: data <= 11'h00b; 
        10'b0101011110: data <= 11'h001; 
        10'b0101011111: data <= 11'h7fb; 
        10'b0101100000: data <= 11'h7f6; 
        10'b0101100001: data <= 11'h7f8; 
        10'b0101100010: data <= 11'h7fa; 
        10'b0101100011: data <= 11'h7f8; 
        10'b0101100100: data <= 11'h7f7; 
        10'b0101100101: data <= 11'h7f1; 
        10'b0101100110: data <= 11'h7ef; 
        10'b0101100111: data <= 11'h7f1; 
        10'b0101101000: data <= 11'h7f6; 
        10'b0101101001: data <= 11'h7fd; 
        10'b0101101010: data <= 11'h000; 
        10'b0101101011: data <= 11'h000; 
        10'b0101101100: data <= 11'h7ff; 
        10'b0101101101: data <= 11'h7ff; 
        10'b0101101110: data <= 11'h7fe; 
        10'b0101101111: data <= 11'h7ff; 
        10'b0101110000: data <= 11'h000; 
        10'b0101110001: data <= 11'h001; 
        10'b0101110010: data <= 11'h003; 
        10'b0101110011: data <= 11'h002; 
        10'b0101110100: data <= 11'h003; 
        10'b0101110101: data <= 11'h002; 
        10'b0101110110: data <= 11'h008; 
        10'b0101110111: data <= 11'h009; 
        10'b0101111000: data <= 11'h006; 
        10'b0101111001: data <= 11'h006; 
        10'b0101111010: data <= 11'h7ff; 
        10'b0101111011: data <= 11'h7f9; 
        10'b0101111100: data <= 11'h7f5; 
        10'b0101111101: data <= 11'h7fa; 
        10'b0101111110: data <= 11'h7fe; 
        10'b0101111111: data <= 11'h7fe; 
        10'b0110000000: data <= 11'h7ff; 
        10'b0110000001: data <= 11'h7fc; 
        10'b0110000010: data <= 11'h7f8; 
        10'b0110000011: data <= 11'h7f5; 
        10'b0110000100: data <= 11'h7f7; 
        10'b0110000101: data <= 11'h7ff; 
        10'b0110000110: data <= 11'h7fe; 
        10'b0110000111: data <= 11'h000; 
        10'b0110001000: data <= 11'h7ff; 
        10'b0110001001: data <= 11'h7fe; 
        10'b0110001010: data <= 11'h7ff; 
        10'b0110001011: data <= 11'h7fe; 
        10'b0110001100: data <= 11'h7ff; 
        10'b0110001101: data <= 11'h7ff; 
        10'b0110001110: data <= 11'h000; 
        10'b0110001111: data <= 11'h000; 
        10'b0110010000: data <= 11'h003; 
        10'b0110010001: data <= 11'h006; 
        10'b0110010010: data <= 11'h007; 
        10'b0110010011: data <= 11'h001; 
        10'b0110010100: data <= 11'h002; 
        10'b0110010101: data <= 11'h000; 
        10'b0110010110: data <= 11'h7fb; 
        10'b0110010111: data <= 11'h7fb; 
        10'b0110011000: data <= 11'h7f8; 
        10'b0110011001: data <= 11'h7f9; 
        10'b0110011010: data <= 11'h7fa; 
        10'b0110011011: data <= 11'h7fd; 
        10'b0110011100: data <= 11'h7fd; 
        10'b0110011101: data <= 11'h7fe; 
        10'b0110011110: data <= 11'h7ff; 
        10'b0110011111: data <= 11'h7fa; 
        10'b0110100000: data <= 11'h7fc; 
        10'b0110100001: data <= 11'h7fe; 
        10'b0110100010: data <= 11'h7ff; 
        10'b0110100011: data <= 11'h7fe; 
        10'b0110100100: data <= 11'h7fe; 
        10'b0110100101: data <= 11'h000; 
        10'b0110100110: data <= 11'h7fe; 
        10'b0110100111: data <= 11'h7ff; 
        10'b0110101000: data <= 11'h7fd; 
        10'b0110101001: data <= 11'h7fc; 
        10'b0110101010: data <= 11'h7fa; 
        10'b0110101011: data <= 11'h7fc; 
        10'b0110101100: data <= 11'h001; 
        10'b0110101101: data <= 11'h006; 
        10'b0110101110: data <= 11'h003; 
        10'b0110101111: data <= 11'h003; 
        10'b0110110000: data <= 11'h002; 
        10'b0110110001: data <= 11'h7fe; 
        10'b0110110010: data <= 11'h7f9; 
        10'b0110110011: data <= 11'h7f8; 
        10'b0110110100: data <= 11'h7f9; 
        10'b0110110101: data <= 11'h7f8; 
        10'b0110110110: data <= 11'h7fb; 
        10'b0110110111: data <= 11'h000; 
        10'b0110111000: data <= 11'h7fe; 
        10'b0110111001: data <= 11'h7fe; 
        10'b0110111010: data <= 11'h7fe; 
        10'b0110111011: data <= 11'h7fe; 
        10'b0110111100: data <= 11'h7ff; 
        10'b0110111101: data <= 11'h000; 
        10'b0110111110: data <= 11'h000; 
        10'b0110111111: data <= 11'h7ff; 
        10'b0111000000: data <= 11'h7ff; 
        10'b0111000001: data <= 11'h7ff; 
        10'b0111000010: data <= 11'h000; 
        10'b0111000011: data <= 11'h7fe; 
        10'b0111000100: data <= 11'h7ff; 
        10'b0111000101: data <= 11'h7fb; 
        10'b0111000110: data <= 11'h7f7; 
        10'b0111000111: data <= 11'h7f5; 
        10'b0111001000: data <= 11'h7f9; 
        10'b0111001001: data <= 11'h7fc; 
        10'b0111001010: data <= 11'h7fe; 
        10'b0111001011: data <= 11'h7fe; 
        10'b0111001100: data <= 11'h7fe; 
        10'b0111001101: data <= 11'h7fb; 
        10'b0111001110: data <= 11'h7f6; 
        10'b0111001111: data <= 11'h7f8; 
        10'b0111010000: data <= 11'h7fa; 
        10'b0111010001: data <= 11'h7fe; 
        10'b0111010010: data <= 11'h7fe; 
        10'b0111010011: data <= 11'h000; 
        10'b0111010100: data <= 11'h002; 
        10'b0111010101: data <= 11'h000; 
        10'b0111010110: data <= 11'h002; 
        10'b0111010111: data <= 11'h000; 
        10'b0111011000: data <= 11'h000; 
        10'b0111011001: data <= 11'h000; 
        10'b0111011010: data <= 11'h7ff; 
        10'b0111011011: data <= 11'h7ff; 
        10'b0111011100: data <= 11'h7ff; 
        10'b0111011101: data <= 11'h000; 
        10'b0111011110: data <= 11'h000; 
        10'b0111011111: data <= 11'h000; 
        10'b0111100000: data <= 11'h7ff; 
        10'b0111100001: data <= 11'h000; 
        10'b0111100010: data <= 11'h001; 
        10'b0111100011: data <= 11'h7f9; 
        10'b0111100100: data <= 11'h7f3; 
        10'b0111100101: data <= 11'h7f4; 
        10'b0111100110: data <= 11'h7f7; 
        10'b0111100111: data <= 11'h7fb; 
        10'b0111101000: data <= 11'h7f8; 
        10'b0111101001: data <= 11'h7f5; 
        10'b0111101010: data <= 11'h7f6; 
        10'b0111101011: data <= 11'h7fb; 
        10'b0111101100: data <= 11'h7fe; 
        10'b0111101101: data <= 11'h003; 
        10'b0111101110: data <= 11'h005; 
        10'b0111101111: data <= 11'h003; 
        10'b0111110000: data <= 11'h003; 
        10'b0111110001: data <= 11'h001; 
        10'b0111110010: data <= 11'h000; 
        10'b0111110011: data <= 11'h002; 
        10'b0111110100: data <= 11'h002; 
        10'b0111110101: data <= 11'h7ff; 
        10'b0111110110: data <= 11'h000; 
        10'b0111110111: data <= 11'h000; 
        10'b0111111000: data <= 11'h000; 
        10'b0111111001: data <= 11'h7ff; 
        10'b0111111010: data <= 11'h7ff; 
        10'b0111111011: data <= 11'h7ff; 
        10'b0111111100: data <= 11'h003; 
        10'b0111111101: data <= 11'h003; 
        10'b0111111110: data <= 11'h008; 
        10'b0111111111: data <= 11'h001; 
        10'b1000000000: data <= 11'h7f8; 
        10'b1000000001: data <= 11'h7f5; 
        10'b1000000010: data <= 11'h7f1; 
        10'b1000000011: data <= 11'h7f3; 
        10'b1000000100: data <= 11'h7f6; 
        10'b1000000101: data <= 11'h7fb; 
        10'b1000000110: data <= 11'h7fd; 
        10'b1000000111: data <= 11'h7ff; 
        10'b1000001000: data <= 11'h000; 
        10'b1000001001: data <= 11'h004; 
        10'b1000001010: data <= 11'h002; 
        10'b1000001011: data <= 11'h003; 
        10'b1000001100: data <= 11'h002; 
        10'b1000001101: data <= 11'h003; 
        10'b1000001110: data <= 11'h003; 
        10'b1000001111: data <= 11'h004; 
        10'b1000010000: data <= 11'h002; 
        10'b1000010001: data <= 11'h000; 
        10'b1000010010: data <= 11'h7ff; 
        10'b1000010011: data <= 11'h000; 
        10'b1000010100: data <= 11'h000; 
        10'b1000010101: data <= 11'h7ff; 
        10'b1000010110: data <= 11'h7ff; 
        10'b1000010111: data <= 11'h000; 
        10'b1000011000: data <= 11'h004; 
        10'b1000011001: data <= 11'h007; 
        10'b1000011010: data <= 11'h009; 
        10'b1000011011: data <= 11'h006; 
        10'b1000011100: data <= 11'h004; 
        10'b1000011101: data <= 11'h001; 
        10'b1000011110: data <= 11'h7fd; 
        10'b1000011111: data <= 11'h7fd; 
        10'b1000100000: data <= 11'h000; 
        10'b1000100001: data <= 11'h004; 
        10'b1000100010: data <= 11'h001; 
        10'b1000100011: data <= 11'h002; 
        10'b1000100100: data <= 11'h002; 
        10'b1000100101: data <= 11'h7ff; 
        10'b1000100110: data <= 11'h001; 
        10'b1000100111: data <= 11'h001; 
        10'b1000101000: data <= 11'h000; 
        10'b1000101001: data <= 11'h002; 
        10'b1000101010: data <= 11'h004; 
        10'b1000101011: data <= 11'h003; 
        10'b1000101100: data <= 11'h000; 
        10'b1000101101: data <= 11'h000; 
        10'b1000101110: data <= 11'h000; 
        10'b1000101111: data <= 11'h7fe; 
        10'b1000110000: data <= 11'h000; 
        10'b1000110001: data <= 11'h7fe; 
        10'b1000110010: data <= 11'h7ff; 
        10'b1000110011: data <= 11'h7ff; 
        10'b1000110100: data <= 11'h001; 
        10'b1000110101: data <= 11'h004; 
        10'b1000110110: data <= 11'h005; 
        10'b1000110111: data <= 11'h006; 
        10'b1000111000: data <= 11'h009; 
        10'b1000111001: data <= 11'h007; 
        10'b1000111010: data <= 11'h006; 
        10'b1000111011: data <= 11'h009; 
        10'b1000111100: data <= 11'h006; 
        10'b1000111101: data <= 11'h004; 
        10'b1000111110: data <= 11'h7ff; 
        10'b1000111111: data <= 11'h7ff; 
        10'b1001000000: data <= 11'h003; 
        10'b1001000001: data <= 11'h002; 
        10'b1001000010: data <= 11'h003; 
        10'b1001000011: data <= 11'h004; 
        10'b1001000100: data <= 11'h003; 
        10'b1001000101: data <= 11'h002; 
        10'b1001000110: data <= 11'h006; 
        10'b1001000111: data <= 11'h004; 
        10'b1001001000: data <= 11'h7ff; 
        10'b1001001001: data <= 11'h7fe; 
        10'b1001001010: data <= 11'h7ff; 
        10'b1001001011: data <= 11'h7ff; 
        10'b1001001100: data <= 11'h7ff; 
        10'b1001001101: data <= 11'h000; 
        10'b1001001110: data <= 11'h7fe; 
        10'b1001001111: data <= 11'h7ff; 
        10'b1001010000: data <= 11'h002; 
        10'b1001010001: data <= 11'h7ff; 
        10'b1001010010: data <= 11'h002; 
        10'b1001010011: data <= 11'h006; 
        10'b1001010100: data <= 11'h008; 
        10'b1001010101: data <= 11'h005; 
        10'b1001010110: data <= 11'h005; 
        10'b1001010111: data <= 11'h002; 
        10'b1001011000: data <= 11'h003; 
        10'b1001011001: data <= 11'h002; 
        10'b1001011010: data <= 11'h002; 
        10'b1001011011: data <= 11'h002; 
        10'b1001011100: data <= 11'h001; 
        10'b1001011101: data <= 11'h002; 
        10'b1001011110: data <= 11'h001; 
        10'b1001011111: data <= 11'h003; 
        10'b1001100000: data <= 11'h003; 
        10'b1001100001: data <= 11'h005; 
        10'b1001100010: data <= 11'h007; 
        10'b1001100011: data <= 11'h001; 
        10'b1001100100: data <= 11'h000; 
        10'b1001100101: data <= 11'h7fe; 
        10'b1001100110: data <= 11'h7ff; 
        10'b1001100111: data <= 11'h7ff; 
        10'b1001101000: data <= 11'h000; 
        10'b1001101001: data <= 11'h7fe; 
        10'b1001101010: data <= 11'h7ff; 
        10'b1001101011: data <= 11'h7ff; 
        10'b1001101100: data <= 11'h001; 
        10'b1001101101: data <= 11'h7ff; 
        10'b1001101110: data <= 11'h7fe; 
        10'b1001101111: data <= 11'h000; 
        10'b1001110000: data <= 11'h003; 
        10'b1001110001: data <= 11'h005; 
        10'b1001110010: data <= 11'h001; 
        10'b1001110011: data <= 11'h004; 
        10'b1001110100: data <= 11'h007; 
        10'b1001110101: data <= 11'h008; 
        10'b1001110110: data <= 11'h004; 
        10'b1001110111: data <= 11'h001; 
        10'b1001111000: data <= 11'h000; 
        10'b1001111001: data <= 11'h001; 
        10'b1001111010: data <= 11'h002; 
        10'b1001111011: data <= 11'h002; 
        10'b1001111100: data <= 11'h004; 
        10'b1001111101: data <= 11'h003; 
        10'b1001111110: data <= 11'h003; 
        10'b1001111111: data <= 11'h001; 
        10'b1010000000: data <= 11'h000; 
        10'b1010000001: data <= 11'h000; 
        10'b1010000010: data <= 11'h7ff; 
        10'b1010000011: data <= 11'h000; 
        10'b1010000100: data <= 11'h7ff; 
        10'b1010000101: data <= 11'h7ff; 
        10'b1010000110: data <= 11'h000; 
        10'b1010000111: data <= 11'h7ff; 
        10'b1010001000: data <= 11'h7ff; 
        10'b1010001001: data <= 11'h7ff; 
        10'b1010001010: data <= 11'h7fd; 
        10'b1010001011: data <= 11'h7ff; 
        10'b1010001100: data <= 11'h003; 
        10'b1010001101: data <= 11'h002; 
        10'b1010001110: data <= 11'h002; 
        10'b1010001111: data <= 11'h004; 
        10'b1010010000: data <= 11'h004; 
        10'b1010010001: data <= 11'h003; 
        10'b1010010010: data <= 11'h003; 
        10'b1010010011: data <= 11'h003; 
        10'b1010010100: data <= 11'h003; 
        10'b1010010101: data <= 11'h001; 
        10'b1010010110: data <= 11'h7fe; 
        10'b1010010111: data <= 11'h000; 
        10'b1010011000: data <= 11'h001; 
        10'b1010011001: data <= 11'h001; 
        10'b1010011010: data <= 11'h002; 
        10'b1010011011: data <= 11'h7ff; 
        10'b1010011100: data <= 11'h000; 
        10'b1010011101: data <= 11'h7ff; 
        10'b1010011110: data <= 11'h7ff; 
        10'b1010011111: data <= 11'h000; 
        10'b1010100000: data <= 11'h000; 
        10'b1010100001: data <= 11'h7ff; 
        10'b1010100010: data <= 11'h7ff; 
        10'b1010100011: data <= 11'h000; 
        10'b1010100100: data <= 11'h7fe; 
        10'b1010100101: data <= 11'h7fe; 
        10'b1010100110: data <= 11'h7ff; 
        10'b1010100111: data <= 11'h000; 
        10'b1010101000: data <= 11'h000; 
        10'b1010101001: data <= 11'h003; 
        10'b1010101010: data <= 11'h004; 
        10'b1010101011: data <= 11'h003; 
        10'b1010101100: data <= 11'h002; 
        10'b1010101101: data <= 11'h003; 
        10'b1010101110: data <= 11'h005; 
        10'b1010101111: data <= 11'h004; 
        10'b1010110000: data <= 11'h003; 
        10'b1010110001: data <= 11'h001; 
        10'b1010110010: data <= 11'h002; 
        10'b1010110011: data <= 11'h002; 
        10'b1010110100: data <= 11'h000; 
        10'b1010110101: data <= 11'h000; 
        10'b1010110110: data <= 11'h7ff; 
        10'b1010110111: data <= 11'h000; 
        10'b1010111000: data <= 11'h7ff; 
        10'b1010111001: data <= 11'h000; 
        10'b1010111010: data <= 11'h000; 
        10'b1010111011: data <= 11'h7fe; 
        10'b1010111100: data <= 11'h7ff; 
        10'b1010111101: data <= 11'h000; 
        10'b1010111110: data <= 11'h000; 
        10'b1010111111: data <= 11'h7fe; 
        10'b1011000000: data <= 11'h000; 
        10'b1011000001: data <= 11'h7ff; 
        10'b1011000010: data <= 11'h7fe; 
        10'b1011000011: data <= 11'h7ff; 
        10'b1011000100: data <= 11'h7fe; 
        10'b1011000101: data <= 11'h001; 
        10'b1011000110: data <= 11'h001; 
        10'b1011000111: data <= 11'h002; 
        10'b1011001000: data <= 11'h002; 
        10'b1011001001: data <= 11'h004; 
        10'b1011001010: data <= 11'h000; 
        10'b1011001011: data <= 11'h001; 
        10'b1011001100: data <= 11'h001; 
        10'b1011001101: data <= 11'h002; 
        10'b1011001110: data <= 11'h7ff; 
        10'b1011001111: data <= 11'h000; 
        10'b1011010000: data <= 11'h7fe; 
        10'b1011010001: data <= 11'h000; 
        10'b1011010010: data <= 11'h7ff; 
        10'b1011010011: data <= 11'h7ff; 
        10'b1011010100: data <= 11'h000; 
        10'b1011010101: data <= 11'h000; 
        10'b1011010110: data <= 11'h7fe; 
        10'b1011010111: data <= 11'h7ff; 
        10'b1011011000: data <= 11'h7ff; 
        10'b1011011001: data <= 11'h7ff; 
        10'b1011011010: data <= 11'h7ff; 
        10'b1011011011: data <= 11'h7ff; 
        10'b1011011100: data <= 11'h7ff; 
        10'b1011011101: data <= 11'h7ff; 
        10'b1011011110: data <= 11'h000; 
        10'b1011011111: data <= 11'h7ff; 
        10'b1011100000: data <= 11'h7fe; 
        10'b1011100001: data <= 11'h7ff; 
        10'b1011100010: data <= 11'h7ff; 
        10'b1011100011: data <= 11'h000; 
        10'b1011100100: data <= 11'h000; 
        10'b1011100101: data <= 11'h000; 
        10'b1011100110: data <= 11'h7ff; 
        10'b1011100111: data <= 11'h7ff; 
        10'b1011101000: data <= 11'h000; 
        10'b1011101001: data <= 11'h7ff; 
        10'b1011101010: data <= 11'h7fd; 
        10'b1011101011: data <= 11'h7fe; 
        10'b1011101100: data <= 11'h000; 
        10'b1011101101: data <= 11'h000; 
        10'b1011101110: data <= 11'h7ff; 
        10'b1011101111: data <= 11'h000; 
        10'b1011110000: data <= 11'h7ff; 
        10'b1011110001: data <= 11'h7ff; 
        10'b1011110010: data <= 11'h7ff; 
        10'b1011110011: data <= 11'h7fe; 
        10'b1011110100: data <= 11'h000; 
        10'b1011110101: data <= 11'h000; 
        10'b1011110110: data <= 11'h000; 
        10'b1011110111: data <= 11'h7ff; 
        10'b1011111000: data <= 11'h7fe; 
        10'b1011111001: data <= 11'h000; 
        10'b1011111010: data <= 11'h7ff; 
        10'b1011111011: data <= 11'h7ff; 
        10'b1011111100: data <= 11'h000; 
        10'b1011111101: data <= 11'h7ff; 
        10'b1011111110: data <= 11'h7ff; 
        10'b1011111111: data <= 11'h000; 
        10'b1100000000: data <= 11'h7ff; 
        10'b1100000001: data <= 11'h7fe; 
        10'b1100000010: data <= 11'h000; 
        10'b1100000011: data <= 11'h7ff; 
        10'b1100000100: data <= 11'h7fe; 
        10'b1100000101: data <= 11'h7fe; 
        10'b1100000110: data <= 11'h7ff; 
        10'b1100000111: data <= 11'h7fe; 
        10'b1100001000: data <= 11'h000; 
        10'b1100001001: data <= 11'h7ff; 
        10'b1100001010: data <= 11'h000; 
        10'b1100001011: data <= 11'h7fe; 
        10'b1100001100: data <= 11'h000; 
        10'b1100001101: data <= 11'h7ff; 
        10'b1100001110: data <= 11'h7fe; 
        10'b1100001111: data <= 11'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 6) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 12'hffe; 
        10'b0000000001: data <= 12'h000; 
        10'b0000000010: data <= 12'h000; 
        10'b0000000011: data <= 12'hffd; 
        10'b0000000100: data <= 12'hfff; 
        10'b0000000101: data <= 12'hffe; 
        10'b0000000110: data <= 12'h000; 
        10'b0000000111: data <= 12'hffe; 
        10'b0000001000: data <= 12'hfff; 
        10'b0000001001: data <= 12'h001; 
        10'b0000001010: data <= 12'hfff; 
        10'b0000001011: data <= 12'hfff; 
        10'b0000001100: data <= 12'hffe; 
        10'b0000001101: data <= 12'h000; 
        10'b0000001110: data <= 12'hffd; 
        10'b0000001111: data <= 12'hffe; 
        10'b0000010000: data <= 12'hffd; 
        10'b0000010001: data <= 12'hffd; 
        10'b0000010010: data <= 12'h000; 
        10'b0000010011: data <= 12'hfff; 
        10'b0000010100: data <= 12'hffd; 
        10'b0000010101: data <= 12'hfff; 
        10'b0000010110: data <= 12'hfff; 
        10'b0000010111: data <= 12'hffe; 
        10'b0000011000: data <= 12'hffd; 
        10'b0000011001: data <= 12'hfff; 
        10'b0000011010: data <= 12'hfff; 
        10'b0000011011: data <= 12'hffe; 
        10'b0000011100: data <= 12'h000; 
        10'b0000011101: data <= 12'hffc; 
        10'b0000011110: data <= 12'h000; 
        10'b0000011111: data <= 12'hffd; 
        10'b0000100000: data <= 12'h000; 
        10'b0000100001: data <= 12'hffe; 
        10'b0000100010: data <= 12'hfff; 
        10'b0000100011: data <= 12'hffe; 
        10'b0000100100: data <= 12'hffd; 
        10'b0000100101: data <= 12'hfff; 
        10'b0000100110: data <= 12'h000; 
        10'b0000100111: data <= 12'hffd; 
        10'b0000101000: data <= 12'hffe; 
        10'b0000101001: data <= 12'hffd; 
        10'b0000101010: data <= 12'hffd; 
        10'b0000101011: data <= 12'hfff; 
        10'b0000101100: data <= 12'hffe; 
        10'b0000101101: data <= 12'hffd; 
        10'b0000101110: data <= 12'hffe; 
        10'b0000101111: data <= 12'hffe; 
        10'b0000110000: data <= 12'hfff; 
        10'b0000110001: data <= 12'hffd; 
        10'b0000110010: data <= 12'h000; 
        10'b0000110011: data <= 12'hffd; 
        10'b0000110100: data <= 12'h000; 
        10'b0000110101: data <= 12'h000; 
        10'b0000110110: data <= 12'hffd; 
        10'b0000110111: data <= 12'hffe; 
        10'b0000111000: data <= 12'hffe; 
        10'b0000111001: data <= 12'hfff; 
        10'b0000111010: data <= 12'hffe; 
        10'b0000111011: data <= 12'hffd; 
        10'b0000111100: data <= 12'hffd; 
        10'b0000111101: data <= 12'hfff; 
        10'b0000111110: data <= 12'h000; 
        10'b0000111111: data <= 12'hfff; 
        10'b0001000000: data <= 12'hffd; 
        10'b0001000001: data <= 12'hffe; 
        10'b0001000010: data <= 12'h000; 
        10'b0001000011: data <= 12'hffc; 
        10'b0001000100: data <= 12'h000; 
        10'b0001000101: data <= 12'hffd; 
        10'b0001000110: data <= 12'hffd; 
        10'b0001000111: data <= 12'hffd; 
        10'b0001001000: data <= 12'hffe; 
        10'b0001001001: data <= 12'hfff; 
        10'b0001001010: data <= 12'hffe; 
        10'b0001001011: data <= 12'hffe; 
        10'b0001001100: data <= 12'h001; 
        10'b0001001101: data <= 12'h000; 
        10'b0001001110: data <= 12'h000; 
        10'b0001001111: data <= 12'hffd; 
        10'b0001010000: data <= 12'hffd; 
        10'b0001010001: data <= 12'hffe; 
        10'b0001010010: data <= 12'h000; 
        10'b0001010011: data <= 12'hfff; 
        10'b0001010100: data <= 12'hfff; 
        10'b0001010101: data <= 12'hfff; 
        10'b0001010110: data <= 12'hffd; 
        10'b0001010111: data <= 12'h000; 
        10'b0001011000: data <= 12'hffd; 
        10'b0001011001: data <= 12'hffe; 
        10'b0001011010: data <= 12'hffc; 
        10'b0001011011: data <= 12'hffe; 
        10'b0001011100: data <= 12'hffd; 
        10'b0001011101: data <= 12'hffe; 
        10'b0001011110: data <= 12'hffa; 
        10'b0001011111: data <= 12'hff8; 
        10'b0001100000: data <= 12'hffc; 
        10'b0001100001: data <= 12'hffc; 
        10'b0001100010: data <= 12'hffb; 
        10'b0001100011: data <= 12'hffe; 
        10'b0001100100: data <= 12'hfff; 
        10'b0001100101: data <= 12'hffc; 
        10'b0001100110: data <= 12'hffe; 
        10'b0001100111: data <= 12'hfff; 
        10'b0001101000: data <= 12'hfff; 
        10'b0001101001: data <= 12'hffe; 
        10'b0001101010: data <= 12'hffc; 
        10'b0001101011: data <= 12'hffd; 
        10'b0001101100: data <= 12'hffb; 
        10'b0001101101: data <= 12'h001; 
        10'b0001101110: data <= 12'h000; 
        10'b0001101111: data <= 12'hffd; 
        10'b0001110000: data <= 12'hffd; 
        10'b0001110001: data <= 12'hffe; 
        10'b0001110010: data <= 12'h000; 
        10'b0001110011: data <= 12'h000; 
        10'b0001110100: data <= 12'h000; 
        10'b0001110101: data <= 12'hffe; 
        10'b0001110110: data <= 12'hffd; 
        10'b0001110111: data <= 12'hffb; 
        10'b0001111000: data <= 12'hff7; 
        10'b0001111001: data <= 12'hff4; 
        10'b0001111010: data <= 12'hfee; 
        10'b0001111011: data <= 12'hff5; 
        10'b0001111100: data <= 12'hff5; 
        10'b0001111101: data <= 12'hff1; 
        10'b0001111110: data <= 12'hff8; 
        10'b0001111111: data <= 12'h000; 
        10'b0010000000: data <= 12'hfff; 
        10'b0010000001: data <= 12'h003; 
        10'b0010000010: data <= 12'hfff; 
        10'b0010000011: data <= 12'hffc; 
        10'b0010000100: data <= 12'hffa; 
        10'b0010000101: data <= 12'hffd; 
        10'b0010000110: data <= 12'hffe; 
        10'b0010000111: data <= 12'hffe; 
        10'b0010001000: data <= 12'hffe; 
        10'b0010001001: data <= 12'h001; 
        10'b0010001010: data <= 12'h000; 
        10'b0010001011: data <= 12'hffe; 
        10'b0010001100: data <= 12'hfff; 
        10'b0010001101: data <= 12'h001; 
        10'b0010001110: data <= 12'hffd; 
        10'b0010001111: data <= 12'hffd; 
        10'b0010010000: data <= 12'hffe; 
        10'b0010010001: data <= 12'hffa; 
        10'b0010010010: data <= 12'hff8; 
        10'b0010010011: data <= 12'hff8; 
        10'b0010010100: data <= 12'hffb; 
        10'b0010010101: data <= 12'hfff; 
        10'b0010010110: data <= 12'h002; 
        10'b0010010111: data <= 12'h002; 
        10'b0010011000: data <= 12'hffd; 
        10'b0010011001: data <= 12'hffc; 
        10'b0010011010: data <= 12'hffe; 
        10'b0010011011: data <= 12'hfff; 
        10'b0010011100: data <= 12'h004; 
        10'b0010011101: data <= 12'h004; 
        10'b0010011110: data <= 12'h008; 
        10'b0010011111: data <= 12'h005; 
        10'b0010100000: data <= 12'h005; 
        10'b0010100001: data <= 12'h006; 
        10'b0010100010: data <= 12'h00b; 
        10'b0010100011: data <= 12'h00a; 
        10'b0010100100: data <= 12'h007; 
        10'b0010100101: data <= 12'h004; 
        10'b0010100110: data <= 12'h002; 
        10'b0010100111: data <= 12'h001; 
        10'b0010101000: data <= 12'hffd; 
        10'b0010101001: data <= 12'hffd; 
        10'b0010101010: data <= 12'h000; 
        10'b0010101011: data <= 12'hffd; 
        10'b0010101100: data <= 12'hffc; 
        10'b0010101101: data <= 12'hff6; 
        10'b0010101110: data <= 12'hffc; 
        10'b0010101111: data <= 12'hfff; 
        10'b0010110000: data <= 12'h000; 
        10'b0010110001: data <= 12'h004; 
        10'b0010110010: data <= 12'h008; 
        10'b0010110011: data <= 12'h007; 
        10'b0010110100: data <= 12'h001; 
        10'b0010110101: data <= 12'h003; 
        10'b0010110110: data <= 12'hfff; 
        10'b0010110111: data <= 12'hffc; 
        10'b0010111000: data <= 12'hffe; 
        10'b0010111001: data <= 12'hffe; 
        10'b0010111010: data <= 12'h000; 
        10'b0010111011: data <= 12'h008; 
        10'b0010111100: data <= 12'h004; 
        10'b0010111101: data <= 12'h005; 
        10'b0010111110: data <= 12'h00f; 
        10'b0010111111: data <= 12'h013; 
        10'b0011000000: data <= 12'h015; 
        10'b0011000001: data <= 12'h00b; 
        10'b0011000010: data <= 12'h005; 
        10'b0011000011: data <= 12'h001; 
        10'b0011000100: data <= 12'hffe; 
        10'b0011000101: data <= 12'hfff; 
        10'b0011000110: data <= 12'hfff; 
        10'b0011000111: data <= 12'hffc; 
        10'b0011001000: data <= 12'hff5; 
        10'b0011001001: data <= 12'hff3; 
        10'b0011001010: data <= 12'hff8; 
        10'b0011001011: data <= 12'h001; 
        10'b0011001100: data <= 12'h005; 
        10'b0011001101: data <= 12'h00a; 
        10'b0011001110: data <= 12'h00a; 
        10'b0011001111: data <= 12'h009; 
        10'b0011010000: data <= 12'h003; 
        10'b0011010001: data <= 12'hfff; 
        10'b0011010010: data <= 12'hffd; 
        10'b0011010011: data <= 12'h000; 
        10'b0011010100: data <= 12'h004; 
        10'b0011010101: data <= 12'h004; 
        10'b0011010110: data <= 12'h005; 
        10'b0011010111: data <= 12'h00b; 
        10'b0011011000: data <= 12'h00a; 
        10'b0011011001: data <= 12'h00c; 
        10'b0011011010: data <= 12'h010; 
        10'b0011011011: data <= 12'h016; 
        10'b0011011100: data <= 12'h01b; 
        10'b0011011101: data <= 12'h013; 
        10'b0011011110: data <= 12'h003; 
        10'b0011011111: data <= 12'h000; 
        10'b0011100000: data <= 12'hfff; 
        10'b0011100001: data <= 12'h001; 
        10'b0011100010: data <= 12'h000; 
        10'b0011100011: data <= 12'hffb; 
        10'b0011100100: data <= 12'hff0; 
        10'b0011100101: data <= 12'hff2; 
        10'b0011100110: data <= 12'hff6; 
        10'b0011100111: data <= 12'h001; 
        10'b0011101000: data <= 12'h008; 
        10'b0011101001: data <= 12'h002; 
        10'b0011101010: data <= 12'h004; 
        10'b0011101011: data <= 12'h008; 
        10'b0011101100: data <= 12'h005; 
        10'b0011101101: data <= 12'hffa; 
        10'b0011101110: data <= 12'hff4; 
        10'b0011101111: data <= 12'hff9; 
        10'b0011110000: data <= 12'hffb; 
        10'b0011110001: data <= 12'h000; 
        10'b0011110010: data <= 12'h001; 
        10'b0011110011: data <= 12'h009; 
        10'b0011110100: data <= 12'h00a; 
        10'b0011110101: data <= 12'h00e; 
        10'b0011110110: data <= 12'h016; 
        10'b0011110111: data <= 12'h01d; 
        10'b0011111000: data <= 12'h027; 
        10'b0011111001: data <= 12'h019; 
        10'b0011111010: data <= 12'h005; 
        10'b0011111011: data <= 12'h000; 
        10'b0011111100: data <= 12'hffd; 
        10'b0011111101: data <= 12'hffe; 
        10'b0011111110: data <= 12'hffd; 
        10'b0011111111: data <= 12'hff8; 
        10'b0100000000: data <= 12'hff7; 
        10'b0100000001: data <= 12'hff8; 
        10'b0100000010: data <= 12'h001; 
        10'b0100000011: data <= 12'hfff; 
        10'b0100000100: data <= 12'h007; 
        10'b0100000101: data <= 12'h006; 
        10'b0100000110: data <= 12'h006; 
        10'b0100000111: data <= 12'h011; 
        10'b0100001000: data <= 12'h00b; 
        10'b0100001001: data <= 12'hffb; 
        10'b0100001010: data <= 12'hff1; 
        10'b0100001011: data <= 12'hfeb; 
        10'b0100001100: data <= 12'hfec; 
        10'b0100001101: data <= 12'hff4; 
        10'b0100001110: data <= 12'hffd; 
        10'b0100001111: data <= 12'h000; 
        10'b0100010000: data <= 12'h009; 
        10'b0100010001: data <= 12'h013; 
        10'b0100010010: data <= 12'h01c; 
        10'b0100010011: data <= 12'h026; 
        10'b0100010100: data <= 12'h030; 
        10'b0100010101: data <= 12'h020; 
        10'b0100010110: data <= 12'h006; 
        10'b0100010111: data <= 12'hffe; 
        10'b0100011000: data <= 12'hfff; 
        10'b0100011001: data <= 12'hffe; 
        10'b0100011010: data <= 12'hffd; 
        10'b0100011011: data <= 12'hffe; 
        10'b0100011100: data <= 12'hffd; 
        10'b0100011101: data <= 12'hffe; 
        10'b0100011110: data <= 12'h005; 
        10'b0100011111: data <= 12'h00a; 
        10'b0100100000: data <= 12'h010; 
        10'b0100100001: data <= 12'h011; 
        10'b0100100010: data <= 12'h011; 
        10'b0100100011: data <= 12'h014; 
        10'b0100100100: data <= 12'h011; 
        10'b0100100101: data <= 12'h00d; 
        10'b0100100110: data <= 12'hffd; 
        10'b0100100111: data <= 12'hff5; 
        10'b0100101000: data <= 12'hfee; 
        10'b0100101001: data <= 12'hfef; 
        10'b0100101010: data <= 12'hfee; 
        10'b0100101011: data <= 12'hfec; 
        10'b0100101100: data <= 12'hff2; 
        10'b0100101101: data <= 12'hffc; 
        10'b0100101110: data <= 12'h002; 
        10'b0100101111: data <= 12'h00d; 
        10'b0100110000: data <= 12'h01a; 
        10'b0100110001: data <= 12'h013; 
        10'b0100110010: data <= 12'h007; 
        10'b0100110011: data <= 12'hffe; 
        10'b0100110100: data <= 12'hffd; 
        10'b0100110101: data <= 12'h000; 
        10'b0100110110: data <= 12'hffe; 
        10'b0100110111: data <= 12'hffe; 
        10'b0100111000: data <= 12'hffe; 
        10'b0100111001: data <= 12'h000; 
        10'b0100111010: data <= 12'h009; 
        10'b0100111011: data <= 12'h00a; 
        10'b0100111100: data <= 12'h00f; 
        10'b0100111101: data <= 12'h00e; 
        10'b0100111110: data <= 12'h00a; 
        10'b0100111111: data <= 12'h00b; 
        10'b0101000000: data <= 12'h013; 
        10'b0101000001: data <= 12'h011; 
        10'b0101000010: data <= 12'h000; 
        10'b0101000011: data <= 12'hff5; 
        10'b0101000100: data <= 12'hff3; 
        10'b0101000101: data <= 12'hff1; 
        10'b0101000110: data <= 12'hfed; 
        10'b0101000111: data <= 12'hfe5; 
        10'b0101001000: data <= 12'hfd9; 
        10'b0101001001: data <= 12'hfdc; 
        10'b0101001010: data <= 12'hfe2; 
        10'b0101001011: data <= 12'hfea; 
        10'b0101001100: data <= 12'hff8; 
        10'b0101001101: data <= 12'h001; 
        10'b0101001110: data <= 12'h002; 
        10'b0101001111: data <= 12'hfff; 
        10'b0101010000: data <= 12'hfff; 
        10'b0101010001: data <= 12'hfff; 
        10'b0101010010: data <= 12'hffe; 
        10'b0101010011: data <= 12'hffe; 
        10'b0101010100: data <= 12'hffe; 
        10'b0101010101: data <= 12'h004; 
        10'b0101010110: data <= 12'h00a; 
        10'b0101010111: data <= 12'h009; 
        10'b0101011000: data <= 12'h006; 
        10'b0101011001: data <= 12'h004; 
        10'b0101011010: data <= 12'h00b; 
        10'b0101011011: data <= 12'h017; 
        10'b0101011100: data <= 12'h015; 
        10'b0101011101: data <= 12'h016; 
        10'b0101011110: data <= 12'h002; 
        10'b0101011111: data <= 12'hff5; 
        10'b0101100000: data <= 12'hfec; 
        10'b0101100001: data <= 12'hfef; 
        10'b0101100010: data <= 12'hff5; 
        10'b0101100011: data <= 12'hff0; 
        10'b0101100100: data <= 12'hfee; 
        10'b0101100101: data <= 12'hfe2; 
        10'b0101100110: data <= 12'hfdd; 
        10'b0101100111: data <= 12'hfe2; 
        10'b0101101000: data <= 12'hfec; 
        10'b0101101001: data <= 12'hffa; 
        10'b0101101010: data <= 12'h000; 
        10'b0101101011: data <= 12'h000; 
        10'b0101101100: data <= 12'hfff; 
        10'b0101101101: data <= 12'hffd; 
        10'b0101101110: data <= 12'hffd; 
        10'b0101101111: data <= 12'hffe; 
        10'b0101110000: data <= 12'hfff; 
        10'b0101110001: data <= 12'h002; 
        10'b0101110010: data <= 12'h007; 
        10'b0101110011: data <= 12'h005; 
        10'b0101110100: data <= 12'h006; 
        10'b0101110101: data <= 12'h005; 
        10'b0101110110: data <= 12'h00f; 
        10'b0101110111: data <= 12'h011; 
        10'b0101111000: data <= 12'h00d; 
        10'b0101111001: data <= 12'h00c; 
        10'b0101111010: data <= 12'hffe; 
        10'b0101111011: data <= 12'hff3; 
        10'b0101111100: data <= 12'hfeb; 
        10'b0101111101: data <= 12'hff5; 
        10'b0101111110: data <= 12'hffc; 
        10'b0101111111: data <= 12'hffb; 
        10'b0110000000: data <= 12'hffe; 
        10'b0110000001: data <= 12'hff7; 
        10'b0110000010: data <= 12'hff0; 
        10'b0110000011: data <= 12'hfe9; 
        10'b0110000100: data <= 12'hfef; 
        10'b0110000101: data <= 12'hffd; 
        10'b0110000110: data <= 12'hffd; 
        10'b0110000111: data <= 12'h000; 
        10'b0110001000: data <= 12'hfff; 
        10'b0110001001: data <= 12'hffd; 
        10'b0110001010: data <= 12'hffe; 
        10'b0110001011: data <= 12'hffc; 
        10'b0110001100: data <= 12'hfff; 
        10'b0110001101: data <= 12'hfff; 
        10'b0110001110: data <= 12'h000; 
        10'b0110001111: data <= 12'hfff; 
        10'b0110010000: data <= 12'h007; 
        10'b0110010001: data <= 12'h00b; 
        10'b0110010010: data <= 12'h00d; 
        10'b0110010011: data <= 12'h003; 
        10'b0110010100: data <= 12'h004; 
        10'b0110010101: data <= 12'hfff; 
        10'b0110010110: data <= 12'hff6; 
        10'b0110010111: data <= 12'hff5; 
        10'b0110011000: data <= 12'hff1; 
        10'b0110011001: data <= 12'hff3; 
        10'b0110011010: data <= 12'hff3; 
        10'b0110011011: data <= 12'hffa; 
        10'b0110011100: data <= 12'hffb; 
        10'b0110011101: data <= 12'hffb; 
        10'b0110011110: data <= 12'hffd; 
        10'b0110011111: data <= 12'hff3; 
        10'b0110100000: data <= 12'hff8; 
        10'b0110100001: data <= 12'hffc; 
        10'b0110100010: data <= 12'hffe; 
        10'b0110100011: data <= 12'hffc; 
        10'b0110100100: data <= 12'hffd; 
        10'b0110100101: data <= 12'h001; 
        10'b0110100110: data <= 12'hffc; 
        10'b0110100111: data <= 12'hfff; 
        10'b0110101000: data <= 12'hffb; 
        10'b0110101001: data <= 12'hff8; 
        10'b0110101010: data <= 12'hff5; 
        10'b0110101011: data <= 12'hff9; 
        10'b0110101100: data <= 12'h003; 
        10'b0110101101: data <= 12'h00c; 
        10'b0110101110: data <= 12'h006; 
        10'b0110101111: data <= 12'h005; 
        10'b0110110000: data <= 12'h005; 
        10'b0110110001: data <= 12'hffc; 
        10'b0110110010: data <= 12'hff2; 
        10'b0110110011: data <= 12'hff0; 
        10'b0110110100: data <= 12'hff1; 
        10'b0110110101: data <= 12'hff1; 
        10'b0110110110: data <= 12'hff5; 
        10'b0110110111: data <= 12'hfff; 
        10'b0110111000: data <= 12'hffc; 
        10'b0110111001: data <= 12'hffd; 
        10'b0110111010: data <= 12'hffc; 
        10'b0110111011: data <= 12'hffc; 
        10'b0110111100: data <= 12'hffd; 
        10'b0110111101: data <= 12'h000; 
        10'b0110111110: data <= 12'h001; 
        10'b0110111111: data <= 12'hffe; 
        10'b0111000000: data <= 12'hffe; 
        10'b0111000001: data <= 12'hfff; 
        10'b0111000010: data <= 12'hfff; 
        10'b0111000011: data <= 12'hffc; 
        10'b0111000100: data <= 12'hffe; 
        10'b0111000101: data <= 12'hff7; 
        10'b0111000110: data <= 12'hfee; 
        10'b0111000111: data <= 12'hfea; 
        10'b0111001000: data <= 12'hff1; 
        10'b0111001001: data <= 12'hff8; 
        10'b0111001010: data <= 12'hffd; 
        10'b0111001011: data <= 12'hffb; 
        10'b0111001100: data <= 12'hffd; 
        10'b0111001101: data <= 12'hff6; 
        10'b0111001110: data <= 12'hfed; 
        10'b0111001111: data <= 12'hff0; 
        10'b0111010000: data <= 12'hff5; 
        10'b0111010001: data <= 12'hffc; 
        10'b0111010010: data <= 12'hffc; 
        10'b0111010011: data <= 12'h001; 
        10'b0111010100: data <= 12'h003; 
        10'b0111010101: data <= 12'h001; 
        10'b0111010110: data <= 12'h003; 
        10'b0111010111: data <= 12'h001; 
        10'b0111011000: data <= 12'h001; 
        10'b0111011001: data <= 12'h000; 
        10'b0111011010: data <= 12'hffe; 
        10'b0111011011: data <= 12'hffe; 
        10'b0111011100: data <= 12'hffe; 
        10'b0111011101: data <= 12'h000; 
        10'b0111011110: data <= 12'h000; 
        10'b0111011111: data <= 12'h000; 
        10'b0111100000: data <= 12'hffe; 
        10'b0111100001: data <= 12'h001; 
        10'b0111100010: data <= 12'h001; 
        10'b0111100011: data <= 12'hff2; 
        10'b0111100100: data <= 12'hfe6; 
        10'b0111100101: data <= 12'hfe8; 
        10'b0111100110: data <= 12'hfef; 
        10'b0111100111: data <= 12'hff6; 
        10'b0111101000: data <= 12'hff0; 
        10'b0111101001: data <= 12'hfeb; 
        10'b0111101010: data <= 12'hfeb; 
        10'b0111101011: data <= 12'hff7; 
        10'b0111101100: data <= 12'hffc; 
        10'b0111101101: data <= 12'h006; 
        10'b0111101110: data <= 12'h009; 
        10'b0111101111: data <= 12'h006; 
        10'b0111110000: data <= 12'h006; 
        10'b0111110001: data <= 12'h002; 
        10'b0111110010: data <= 12'h000; 
        10'b0111110011: data <= 12'h003; 
        10'b0111110100: data <= 12'h004; 
        10'b0111110101: data <= 12'hffd; 
        10'b0111110110: data <= 12'h000; 
        10'b0111110111: data <= 12'h000; 
        10'b0111111000: data <= 12'h000; 
        10'b0111111001: data <= 12'hffd; 
        10'b0111111010: data <= 12'hffe; 
        10'b0111111011: data <= 12'hffe; 
        10'b0111111100: data <= 12'h005; 
        10'b0111111101: data <= 12'h007; 
        10'b0111111110: data <= 12'h010; 
        10'b0111111111: data <= 12'h003; 
        10'b1000000000: data <= 12'hff0; 
        10'b1000000001: data <= 12'hfe9; 
        10'b1000000010: data <= 12'hfe2; 
        10'b1000000011: data <= 12'hfe5; 
        10'b1000000100: data <= 12'hfed; 
        10'b1000000101: data <= 12'hff5; 
        10'b1000000110: data <= 12'hffb; 
        10'b1000000111: data <= 12'hffe; 
        10'b1000001000: data <= 12'h000; 
        10'b1000001001: data <= 12'h007; 
        10'b1000001010: data <= 12'h004; 
        10'b1000001011: data <= 12'h006; 
        10'b1000001100: data <= 12'h004; 
        10'b1000001101: data <= 12'h006; 
        10'b1000001110: data <= 12'h005; 
        10'b1000001111: data <= 12'h007; 
        10'b1000010000: data <= 12'h004; 
        10'b1000010001: data <= 12'h000; 
        10'b1000010010: data <= 12'hffd; 
        10'b1000010011: data <= 12'hfff; 
        10'b1000010100: data <= 12'h000; 
        10'b1000010101: data <= 12'hffd; 
        10'b1000010110: data <= 12'hfff; 
        10'b1000010111: data <= 12'h001; 
        10'b1000011000: data <= 12'h008; 
        10'b1000011001: data <= 12'h00d; 
        10'b1000011010: data <= 12'h012; 
        10'b1000011011: data <= 12'h00c; 
        10'b1000011100: data <= 12'h008; 
        10'b1000011101: data <= 12'h002; 
        10'b1000011110: data <= 12'hffa; 
        10'b1000011111: data <= 12'hffa; 
        10'b1000100000: data <= 12'h001; 
        10'b1000100001: data <= 12'h007; 
        10'b1000100010: data <= 12'h003; 
        10'b1000100011: data <= 12'h004; 
        10'b1000100100: data <= 12'h004; 
        10'b1000100101: data <= 12'hfff; 
        10'b1000100110: data <= 12'h003; 
        10'b1000100111: data <= 12'h003; 
        10'b1000101000: data <= 12'h001; 
        10'b1000101001: data <= 12'h005; 
        10'b1000101010: data <= 12'h008; 
        10'b1000101011: data <= 12'h006; 
        10'b1000101100: data <= 12'h000; 
        10'b1000101101: data <= 12'h000; 
        10'b1000101110: data <= 12'h000; 
        10'b1000101111: data <= 12'hffd; 
        10'b1000110000: data <= 12'h000; 
        10'b1000110001: data <= 12'hffc; 
        10'b1000110010: data <= 12'hffe; 
        10'b1000110011: data <= 12'hffd; 
        10'b1000110100: data <= 12'h001; 
        10'b1000110101: data <= 12'h009; 
        10'b1000110110: data <= 12'h00a; 
        10'b1000110111: data <= 12'h00c; 
        10'b1000111000: data <= 12'h011; 
        10'b1000111001: data <= 12'h00f; 
        10'b1000111010: data <= 12'h00d; 
        10'b1000111011: data <= 12'h013; 
        10'b1000111100: data <= 12'h00c; 
        10'b1000111101: data <= 12'h009; 
        10'b1000111110: data <= 12'hffe; 
        10'b1000111111: data <= 12'hffe; 
        10'b1001000000: data <= 12'h006; 
        10'b1001000001: data <= 12'h003; 
        10'b1001000010: data <= 12'h005; 
        10'b1001000011: data <= 12'h007; 
        10'b1001000100: data <= 12'h006; 
        10'b1001000101: data <= 12'h005; 
        10'b1001000110: data <= 12'h00c; 
        10'b1001000111: data <= 12'h009; 
        10'b1001001000: data <= 12'hfff; 
        10'b1001001001: data <= 12'hffc; 
        10'b1001001010: data <= 12'hfff; 
        10'b1001001011: data <= 12'hffe; 
        10'b1001001100: data <= 12'hffd; 
        10'b1001001101: data <= 12'h000; 
        10'b1001001110: data <= 12'hffc; 
        10'b1001001111: data <= 12'hfff; 
        10'b1001010000: data <= 12'h003; 
        10'b1001010001: data <= 12'hfff; 
        10'b1001010010: data <= 12'h004; 
        10'b1001010011: data <= 12'h00b; 
        10'b1001010100: data <= 12'h010; 
        10'b1001010101: data <= 12'h00b; 
        10'b1001010110: data <= 12'h009; 
        10'b1001010111: data <= 12'h005; 
        10'b1001011000: data <= 12'h006; 
        10'b1001011001: data <= 12'h004; 
        10'b1001011010: data <= 12'h004; 
        10'b1001011011: data <= 12'h005; 
        10'b1001011100: data <= 12'h001; 
        10'b1001011101: data <= 12'h004; 
        10'b1001011110: data <= 12'h002; 
        10'b1001011111: data <= 12'h006; 
        10'b1001100000: data <= 12'h006; 
        10'b1001100001: data <= 12'h00b; 
        10'b1001100010: data <= 12'h00d; 
        10'b1001100011: data <= 12'h003; 
        10'b1001100100: data <= 12'h000; 
        10'b1001100101: data <= 12'hffd; 
        10'b1001100110: data <= 12'hffe; 
        10'b1001100111: data <= 12'hffe; 
        10'b1001101000: data <= 12'hfff; 
        10'b1001101001: data <= 12'hffc; 
        10'b1001101010: data <= 12'hffe; 
        10'b1001101011: data <= 12'hffe; 
        10'b1001101100: data <= 12'h001; 
        10'b1001101101: data <= 12'hffe; 
        10'b1001101110: data <= 12'hffc; 
        10'b1001101111: data <= 12'hfff; 
        10'b1001110000: data <= 12'h006; 
        10'b1001110001: data <= 12'h009; 
        10'b1001110010: data <= 12'h002; 
        10'b1001110011: data <= 12'h008; 
        10'b1001110100: data <= 12'h00d; 
        10'b1001110101: data <= 12'h010; 
        10'b1001110110: data <= 12'h008; 
        10'b1001110111: data <= 12'h001; 
        10'b1001111000: data <= 12'h001; 
        10'b1001111001: data <= 12'h002; 
        10'b1001111010: data <= 12'h004; 
        10'b1001111011: data <= 12'h004; 
        10'b1001111100: data <= 12'h007; 
        10'b1001111101: data <= 12'h007; 
        10'b1001111110: data <= 12'h007; 
        10'b1001111111: data <= 12'h002; 
        10'b1010000000: data <= 12'h000; 
        10'b1010000001: data <= 12'h000; 
        10'b1010000010: data <= 12'hfff; 
        10'b1010000011: data <= 12'hfff; 
        10'b1010000100: data <= 12'hffd; 
        10'b1010000101: data <= 12'hfff; 
        10'b1010000110: data <= 12'hfff; 
        10'b1010000111: data <= 12'hfff; 
        10'b1010001000: data <= 12'hffd; 
        10'b1010001001: data <= 12'hffe; 
        10'b1010001010: data <= 12'hffa; 
        10'b1010001011: data <= 12'hffd; 
        10'b1010001100: data <= 12'h005; 
        10'b1010001101: data <= 12'h005; 
        10'b1010001110: data <= 12'h005; 
        10'b1010001111: data <= 12'h009; 
        10'b1010010000: data <= 12'h008; 
        10'b1010010001: data <= 12'h006; 
        10'b1010010010: data <= 12'h007; 
        10'b1010010011: data <= 12'h006; 
        10'b1010010100: data <= 12'h006; 
        10'b1010010101: data <= 12'h003; 
        10'b1010010110: data <= 12'hffd; 
        10'b1010010111: data <= 12'h000; 
        10'b1010011000: data <= 12'h003; 
        10'b1010011001: data <= 12'h001; 
        10'b1010011010: data <= 12'h004; 
        10'b1010011011: data <= 12'hffe; 
        10'b1010011100: data <= 12'h001; 
        10'b1010011101: data <= 12'hffe; 
        10'b1010011110: data <= 12'hffe; 
        10'b1010011111: data <= 12'h001; 
        10'b1010100000: data <= 12'h000; 
        10'b1010100001: data <= 12'hffe; 
        10'b1010100010: data <= 12'hffe; 
        10'b1010100011: data <= 12'h001; 
        10'b1010100100: data <= 12'hffc; 
        10'b1010100101: data <= 12'hffc; 
        10'b1010100110: data <= 12'hfff; 
        10'b1010100111: data <= 12'hfff; 
        10'b1010101000: data <= 12'h000; 
        10'b1010101001: data <= 12'h007; 
        10'b1010101010: data <= 12'h008; 
        10'b1010101011: data <= 12'h007; 
        10'b1010101100: data <= 12'h004; 
        10'b1010101101: data <= 12'h006; 
        10'b1010101110: data <= 12'h00b; 
        10'b1010101111: data <= 12'h009; 
        10'b1010110000: data <= 12'h005; 
        10'b1010110001: data <= 12'h003; 
        10'b1010110010: data <= 12'h005; 
        10'b1010110011: data <= 12'h003; 
        10'b1010110100: data <= 12'h000; 
        10'b1010110101: data <= 12'h000; 
        10'b1010110110: data <= 12'hfff; 
        10'b1010110111: data <= 12'h000; 
        10'b1010111000: data <= 12'hffd; 
        10'b1010111001: data <= 12'hfff; 
        10'b1010111010: data <= 12'h000; 
        10'b1010111011: data <= 12'hffd; 
        10'b1010111100: data <= 12'hfff; 
        10'b1010111101: data <= 12'h000; 
        10'b1010111110: data <= 12'h000; 
        10'b1010111111: data <= 12'hffd; 
        10'b1011000000: data <= 12'h000; 
        10'b1011000001: data <= 12'hfff; 
        10'b1011000010: data <= 12'hffc; 
        10'b1011000011: data <= 12'hfff; 
        10'b1011000100: data <= 12'hffc; 
        10'b1011000101: data <= 12'h002; 
        10'b1011000110: data <= 12'h002; 
        10'b1011000111: data <= 12'h004; 
        10'b1011001000: data <= 12'h004; 
        10'b1011001001: data <= 12'h008; 
        10'b1011001010: data <= 12'h000; 
        10'b1011001011: data <= 12'h002; 
        10'b1011001100: data <= 12'h002; 
        10'b1011001101: data <= 12'h004; 
        10'b1011001110: data <= 12'hffd; 
        10'b1011001111: data <= 12'h000; 
        10'b1011010000: data <= 12'hffc; 
        10'b1011010001: data <= 12'h000; 
        10'b1011010010: data <= 12'hffe; 
        10'b1011010011: data <= 12'hffd; 
        10'b1011010100: data <= 12'h000; 
        10'b1011010101: data <= 12'h000; 
        10'b1011010110: data <= 12'hffc; 
        10'b1011010111: data <= 12'hffe; 
        10'b1011011000: data <= 12'hfff; 
        10'b1011011001: data <= 12'hfff; 
        10'b1011011010: data <= 12'hffd; 
        10'b1011011011: data <= 12'hffe; 
        10'b1011011100: data <= 12'hffe; 
        10'b1011011101: data <= 12'hffe; 
        10'b1011011110: data <= 12'hfff; 
        10'b1011011111: data <= 12'hffd; 
        10'b1011100000: data <= 12'hffd; 
        10'b1011100001: data <= 12'hffe; 
        10'b1011100010: data <= 12'hffe; 
        10'b1011100011: data <= 12'h000; 
        10'b1011100100: data <= 12'h000; 
        10'b1011100101: data <= 12'hfff; 
        10'b1011100110: data <= 12'hffd; 
        10'b1011100111: data <= 12'hfff; 
        10'b1011101000: data <= 12'hfff; 
        10'b1011101001: data <= 12'hffd; 
        10'b1011101010: data <= 12'hffb; 
        10'b1011101011: data <= 12'hffc; 
        10'b1011101100: data <= 12'hfff; 
        10'b1011101101: data <= 12'hfff; 
        10'b1011101110: data <= 12'hffe; 
        10'b1011101111: data <= 12'hfff; 
        10'b1011110000: data <= 12'hffe; 
        10'b1011110001: data <= 12'hfff; 
        10'b1011110010: data <= 12'hffe; 
        10'b1011110011: data <= 12'hffc; 
        10'b1011110100: data <= 12'hfff; 
        10'b1011110101: data <= 12'h000; 
        10'b1011110110: data <= 12'h000; 
        10'b1011110111: data <= 12'hfff; 
        10'b1011111000: data <= 12'hffd; 
        10'b1011111001: data <= 12'h000; 
        10'b1011111010: data <= 12'hffe; 
        10'b1011111011: data <= 12'hffe; 
        10'b1011111100: data <= 12'h001; 
        10'b1011111101: data <= 12'hffe; 
        10'b1011111110: data <= 12'hffe; 
        10'b1011111111: data <= 12'h000; 
        10'b1100000000: data <= 12'hfff; 
        10'b1100000001: data <= 12'hffc; 
        10'b1100000010: data <= 12'h000; 
        10'b1100000011: data <= 12'hfff; 
        10'b1100000100: data <= 12'hffd; 
        10'b1100000101: data <= 12'hffc; 
        10'b1100000110: data <= 12'hffd; 
        10'b1100000111: data <= 12'hffc; 
        10'b1100001000: data <= 12'h000; 
        10'b1100001001: data <= 12'hffe; 
        10'b1100001010: data <= 12'h001; 
        10'b1100001011: data <= 12'hffd; 
        10'b1100001100: data <= 12'hfff; 
        10'b1100001101: data <= 12'hffe; 
        10'b1100001110: data <= 12'hffd; 
        10'b1100001111: data <= 12'h000; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 7) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 13'h1ffc; 
        10'b0000000001: data <= 13'h1fff; 
        10'b0000000010: data <= 13'h1fff; 
        10'b0000000011: data <= 13'h1ffa; 
        10'b0000000100: data <= 13'h1ffd; 
        10'b0000000101: data <= 13'h1ffc; 
        10'b0000000110: data <= 13'h0000; 
        10'b0000000111: data <= 13'h1ffc; 
        10'b0000001000: data <= 13'h1ffe; 
        10'b0000001001: data <= 13'h0001; 
        10'b0000001010: data <= 13'h1ffe; 
        10'b0000001011: data <= 13'h1ffe; 
        10'b0000001100: data <= 13'h1ffb; 
        10'b0000001101: data <= 13'h0000; 
        10'b0000001110: data <= 13'h1ffa; 
        10'b0000001111: data <= 13'h1ffb; 
        10'b0000010000: data <= 13'h1ff9; 
        10'b0000010001: data <= 13'h1ffa; 
        10'b0000010010: data <= 13'h1fff; 
        10'b0000010011: data <= 13'h1ffe; 
        10'b0000010100: data <= 13'h1ff9; 
        10'b0000010101: data <= 13'h1ffd; 
        10'b0000010110: data <= 13'h1ffe; 
        10'b0000010111: data <= 13'h1ffd; 
        10'b0000011000: data <= 13'h1ff9; 
        10'b0000011001: data <= 13'h1ffe; 
        10'b0000011010: data <= 13'h1ffe; 
        10'b0000011011: data <= 13'h1ffc; 
        10'b0000011100: data <= 13'h0000; 
        10'b0000011101: data <= 13'h1ff9; 
        10'b0000011110: data <= 13'h0000; 
        10'b0000011111: data <= 13'h1ffa; 
        10'b0000100000: data <= 13'h0000; 
        10'b0000100001: data <= 13'h1ffc; 
        10'b0000100010: data <= 13'h1ffe; 
        10'b0000100011: data <= 13'h1ffc; 
        10'b0000100100: data <= 13'h1ffb; 
        10'b0000100101: data <= 13'h1ffe; 
        10'b0000100110: data <= 13'h0001; 
        10'b0000100111: data <= 13'h1ffa; 
        10'b0000101000: data <= 13'h1ffc; 
        10'b0000101001: data <= 13'h1ffb; 
        10'b0000101010: data <= 13'h1ff9; 
        10'b0000101011: data <= 13'h1fff; 
        10'b0000101100: data <= 13'h1ffb; 
        10'b0000101101: data <= 13'h1ffa; 
        10'b0000101110: data <= 13'h1ffb; 
        10'b0000101111: data <= 13'h1ffb; 
        10'b0000110000: data <= 13'h1ffe; 
        10'b0000110001: data <= 13'h1ffa; 
        10'b0000110010: data <= 13'h0000; 
        10'b0000110011: data <= 13'h1ffa; 
        10'b0000110100: data <= 13'h0000; 
        10'b0000110101: data <= 13'h0000; 
        10'b0000110110: data <= 13'h1ffa; 
        10'b0000110111: data <= 13'h1ffd; 
        10'b0000111000: data <= 13'h1ffd; 
        10'b0000111001: data <= 13'h1fff; 
        10'b0000111010: data <= 13'h1ffc; 
        10'b0000111011: data <= 13'h1ff9; 
        10'b0000111100: data <= 13'h1ffa; 
        10'b0000111101: data <= 13'h1ffe; 
        10'b0000111110: data <= 13'h0000; 
        10'b0000111111: data <= 13'h1ffe; 
        10'b0001000000: data <= 13'h1ffb; 
        10'b0001000001: data <= 13'h1ffc; 
        10'b0001000010: data <= 13'h0001; 
        10'b0001000011: data <= 13'h1ff9; 
        10'b0001000100: data <= 13'h0000; 
        10'b0001000101: data <= 13'h1ffb; 
        10'b0001000110: data <= 13'h1ff9; 
        10'b0001000111: data <= 13'h1ffa; 
        10'b0001001000: data <= 13'h1ffc; 
        10'b0001001001: data <= 13'h1ffd; 
        10'b0001001010: data <= 13'h1ffc; 
        10'b0001001011: data <= 13'h1ffc; 
        10'b0001001100: data <= 13'h0002; 
        10'b0001001101: data <= 13'h0000; 
        10'b0001001110: data <= 13'h0001; 
        10'b0001001111: data <= 13'h1ffb; 
        10'b0001010000: data <= 13'h1ff9; 
        10'b0001010001: data <= 13'h1ffd; 
        10'b0001010010: data <= 13'h0000; 
        10'b0001010011: data <= 13'h1ffe; 
        10'b0001010100: data <= 13'h1fff; 
        10'b0001010101: data <= 13'h1ffe; 
        10'b0001010110: data <= 13'h1ffa; 
        10'b0001010111: data <= 13'h0000; 
        10'b0001011000: data <= 13'h1ffa; 
        10'b0001011001: data <= 13'h1ffc; 
        10'b0001011010: data <= 13'h1ff9; 
        10'b0001011011: data <= 13'h1ffb; 
        10'b0001011100: data <= 13'h1ff9; 
        10'b0001011101: data <= 13'h1ffb; 
        10'b0001011110: data <= 13'h1ff4; 
        10'b0001011111: data <= 13'h1ff1; 
        10'b0001100000: data <= 13'h1ff7; 
        10'b0001100001: data <= 13'h1ff8; 
        10'b0001100010: data <= 13'h1ff6; 
        10'b0001100011: data <= 13'h1ffd; 
        10'b0001100100: data <= 13'h1fff; 
        10'b0001100101: data <= 13'h1ff8; 
        10'b0001100110: data <= 13'h1ffb; 
        10'b0001100111: data <= 13'h1fff; 
        10'b0001101000: data <= 13'h1fff; 
        10'b0001101001: data <= 13'h1ffd; 
        10'b0001101010: data <= 13'h1ff8; 
        10'b0001101011: data <= 13'h1ffb; 
        10'b0001101100: data <= 13'h1ff6; 
        10'b0001101101: data <= 13'h0001; 
        10'b0001101110: data <= 13'h0001; 
        10'b0001101111: data <= 13'h1ffa; 
        10'b0001110000: data <= 13'h1ff9; 
        10'b0001110001: data <= 13'h1ffc; 
        10'b0001110010: data <= 13'h0001; 
        10'b0001110011: data <= 13'h0000; 
        10'b0001110100: data <= 13'h0001; 
        10'b0001110101: data <= 13'h1ffb; 
        10'b0001110110: data <= 13'h1ffb; 
        10'b0001110111: data <= 13'h1ff5; 
        10'b0001111000: data <= 13'h1fee; 
        10'b0001111001: data <= 13'h1fe8; 
        10'b0001111010: data <= 13'h1fdd; 
        10'b0001111011: data <= 13'h1fe9; 
        10'b0001111100: data <= 13'h1fe9; 
        10'b0001111101: data <= 13'h1fe1; 
        10'b0001111110: data <= 13'h1fef; 
        10'b0001111111: data <= 13'h0000; 
        10'b0010000000: data <= 13'h1ffe; 
        10'b0010000001: data <= 13'h0006; 
        10'b0010000010: data <= 13'h1ffe; 
        10'b0010000011: data <= 13'h1ff7; 
        10'b0010000100: data <= 13'h1ff5; 
        10'b0010000101: data <= 13'h1ffa; 
        10'b0010000110: data <= 13'h1ffb; 
        10'b0010000111: data <= 13'h1ffd; 
        10'b0010001000: data <= 13'h1ffc; 
        10'b0010001001: data <= 13'h0002; 
        10'b0010001010: data <= 13'h0001; 
        10'b0010001011: data <= 13'h1ffd; 
        10'b0010001100: data <= 13'h1ffd; 
        10'b0010001101: data <= 13'h0002; 
        10'b0010001110: data <= 13'h1ffb; 
        10'b0010001111: data <= 13'h1ffa; 
        10'b0010010000: data <= 13'h1ffb; 
        10'b0010010001: data <= 13'h1ff5; 
        10'b0010010010: data <= 13'h1fef; 
        10'b0010010011: data <= 13'h1ff0; 
        10'b0010010100: data <= 13'h1ff5; 
        10'b0010010101: data <= 13'h1ffe; 
        10'b0010010110: data <= 13'h0004; 
        10'b0010010111: data <= 13'h0004; 
        10'b0010011000: data <= 13'h1ffa; 
        10'b0010011001: data <= 13'h1ff8; 
        10'b0010011010: data <= 13'h1ffb; 
        10'b0010011011: data <= 13'h1ffe; 
        10'b0010011100: data <= 13'h0008; 
        10'b0010011101: data <= 13'h0008; 
        10'b0010011110: data <= 13'h0010; 
        10'b0010011111: data <= 13'h000a; 
        10'b0010100000: data <= 13'h000a; 
        10'b0010100001: data <= 13'h000c; 
        10'b0010100010: data <= 13'h0017; 
        10'b0010100011: data <= 13'h0013; 
        10'b0010100100: data <= 13'h000e; 
        10'b0010100101: data <= 13'h0007; 
        10'b0010100110: data <= 13'h0005; 
        10'b0010100111: data <= 13'h0002; 
        10'b0010101000: data <= 13'h1ffa; 
        10'b0010101001: data <= 13'h1ff9; 
        10'b0010101010: data <= 13'h0001; 
        10'b0010101011: data <= 13'h1ffa; 
        10'b0010101100: data <= 13'h1ff8; 
        10'b0010101101: data <= 13'h1fed; 
        10'b0010101110: data <= 13'h1ff7; 
        10'b0010101111: data <= 13'h1fff; 
        10'b0010110000: data <= 13'h1fff; 
        10'b0010110001: data <= 13'h0008; 
        10'b0010110010: data <= 13'h0010; 
        10'b0010110011: data <= 13'h000e; 
        10'b0010110100: data <= 13'h0002; 
        10'b0010110101: data <= 13'h0005; 
        10'b0010110110: data <= 13'h1ffe; 
        10'b0010110111: data <= 13'h1ff8; 
        10'b0010111000: data <= 13'h1ffb; 
        10'b0010111001: data <= 13'h1ffc; 
        10'b0010111010: data <= 13'h0000; 
        10'b0010111011: data <= 13'h0010; 
        10'b0010111100: data <= 13'h0009; 
        10'b0010111101: data <= 13'h000a; 
        10'b0010111110: data <= 13'h001f; 
        10'b0010111111: data <= 13'h0025; 
        10'b0011000000: data <= 13'h002a; 
        10'b0011000001: data <= 13'h0016; 
        10'b0011000010: data <= 13'h000b; 
        10'b0011000011: data <= 13'h0003; 
        10'b0011000100: data <= 13'h1ffd; 
        10'b0011000101: data <= 13'h1ffe; 
        10'b0011000110: data <= 13'h1ffd; 
        10'b0011000111: data <= 13'h1ff8; 
        10'b0011001000: data <= 13'h1fe9; 
        10'b0011001001: data <= 13'h1fe5; 
        10'b0011001010: data <= 13'h1ff0; 
        10'b0011001011: data <= 13'h0002; 
        10'b0011001100: data <= 13'h000b; 
        10'b0011001101: data <= 13'h0015; 
        10'b0011001110: data <= 13'h0014; 
        10'b0011001111: data <= 13'h0012; 
        10'b0011010000: data <= 13'h0005; 
        10'b0011010001: data <= 13'h1ffe; 
        10'b0011010010: data <= 13'h1ffa; 
        10'b0011010011: data <= 13'h0000; 
        10'b0011010100: data <= 13'h0009; 
        10'b0011010101: data <= 13'h0008; 
        10'b0011010110: data <= 13'h000a; 
        10'b0011010111: data <= 13'h0016; 
        10'b0011011000: data <= 13'h0013; 
        10'b0011011001: data <= 13'h0017; 
        10'b0011011010: data <= 13'h0020; 
        10'b0011011011: data <= 13'h002b; 
        10'b0011011100: data <= 13'h0035; 
        10'b0011011101: data <= 13'h0026; 
        10'b0011011110: data <= 13'h0006; 
        10'b0011011111: data <= 13'h1fff; 
        10'b0011100000: data <= 13'h1ffe; 
        10'b0011100001: data <= 13'h0001; 
        10'b0011100010: data <= 13'h0000; 
        10'b0011100011: data <= 13'h1ff5; 
        10'b0011100100: data <= 13'h1fdf; 
        10'b0011100101: data <= 13'h1fe4; 
        10'b0011100110: data <= 13'h1fec; 
        10'b0011100111: data <= 13'h0001; 
        10'b0011101000: data <= 13'h0010; 
        10'b0011101001: data <= 13'h0005; 
        10'b0011101010: data <= 13'h0008; 
        10'b0011101011: data <= 13'h0010; 
        10'b0011101100: data <= 13'h000a; 
        10'b0011101101: data <= 13'h1ff5; 
        10'b0011101110: data <= 13'h1fe7; 
        10'b0011101111: data <= 13'h1ff1; 
        10'b0011110000: data <= 13'h1ff7; 
        10'b0011110001: data <= 13'h0001; 
        10'b0011110010: data <= 13'h0003; 
        10'b0011110011: data <= 13'h0013; 
        10'b0011110100: data <= 13'h0014; 
        10'b0011110101: data <= 13'h001c; 
        10'b0011110110: data <= 13'h002c; 
        10'b0011110111: data <= 13'h003a; 
        10'b0011111000: data <= 13'h004d; 
        10'b0011111001: data <= 13'h0032; 
        10'b0011111010: data <= 13'h0009; 
        10'b0011111011: data <= 13'h1fff; 
        10'b0011111100: data <= 13'h1ffa; 
        10'b0011111101: data <= 13'h1ffc; 
        10'b0011111110: data <= 13'h1ff9; 
        10'b0011111111: data <= 13'h1ff1; 
        10'b0100000000: data <= 13'h1fef; 
        10'b0100000001: data <= 13'h1ff0; 
        10'b0100000010: data <= 13'h0002; 
        10'b0100000011: data <= 13'h1fff; 
        10'b0100000100: data <= 13'h000d; 
        10'b0100000101: data <= 13'h000c; 
        10'b0100000110: data <= 13'h000d; 
        10'b0100000111: data <= 13'h0022; 
        10'b0100001000: data <= 13'h0016; 
        10'b0100001001: data <= 13'h1ff7; 
        10'b0100001010: data <= 13'h1fe2; 
        10'b0100001011: data <= 13'h1fd5; 
        10'b0100001100: data <= 13'h1fd8; 
        10'b0100001101: data <= 13'h1fe9; 
        10'b0100001110: data <= 13'h1ffb; 
        10'b0100001111: data <= 13'h0000; 
        10'b0100010000: data <= 13'h0012; 
        10'b0100010001: data <= 13'h0027; 
        10'b0100010010: data <= 13'h0038; 
        10'b0100010011: data <= 13'h004d; 
        10'b0100010100: data <= 13'h0060; 
        10'b0100010101: data <= 13'h003f; 
        10'b0100010110: data <= 13'h000b; 
        10'b0100010111: data <= 13'h1ffc; 
        10'b0100011000: data <= 13'h1fff; 
        10'b0100011001: data <= 13'h1ffc; 
        10'b0100011010: data <= 13'h1ffa; 
        10'b0100011011: data <= 13'h1ffb; 
        10'b0100011100: data <= 13'h1ffb; 
        10'b0100011101: data <= 13'h1ffd; 
        10'b0100011110: data <= 13'h000b; 
        10'b0100011111: data <= 13'h0014; 
        10'b0100100000: data <= 13'h001f; 
        10'b0100100001: data <= 13'h0023; 
        10'b0100100010: data <= 13'h0021; 
        10'b0100100011: data <= 13'h0028; 
        10'b0100100100: data <= 13'h0022; 
        10'b0100100101: data <= 13'h001a; 
        10'b0100100110: data <= 13'h1ffa; 
        10'b0100100111: data <= 13'h1feb; 
        10'b0100101000: data <= 13'h1fdd; 
        10'b0100101001: data <= 13'h1fde; 
        10'b0100101010: data <= 13'h1fdd; 
        10'b0100101011: data <= 13'h1fd8; 
        10'b0100101100: data <= 13'h1fe5; 
        10'b0100101101: data <= 13'h1ff7; 
        10'b0100101110: data <= 13'h0005; 
        10'b0100101111: data <= 13'h001a; 
        10'b0100110000: data <= 13'h0033; 
        10'b0100110001: data <= 13'h0027; 
        10'b0100110010: data <= 13'h000d; 
        10'b0100110011: data <= 13'h1ffc; 
        10'b0100110100: data <= 13'h1ffa; 
        10'b0100110101: data <= 13'h0000; 
        10'b0100110110: data <= 13'h1ffb; 
        10'b0100110111: data <= 13'h1ffd; 
        10'b0100111000: data <= 13'h1ffb; 
        10'b0100111001: data <= 13'h1fff; 
        10'b0100111010: data <= 13'h0011; 
        10'b0100111011: data <= 13'h0015; 
        10'b0100111100: data <= 13'h001e; 
        10'b0100111101: data <= 13'h001c; 
        10'b0100111110: data <= 13'h0015; 
        10'b0100111111: data <= 13'h0017; 
        10'b0101000000: data <= 13'h0025; 
        10'b0101000001: data <= 13'h0023; 
        10'b0101000010: data <= 13'h0001; 
        10'b0101000011: data <= 13'h1fea; 
        10'b0101000100: data <= 13'h1fe5; 
        10'b0101000101: data <= 13'h1fe3; 
        10'b0101000110: data <= 13'h1fd9; 
        10'b0101000111: data <= 13'h1fca; 
        10'b0101001000: data <= 13'h1fb1; 
        10'b0101001001: data <= 13'h1fb8; 
        10'b0101001010: data <= 13'h1fc5; 
        10'b0101001011: data <= 13'h1fd5; 
        10'b0101001100: data <= 13'h1ff1; 
        10'b0101001101: data <= 13'h0002; 
        10'b0101001110: data <= 13'h0004; 
        10'b0101001111: data <= 13'h1ffd; 
        10'b0101010000: data <= 13'h1ffd; 
        10'b0101010001: data <= 13'h1ffe; 
        10'b0101010010: data <= 13'h1ffd; 
        10'b0101010011: data <= 13'h1ffb; 
        10'b0101010100: data <= 13'h1ffd; 
        10'b0101010101: data <= 13'h0009; 
        10'b0101010110: data <= 13'h0014; 
        10'b0101010111: data <= 13'h0012; 
        10'b0101011000: data <= 13'h000d; 
        10'b0101011001: data <= 13'h0007; 
        10'b0101011010: data <= 13'h0016; 
        10'b0101011011: data <= 13'h002d; 
        10'b0101011100: data <= 13'h002a; 
        10'b0101011101: data <= 13'h002b; 
        10'b0101011110: data <= 13'h0004; 
        10'b0101011111: data <= 13'h1fea; 
        10'b0101100000: data <= 13'h1fd7; 
        10'b0101100001: data <= 13'h1fdf; 
        10'b0101100010: data <= 13'h1fea; 
        10'b0101100011: data <= 13'h1fe0; 
        10'b0101100100: data <= 13'h1fdb; 
        10'b0101100101: data <= 13'h1fc3; 
        10'b0101100110: data <= 13'h1fba; 
        10'b0101100111: data <= 13'h1fc4; 
        10'b0101101000: data <= 13'h1fd8; 
        10'b0101101001: data <= 13'h1ff5; 
        10'b0101101010: data <= 13'h0001; 
        10'b0101101011: data <= 13'h0000; 
        10'b0101101100: data <= 13'h1ffe; 
        10'b0101101101: data <= 13'h1ffa; 
        10'b0101101110: data <= 13'h1ffa; 
        10'b0101101111: data <= 13'h1ffc; 
        10'b0101110000: data <= 13'h1fff; 
        10'b0101110001: data <= 13'h0005; 
        10'b0101110010: data <= 13'h000d; 
        10'b0101110011: data <= 13'h000a; 
        10'b0101110100: data <= 13'h000b; 
        10'b0101110101: data <= 13'h0009; 
        10'b0101110110: data <= 13'h001e; 
        10'b0101110111: data <= 13'h0022; 
        10'b0101111000: data <= 13'h0019; 
        10'b0101111001: data <= 13'h0018; 
        10'b0101111010: data <= 13'h1ffb; 
        10'b0101111011: data <= 13'h1fe6; 
        10'b0101111100: data <= 13'h1fd5; 
        10'b0101111101: data <= 13'h1fe9; 
        10'b0101111110: data <= 13'h1ff8; 
        10'b0101111111: data <= 13'h1ff7; 
        10'b0110000000: data <= 13'h1ffc; 
        10'b0110000001: data <= 13'h1fef; 
        10'b0110000010: data <= 13'h1fe1; 
        10'b0110000011: data <= 13'h1fd2; 
        10'b0110000100: data <= 13'h1fde; 
        10'b0110000101: data <= 13'h1ffa; 
        10'b0110000110: data <= 13'h1ffa; 
        10'b0110000111: data <= 13'h1fff; 
        10'b0110001000: data <= 13'h1ffe; 
        10'b0110001001: data <= 13'h1ffa; 
        10'b0110001010: data <= 13'h1ffd; 
        10'b0110001011: data <= 13'h1ff8; 
        10'b0110001100: data <= 13'h1ffd; 
        10'b0110001101: data <= 13'h1ffd; 
        10'b0110001110: data <= 13'h0000; 
        10'b0110001111: data <= 13'h1fff; 
        10'b0110010000: data <= 13'h000e; 
        10'b0110010001: data <= 13'h0016; 
        10'b0110010010: data <= 13'h001b; 
        10'b0110010011: data <= 13'h0005; 
        10'b0110010100: data <= 13'h0009; 
        10'b0110010101: data <= 13'h1ffe; 
        10'b0110010110: data <= 13'h1fed; 
        10'b0110010111: data <= 13'h1fea; 
        10'b0110011000: data <= 13'h1fe2; 
        10'b0110011001: data <= 13'h1fe5; 
        10'b0110011010: data <= 13'h1fe7; 
        10'b0110011011: data <= 13'h1ff4; 
        10'b0110011100: data <= 13'h1ff5; 
        10'b0110011101: data <= 13'h1ff6; 
        10'b0110011110: data <= 13'h1ffa; 
        10'b0110011111: data <= 13'h1fe7; 
        10'b0110100000: data <= 13'h1fef; 
        10'b0110100001: data <= 13'h1ff8; 
        10'b0110100010: data <= 13'h1ffd; 
        10'b0110100011: data <= 13'h1ff9; 
        10'b0110100100: data <= 13'h1ff9; 
        10'b0110100101: data <= 13'h0001; 
        10'b0110100110: data <= 13'h1ff9; 
        10'b0110100111: data <= 13'h1ffd; 
        10'b0110101000: data <= 13'h1ff5; 
        10'b0110101001: data <= 13'h1ff0; 
        10'b0110101010: data <= 13'h1fe9; 
        10'b0110101011: data <= 13'h1ff1; 
        10'b0110101100: data <= 13'h0005; 
        10'b0110101101: data <= 13'h0019; 
        10'b0110101110: data <= 13'h000c; 
        10'b0110101111: data <= 13'h000b; 
        10'b0110110000: data <= 13'h0009; 
        10'b0110110001: data <= 13'h1ff7; 
        10'b0110110010: data <= 13'h1fe4; 
        10'b0110110011: data <= 13'h1fe0; 
        10'b0110110100: data <= 13'h1fe3; 
        10'b0110110101: data <= 13'h1fe2; 
        10'b0110110110: data <= 13'h1feb; 
        10'b0110110111: data <= 13'h1fff; 
        10'b0110111000: data <= 13'h1ff9; 
        10'b0110111001: data <= 13'h1ffa; 
        10'b0110111010: data <= 13'h1ff9; 
        10'b0110111011: data <= 13'h1ff8; 
        10'b0110111100: data <= 13'h1ffa; 
        10'b0110111101: data <= 13'h0000; 
        10'b0110111110: data <= 13'h0001; 
        10'b0110111111: data <= 13'h1ffc; 
        10'b0111000000: data <= 13'h1ffc; 
        10'b0111000001: data <= 13'h1ffd; 
        10'b0111000010: data <= 13'h1ffe; 
        10'b0111000011: data <= 13'h1ff9; 
        10'b0111000100: data <= 13'h1ffc; 
        10'b0111000101: data <= 13'h1fee; 
        10'b0111000110: data <= 13'h1fdb; 
        10'b0111000111: data <= 13'h1fd5; 
        10'b0111001000: data <= 13'h1fe3; 
        10'b0111001001: data <= 13'h1ff0; 
        10'b0111001010: data <= 13'h1ffa; 
        10'b0111001011: data <= 13'h1ff7; 
        10'b0111001100: data <= 13'h1ffa; 
        10'b0111001101: data <= 13'h1fec; 
        10'b0111001110: data <= 13'h1fd9; 
        10'b0111001111: data <= 13'h1fe1; 
        10'b0111010000: data <= 13'h1fe9; 
        10'b0111010001: data <= 13'h1ff8; 
        10'b0111010010: data <= 13'h1ff8; 
        10'b0111010011: data <= 13'h0001; 
        10'b0111010100: data <= 13'h0006; 
        10'b0111010101: data <= 13'h0001; 
        10'b0111010110: data <= 13'h0007; 
        10'b0111010111: data <= 13'h0002; 
        10'b0111011000: data <= 13'h0001; 
        10'b0111011001: data <= 13'h0001; 
        10'b0111011010: data <= 13'h1ffc; 
        10'b0111011011: data <= 13'h1ffc; 
        10'b0111011100: data <= 13'h1ffb; 
        10'b0111011101: data <= 13'h0000; 
        10'b0111011110: data <= 13'h0000; 
        10'b0111011111: data <= 13'h0001; 
        10'b0111100000: data <= 13'h1ffb; 
        10'b0111100001: data <= 13'h0001; 
        10'b0111100010: data <= 13'h0003; 
        10'b0111100011: data <= 13'h1fe3; 
        10'b0111100100: data <= 13'h1fcc; 
        10'b0111100101: data <= 13'h1fcf; 
        10'b0111100110: data <= 13'h1fdd; 
        10'b0111100111: data <= 13'h1feb; 
        10'b0111101000: data <= 13'h1fdf; 
        10'b0111101001: data <= 13'h1fd6; 
        10'b0111101010: data <= 13'h1fd7; 
        10'b0111101011: data <= 13'h1fed; 
        10'b0111101100: data <= 13'h1ff8; 
        10'b0111101101: data <= 13'h000c; 
        10'b0111101110: data <= 13'h0013; 
        10'b0111101111: data <= 13'h000c; 
        10'b0111110000: data <= 13'h000c; 
        10'b0111110001: data <= 13'h0004; 
        10'b0111110010: data <= 13'h0000; 
        10'b0111110011: data <= 13'h0007; 
        10'b0111110100: data <= 13'h0007; 
        10'b0111110101: data <= 13'h1ffa; 
        10'b0111110110: data <= 13'h0000; 
        10'b0111110111: data <= 13'h0000; 
        10'b0111111000: data <= 13'h0001; 
        10'b0111111001: data <= 13'h1ffb; 
        10'b0111111010: data <= 13'h1ffd; 
        10'b0111111011: data <= 13'h1ffc; 
        10'b0111111100: data <= 13'h000a; 
        10'b0111111101: data <= 13'h000e; 
        10'b0111111110: data <= 13'h0020; 
        10'b0111111111: data <= 13'h0006; 
        10'b1000000000: data <= 13'h1fe1; 
        10'b1000000001: data <= 13'h1fd3; 
        10'b1000000010: data <= 13'h1fc5; 
        10'b1000000011: data <= 13'h1fcb; 
        10'b1000000100: data <= 13'h1fda; 
        10'b1000000101: data <= 13'h1fea; 
        10'b1000000110: data <= 13'h1ff5; 
        10'b1000000111: data <= 13'h1ffb; 
        10'b1000001000: data <= 13'h1fff; 
        10'b1000001001: data <= 13'h000f; 
        10'b1000001010: data <= 13'h0007; 
        10'b1000001011: data <= 13'h000d; 
        10'b1000001100: data <= 13'h0009; 
        10'b1000001101: data <= 13'h000d; 
        10'b1000001110: data <= 13'h000a; 
        10'b1000001111: data <= 13'h000e; 
        10'b1000010000: data <= 13'h0007; 
        10'b1000010001: data <= 13'h0001; 
        10'b1000010010: data <= 13'h1ffb; 
        10'b1000010011: data <= 13'h1ffe; 
        10'b1000010100: data <= 13'h0000; 
        10'b1000010101: data <= 13'h1ffb; 
        10'b1000010110: data <= 13'h1ffd; 
        10'b1000010111: data <= 13'h0001; 
        10'b1000011000: data <= 13'h0010; 
        10'b1000011001: data <= 13'h001b; 
        10'b1000011010: data <= 13'h0024; 
        10'b1000011011: data <= 13'h0018; 
        10'b1000011100: data <= 13'h000f; 
        10'b1000011101: data <= 13'h0005; 
        10'b1000011110: data <= 13'h1ff5; 
        10'b1000011111: data <= 13'h1ff4; 
        10'b1000100000: data <= 13'h0001; 
        10'b1000100001: data <= 13'h000f; 
        10'b1000100010: data <= 13'h0005; 
        10'b1000100011: data <= 13'h0008; 
        10'b1000100100: data <= 13'h0008; 
        10'b1000100101: data <= 13'h1ffe; 
        10'b1000100110: data <= 13'h0006; 
        10'b1000100111: data <= 13'h0006; 
        10'b1000101000: data <= 13'h0001; 
        10'b1000101001: data <= 13'h0009; 
        10'b1000101010: data <= 13'h0010; 
        10'b1000101011: data <= 13'h000c; 
        10'b1000101100: data <= 13'h0001; 
        10'b1000101101: data <= 13'h0000; 
        10'b1000101110: data <= 13'h0000; 
        10'b1000101111: data <= 13'h1ffa; 
        10'b1000110000: data <= 13'h0000; 
        10'b1000110001: data <= 13'h1ff9; 
        10'b1000110010: data <= 13'h1ffc; 
        10'b1000110011: data <= 13'h1ffa; 
        10'b1000110100: data <= 13'h0002; 
        10'b1000110101: data <= 13'h0011; 
        10'b1000110110: data <= 13'h0014; 
        10'b1000110111: data <= 13'h0019; 
        10'b1000111000: data <= 13'h0023; 
        10'b1000111001: data <= 13'h001d; 
        10'b1000111010: data <= 13'h001a; 
        10'b1000111011: data <= 13'h0026; 
        10'b1000111100: data <= 13'h0017; 
        10'b1000111101: data <= 13'h0012; 
        10'b1000111110: data <= 13'h1ffb; 
        10'b1000111111: data <= 13'h1ffb; 
        10'b1001000000: data <= 13'h000d; 
        10'b1001000001: data <= 13'h0007; 
        10'b1001000010: data <= 13'h000b; 
        10'b1001000011: data <= 13'h000e; 
        10'b1001000100: data <= 13'h000c; 
        10'b1001000101: data <= 13'h000a; 
        10'b1001000110: data <= 13'h0017; 
        10'b1001000111: data <= 13'h0012; 
        10'b1001001000: data <= 13'h1ffe; 
        10'b1001001001: data <= 13'h1ff9; 
        10'b1001001010: data <= 13'h1ffd; 
        10'b1001001011: data <= 13'h1ffb; 
        10'b1001001100: data <= 13'h1ffb; 
        10'b1001001101: data <= 13'h0000; 
        10'b1001001110: data <= 13'h1ff8; 
        10'b1001001111: data <= 13'h1ffd; 
        10'b1001010000: data <= 13'h0007; 
        10'b1001010001: data <= 13'h1ffe; 
        10'b1001010010: data <= 13'h0008; 
        10'b1001010011: data <= 13'h0017; 
        10'b1001010100: data <= 13'h0021; 
        10'b1001010101: data <= 13'h0015; 
        10'b1001010110: data <= 13'h0012; 
        10'b1001010111: data <= 13'h000a; 
        10'b1001011000: data <= 13'h000d; 
        10'b1001011001: data <= 13'h0008; 
        10'b1001011010: data <= 13'h0008; 
        10'b1001011011: data <= 13'h000a; 
        10'b1001011100: data <= 13'h0003; 
        10'b1001011101: data <= 13'h0008; 
        10'b1001011110: data <= 13'h0004; 
        10'b1001011111: data <= 13'h000d; 
        10'b1001100000: data <= 13'h000d; 
        10'b1001100001: data <= 13'h0015; 
        10'b1001100010: data <= 13'h001a; 
        10'b1001100011: data <= 13'h0006; 
        10'b1001100100: data <= 13'h0000; 
        10'b1001100101: data <= 13'h1ffa; 
        10'b1001100110: data <= 13'h1ffb; 
        10'b1001100111: data <= 13'h1ffb; 
        10'b1001101000: data <= 13'h1ffe; 
        10'b1001101001: data <= 13'h1ff9; 
        10'b1001101010: data <= 13'h1ffc; 
        10'b1001101011: data <= 13'h1ffb; 
        10'b1001101100: data <= 13'h0002; 
        10'b1001101101: data <= 13'h1ffd; 
        10'b1001101110: data <= 13'h1ff8; 
        10'b1001101111: data <= 13'h1fff; 
        10'b1001110000: data <= 13'h000d; 
        10'b1001110001: data <= 13'h0013; 
        10'b1001110010: data <= 13'h0003; 
        10'b1001110011: data <= 13'h0010; 
        10'b1001110100: data <= 13'h001b; 
        10'b1001110101: data <= 13'h0021; 
        10'b1001110110: data <= 13'h0011; 
        10'b1001110111: data <= 13'h0003; 
        10'b1001111000: data <= 13'h0002; 
        10'b1001111001: data <= 13'h0004; 
        10'b1001111010: data <= 13'h0009; 
        10'b1001111011: data <= 13'h0009; 
        10'b1001111100: data <= 13'h000f; 
        10'b1001111101: data <= 13'h000d; 
        10'b1001111110: data <= 13'h000e; 
        10'b1001111111: data <= 13'h0005; 
        10'b1010000000: data <= 13'h1fff; 
        10'b1010000001: data <= 13'h0001; 
        10'b1010000010: data <= 13'h1ffd; 
        10'b1010000011: data <= 13'h1ffe; 
        10'b1010000100: data <= 13'h1ffa; 
        10'b1010000101: data <= 13'h1ffd; 
        10'b1010000110: data <= 13'h1ffe; 
        10'b1010000111: data <= 13'h1ffe; 
        10'b1010001000: data <= 13'h1ffa; 
        10'b1010001001: data <= 13'h1ffc; 
        10'b1010001010: data <= 13'h1ff5; 
        10'b1010001011: data <= 13'h1ffb; 
        10'b1010001100: data <= 13'h000a; 
        10'b1010001101: data <= 13'h000a; 
        10'b1010001110: data <= 13'h000a; 
        10'b1010001111: data <= 13'h0012; 
        10'b1010010000: data <= 13'h0011; 
        10'b1010010001: data <= 13'h000c; 
        10'b1010010010: data <= 13'h000d; 
        10'b1010010011: data <= 13'h000c; 
        10'b1010010100: data <= 13'h000c; 
        10'b1010010101: data <= 13'h0005; 
        10'b1010010110: data <= 13'h1ffa; 
        10'b1010010111: data <= 13'h1fff; 
        10'b1010011000: data <= 13'h0006; 
        10'b1010011001: data <= 13'h0002; 
        10'b1010011010: data <= 13'h0008; 
        10'b1010011011: data <= 13'h1ffb; 
        10'b1010011100: data <= 13'h0001; 
        10'b1010011101: data <= 13'h1ffc; 
        10'b1010011110: data <= 13'h1ffc; 
        10'b1010011111: data <= 13'h0001; 
        10'b1010100000: data <= 13'h1fff; 
        10'b1010100001: data <= 13'h1ffc; 
        10'b1010100010: data <= 13'h1ffc; 
        10'b1010100011: data <= 13'h0001; 
        10'b1010100100: data <= 13'h1ff8; 
        10'b1010100101: data <= 13'h1ff8; 
        10'b1010100110: data <= 13'h1ffd; 
        10'b1010100111: data <= 13'h1fff; 
        10'b1010101000: data <= 13'h0000; 
        10'b1010101001: data <= 13'h000d; 
        10'b1010101010: data <= 13'h0011; 
        10'b1010101011: data <= 13'h000d; 
        10'b1010101100: data <= 13'h0008; 
        10'b1010101101: data <= 13'h000c; 
        10'b1010101110: data <= 13'h0016; 
        10'b1010101111: data <= 13'h0012; 
        10'b1010110000: data <= 13'h000b; 
        10'b1010110001: data <= 13'h0005; 
        10'b1010110010: data <= 13'h000a; 
        10'b1010110011: data <= 13'h0006; 
        10'b1010110100: data <= 13'h0000; 
        10'b1010110101: data <= 13'h1fff; 
        10'b1010110110: data <= 13'h1ffe; 
        10'b1010110111: data <= 13'h0000; 
        10'b1010111000: data <= 13'h1ffb; 
        10'b1010111001: data <= 13'h1ffe; 
        10'b1010111010: data <= 13'h0001; 
        10'b1010111011: data <= 13'h1ffa; 
        10'b1010111100: data <= 13'h1ffd; 
        10'b1010111101: data <= 13'h0000; 
        10'b1010111110: data <= 13'h0001; 
        10'b1010111111: data <= 13'h1ff9; 
        10'b1011000000: data <= 13'h0000; 
        10'b1011000001: data <= 13'h1ffe; 
        10'b1011000010: data <= 13'h1ff8; 
        10'b1011000011: data <= 13'h1ffd; 
        10'b1011000100: data <= 13'h1ff9; 
        10'b1011000101: data <= 13'h0004; 
        10'b1011000110: data <= 13'h0003; 
        10'b1011000111: data <= 13'h0009; 
        10'b1011001000: data <= 13'h0009; 
        10'b1011001001: data <= 13'h000f; 
        10'b1011001010: data <= 13'h0001; 
        10'b1011001011: data <= 13'h0005; 
        10'b1011001100: data <= 13'h0004; 
        10'b1011001101: data <= 13'h0008; 
        10'b1011001110: data <= 13'h1ffb; 
        10'b1011001111: data <= 13'h0000; 
        10'b1011010000: data <= 13'h1ff8; 
        10'b1011010001: data <= 13'h0001; 
        10'b1011010010: data <= 13'h1ffd; 
        10'b1011010011: data <= 13'h1ffa; 
        10'b1011010100: data <= 13'h1fff; 
        10'b1011010101: data <= 13'h0000; 
        10'b1011010110: data <= 13'h1ff9; 
        10'b1011010111: data <= 13'h1ffc; 
        10'b1011011000: data <= 13'h1ffe; 
        10'b1011011001: data <= 13'h1ffe; 
        10'b1011011010: data <= 13'h1ffb; 
        10'b1011011011: data <= 13'h1ffc; 
        10'b1011011100: data <= 13'h1ffc; 
        10'b1011011101: data <= 13'h1ffc; 
        10'b1011011110: data <= 13'h1fff; 
        10'b1011011111: data <= 13'h1ffb; 
        10'b1011100000: data <= 13'h1ff9; 
        10'b1011100001: data <= 13'h1ffc; 
        10'b1011100010: data <= 13'h1ffb; 
        10'b1011100011: data <= 13'h1fff; 
        10'b1011100100: data <= 13'h0000; 
        10'b1011100101: data <= 13'h1ffe; 
        10'b1011100110: data <= 13'h1ffb; 
        10'b1011100111: data <= 13'h1ffd; 
        10'b1011101000: data <= 13'h1fff; 
        10'b1011101001: data <= 13'h1ffb; 
        10'b1011101010: data <= 13'h1ff6; 
        10'b1011101011: data <= 13'h1ff8; 
        10'b1011101100: data <= 13'h1ffe; 
        10'b1011101101: data <= 13'h1ffe; 
        10'b1011101110: data <= 13'h1ffb; 
        10'b1011101111: data <= 13'h1fff; 
        10'b1011110000: data <= 13'h1ffd; 
        10'b1011110001: data <= 13'h1ffe; 
        10'b1011110010: data <= 13'h1ffc; 
        10'b1011110011: data <= 13'h1ff9; 
        10'b1011110100: data <= 13'h1ffe; 
        10'b1011110101: data <= 13'h1fff; 
        10'b1011110110: data <= 13'h1fff; 
        10'b1011110111: data <= 13'h1ffe; 
        10'b1011111000: data <= 13'h1ffa; 
        10'b1011111001: data <= 13'h0000; 
        10'b1011111010: data <= 13'h1ffc; 
        10'b1011111011: data <= 13'h1ffb; 
        10'b1011111100: data <= 13'h0001; 
        10'b1011111101: data <= 13'h1ffc; 
        10'b1011111110: data <= 13'h1ffb; 
        10'b1011111111: data <= 13'h1fff; 
        10'b1100000000: data <= 13'h1ffd; 
        10'b1100000001: data <= 13'h1ff9; 
        10'b1100000010: data <= 13'h0000; 
        10'b1100000011: data <= 13'h1ffe; 
        10'b1100000100: data <= 13'h1ff9; 
        10'b1100000101: data <= 13'h1ff8; 
        10'b1100000110: data <= 13'h1ffa; 
        10'b1100000111: data <= 13'h1ff8; 
        10'b1100001000: data <= 13'h0000; 
        10'b1100001001: data <= 13'h1ffc; 
        10'b1100001010: data <= 13'h0001; 
        10'b1100001011: data <= 13'h1ff9; 
        10'b1100001100: data <= 13'h1ffe; 
        10'b1100001101: data <= 13'h1ffd; 
        10'b1100001110: data <= 13'h1ffa; 
        10'b1100001111: data <= 13'h1fff; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 8) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 14'h3ff7; 
        10'b0000000001: data <= 14'h3fff; 
        10'b0000000010: data <= 14'h3fff; 
        10'b0000000011: data <= 14'h3ff4; 
        10'b0000000100: data <= 14'h3ffa; 
        10'b0000000101: data <= 14'h3ff9; 
        10'b0000000110: data <= 14'h0000; 
        10'b0000000111: data <= 14'h3ff8; 
        10'b0000001000: data <= 14'h3ffd; 
        10'b0000001001: data <= 14'h0003; 
        10'b0000001010: data <= 14'h3ffd; 
        10'b0000001011: data <= 14'h3ffd; 
        10'b0000001100: data <= 14'h3ff7; 
        10'b0000001101: data <= 14'h3fff; 
        10'b0000001110: data <= 14'h3ff4; 
        10'b0000001111: data <= 14'h3ff6; 
        10'b0000010000: data <= 14'h3ff2; 
        10'b0000010001: data <= 14'h3ff5; 
        10'b0000010010: data <= 14'h3ffe; 
        10'b0000010011: data <= 14'h3ffd; 
        10'b0000010100: data <= 14'h3ff2; 
        10'b0000010101: data <= 14'h3ffb; 
        10'b0000010110: data <= 14'h3ffc; 
        10'b0000010111: data <= 14'h3ff9; 
        10'b0000011000: data <= 14'h3ff3; 
        10'b0000011001: data <= 14'h3ffb; 
        10'b0000011010: data <= 14'h3ffc; 
        10'b0000011011: data <= 14'h3ff8; 
        10'b0000011100: data <= 14'h3fff; 
        10'b0000011101: data <= 14'h3ff1; 
        10'b0000011110: data <= 14'h0000; 
        10'b0000011111: data <= 14'h3ff3; 
        10'b0000100000: data <= 14'h3fff; 
        10'b0000100001: data <= 14'h3ff8; 
        10'b0000100010: data <= 14'h3ffc; 
        10'b0000100011: data <= 14'h3ff8; 
        10'b0000100100: data <= 14'h3ff6; 
        10'b0000100101: data <= 14'h3ffc; 
        10'b0000100110: data <= 14'h0001; 
        10'b0000100111: data <= 14'h3ff4; 
        10'b0000101000: data <= 14'h3ff8; 
        10'b0000101001: data <= 14'h3ff5; 
        10'b0000101010: data <= 14'h3ff2; 
        10'b0000101011: data <= 14'h3ffe; 
        10'b0000101100: data <= 14'h3ff7; 
        10'b0000101101: data <= 14'h3ff5; 
        10'b0000101110: data <= 14'h3ff7; 
        10'b0000101111: data <= 14'h3ff6; 
        10'b0000110000: data <= 14'h3ffd; 
        10'b0000110001: data <= 14'h3ff3; 
        10'b0000110010: data <= 14'h0000; 
        10'b0000110011: data <= 14'h3ff4; 
        10'b0000110100: data <= 14'h0000; 
        10'b0000110101: data <= 14'h3fff; 
        10'b0000110110: data <= 14'h3ff5; 
        10'b0000110111: data <= 14'h3ffa; 
        10'b0000111000: data <= 14'h3ffa; 
        10'b0000111001: data <= 14'h3ffd; 
        10'b0000111010: data <= 14'h3ff8; 
        10'b0000111011: data <= 14'h3ff2; 
        10'b0000111100: data <= 14'h3ff5; 
        10'b0000111101: data <= 14'h3ffb; 
        10'b0000111110: data <= 14'h0000; 
        10'b0000111111: data <= 14'h3ffc; 
        10'b0001000000: data <= 14'h3ff6; 
        10'b0001000001: data <= 14'h3ff8; 
        10'b0001000010: data <= 14'h0002; 
        10'b0001000011: data <= 14'h3ff1; 
        10'b0001000100: data <= 14'h3fff; 
        10'b0001000101: data <= 14'h3ff6; 
        10'b0001000110: data <= 14'h3ff2; 
        10'b0001000111: data <= 14'h3ff5; 
        10'b0001001000: data <= 14'h3ff7; 
        10'b0001001001: data <= 14'h3ffb; 
        10'b0001001010: data <= 14'h3ff8; 
        10'b0001001011: data <= 14'h3ff8; 
        10'b0001001100: data <= 14'h0003; 
        10'b0001001101: data <= 14'h0000; 
        10'b0001001110: data <= 14'h0001; 
        10'b0001001111: data <= 14'h3ff5; 
        10'b0001010000: data <= 14'h3ff2; 
        10'b0001010001: data <= 14'h3ff9; 
        10'b0001010010: data <= 14'h3fff; 
        10'b0001010011: data <= 14'h3ffc; 
        10'b0001010100: data <= 14'h3ffd; 
        10'b0001010101: data <= 14'h3ffc; 
        10'b0001010110: data <= 14'h3ff5; 
        10'b0001010111: data <= 14'h3fff; 
        10'b0001011000: data <= 14'h3ff4; 
        10'b0001011001: data <= 14'h3ff8; 
        10'b0001011010: data <= 14'h3ff1; 
        10'b0001011011: data <= 14'h3ff6; 
        10'b0001011100: data <= 14'h3ff2; 
        10'b0001011101: data <= 14'h3ff6; 
        10'b0001011110: data <= 14'h3fe8; 
        10'b0001011111: data <= 14'h3fe1; 
        10'b0001100000: data <= 14'h3fef; 
        10'b0001100001: data <= 14'h3ff0; 
        10'b0001100010: data <= 14'h3fec; 
        10'b0001100011: data <= 14'h3ff9; 
        10'b0001100100: data <= 14'h3ffd; 
        10'b0001100101: data <= 14'h3ff0; 
        10'b0001100110: data <= 14'h3ff7; 
        10'b0001100111: data <= 14'h3ffd; 
        10'b0001101000: data <= 14'h3ffe; 
        10'b0001101001: data <= 14'h3ff9; 
        10'b0001101010: data <= 14'h3ff0; 
        10'b0001101011: data <= 14'h3ff5; 
        10'b0001101100: data <= 14'h3fed; 
        10'b0001101101: data <= 14'h0002; 
        10'b0001101110: data <= 14'h0001; 
        10'b0001101111: data <= 14'h3ff3; 
        10'b0001110000: data <= 14'h3ff3; 
        10'b0001110001: data <= 14'h3ff8; 
        10'b0001110010: data <= 14'h0001; 
        10'b0001110011: data <= 14'h0001; 
        10'b0001110100: data <= 14'h0002; 
        10'b0001110101: data <= 14'h3ff6; 
        10'b0001110110: data <= 14'h3ff6; 
        10'b0001110111: data <= 14'h3fea; 
        10'b0001111000: data <= 14'h3fdc; 
        10'b0001111001: data <= 14'h3fd0; 
        10'b0001111010: data <= 14'h3fb9; 
        10'b0001111011: data <= 14'h3fd3; 
        10'b0001111100: data <= 14'h3fd2; 
        10'b0001111101: data <= 14'h3fc3; 
        10'b0001111110: data <= 14'h3fde; 
        10'b0001111111: data <= 14'h0000; 
        10'b0010000000: data <= 14'h3ffc; 
        10'b0010000001: data <= 14'h000b; 
        10'b0010000010: data <= 14'h3ffd; 
        10'b0010000011: data <= 14'h3fef; 
        10'b0010000100: data <= 14'h3fe9; 
        10'b0010000101: data <= 14'h3ff4; 
        10'b0010000110: data <= 14'h3ff6; 
        10'b0010000111: data <= 14'h3ff9; 
        10'b0010001000: data <= 14'h3ff7; 
        10'b0010001001: data <= 14'h0003; 
        10'b0010001010: data <= 14'h0002; 
        10'b0010001011: data <= 14'h3ffa; 
        10'b0010001100: data <= 14'h3ffb; 
        10'b0010001101: data <= 14'h0003; 
        10'b0010001110: data <= 14'h3ff5; 
        10'b0010001111: data <= 14'h3ff3; 
        10'b0010010000: data <= 14'h3ff7; 
        10'b0010010001: data <= 14'h3fea; 
        10'b0010010010: data <= 14'h3fdf; 
        10'b0010010011: data <= 14'h3fe0; 
        10'b0010010100: data <= 14'h3feb; 
        10'b0010010101: data <= 14'h3ffc; 
        10'b0010010110: data <= 14'h0007; 
        10'b0010010111: data <= 14'h0008; 
        10'b0010011000: data <= 14'h3ff5; 
        10'b0010011001: data <= 14'h3ff0; 
        10'b0010011010: data <= 14'h3ff6; 
        10'b0010011011: data <= 14'h3ffb; 
        10'b0010011100: data <= 14'h0010; 
        10'b0010011101: data <= 14'h0011; 
        10'b0010011110: data <= 14'h0020; 
        10'b0010011111: data <= 14'h0014; 
        10'b0010100000: data <= 14'h0013; 
        10'b0010100001: data <= 14'h0019; 
        10'b0010100010: data <= 14'h002d; 
        10'b0010100011: data <= 14'h0027; 
        10'b0010100100: data <= 14'h001b; 
        10'b0010100101: data <= 14'h000f; 
        10'b0010100110: data <= 14'h0009; 
        10'b0010100111: data <= 14'h0003; 
        10'b0010101000: data <= 14'h3ff4; 
        10'b0010101001: data <= 14'h3ff3; 
        10'b0010101010: data <= 14'h0002; 
        10'b0010101011: data <= 14'h3ff3; 
        10'b0010101100: data <= 14'h3ff0; 
        10'b0010101101: data <= 14'h3fd9; 
        10'b0010101110: data <= 14'h3fef; 
        10'b0010101111: data <= 14'h3ffe; 
        10'b0010110000: data <= 14'h3fff; 
        10'b0010110001: data <= 14'h0010; 
        10'b0010110010: data <= 14'h0021; 
        10'b0010110011: data <= 14'h001b; 
        10'b0010110100: data <= 14'h0005; 
        10'b0010110101: data <= 14'h000a; 
        10'b0010110110: data <= 14'h3ffb; 
        10'b0010110111: data <= 14'h3ff0; 
        10'b0010111000: data <= 14'h3ff7; 
        10'b0010111001: data <= 14'h3ff8; 
        10'b0010111010: data <= 14'h0000; 
        10'b0010111011: data <= 14'h001f; 
        10'b0010111100: data <= 14'h0012; 
        10'b0010111101: data <= 14'h0014; 
        10'b0010111110: data <= 14'h003e; 
        10'b0010111111: data <= 14'h004a; 
        10'b0011000000: data <= 14'h0054; 
        10'b0011000001: data <= 14'h002c; 
        10'b0011000010: data <= 14'h0016; 
        10'b0011000011: data <= 14'h0005; 
        10'b0011000100: data <= 14'h3ff9; 
        10'b0011000101: data <= 14'h3ffc; 
        10'b0011000110: data <= 14'h3ffb; 
        10'b0011000111: data <= 14'h3ff0; 
        10'b0011001000: data <= 14'h3fd3; 
        10'b0011001001: data <= 14'h3fcb; 
        10'b0011001010: data <= 14'h3fe0; 
        10'b0011001011: data <= 14'h0004; 
        10'b0011001100: data <= 14'h0015; 
        10'b0011001101: data <= 14'h002a; 
        10'b0011001110: data <= 14'h0028; 
        10'b0011001111: data <= 14'h0023; 
        10'b0011010000: data <= 14'h000a; 
        10'b0011010001: data <= 14'h3ffd; 
        10'b0011010010: data <= 14'h3ff5; 
        10'b0011010011: data <= 14'h0001; 
        10'b0011010100: data <= 14'h0011; 
        10'b0011010101: data <= 14'h0010; 
        10'b0011010110: data <= 14'h0014; 
        10'b0011010111: data <= 14'h002d; 
        10'b0011011000: data <= 14'h0027; 
        10'b0011011001: data <= 14'h002e; 
        10'b0011011010: data <= 14'h0041; 
        10'b0011011011: data <= 14'h0057; 
        10'b0011011100: data <= 14'h006a; 
        10'b0011011101: data <= 14'h004d; 
        10'b0011011110: data <= 14'h000c; 
        10'b0011011111: data <= 14'h3ffe; 
        10'b0011100000: data <= 14'h3ffd; 
        10'b0011100001: data <= 14'h0003; 
        10'b0011100010: data <= 14'h0000; 
        10'b0011100011: data <= 14'h3fea; 
        10'b0011100100: data <= 14'h3fbf; 
        10'b0011100101: data <= 14'h3fc8; 
        10'b0011100110: data <= 14'h3fd8; 
        10'b0011100111: data <= 14'h0002; 
        10'b0011101000: data <= 14'h001f; 
        10'b0011101001: data <= 14'h0009; 
        10'b0011101010: data <= 14'h0011; 
        10'b0011101011: data <= 14'h0021; 
        10'b0011101100: data <= 14'h0014; 
        10'b0011101101: data <= 14'h3fe9; 
        10'b0011101110: data <= 14'h3fcf; 
        10'b0011101111: data <= 14'h3fe2; 
        10'b0011110000: data <= 14'h3fee; 
        10'b0011110001: data <= 14'h0002; 
        10'b0011110010: data <= 14'h0005; 
        10'b0011110011: data <= 14'h0025; 
        10'b0011110100: data <= 14'h0027; 
        10'b0011110101: data <= 14'h0038; 
        10'b0011110110: data <= 14'h0059; 
        10'b0011110111: data <= 14'h0074; 
        10'b0011111000: data <= 14'h009b; 
        10'b0011111001: data <= 14'h0064; 
        10'b0011111010: data <= 14'h0012; 
        10'b0011111011: data <= 14'h3ffe; 
        10'b0011111100: data <= 14'h3ff3; 
        10'b0011111101: data <= 14'h3ff8; 
        10'b0011111110: data <= 14'h3ff2; 
        10'b0011111111: data <= 14'h3fe2; 
        10'b0100000000: data <= 14'h3fdd; 
        10'b0100000001: data <= 14'h3fe0; 
        10'b0100000010: data <= 14'h0004; 
        10'b0100000011: data <= 14'h3ffe; 
        10'b0100000100: data <= 14'h001b; 
        10'b0100000101: data <= 14'h0017; 
        10'b0100000110: data <= 14'h0019; 
        10'b0100000111: data <= 14'h0044; 
        10'b0100001000: data <= 14'h002c; 
        10'b0100001001: data <= 14'h3fee; 
        10'b0100001010: data <= 14'h3fc4; 
        10'b0100001011: data <= 14'h3fab; 
        10'b0100001100: data <= 14'h3fb0; 
        10'b0100001101: data <= 14'h3fd2; 
        10'b0100001110: data <= 14'h3ff5; 
        10'b0100001111: data <= 14'h0000; 
        10'b0100010000: data <= 14'h0024; 
        10'b0100010001: data <= 14'h004e; 
        10'b0100010010: data <= 14'h0070; 
        10'b0100010011: data <= 14'h009a; 
        10'b0100010100: data <= 14'h00c1; 
        10'b0100010101: data <= 14'h007f; 
        10'b0100010110: data <= 14'h0017; 
        10'b0100010111: data <= 14'h3ff7; 
        10'b0100011000: data <= 14'h3ffd; 
        10'b0100011001: data <= 14'h3ff7; 
        10'b0100011010: data <= 14'h3ff4; 
        10'b0100011011: data <= 14'h3ff6; 
        10'b0100011100: data <= 14'h3ff6; 
        10'b0100011101: data <= 14'h3ff9; 
        10'b0100011110: data <= 14'h0016; 
        10'b0100011111: data <= 14'h0028; 
        10'b0100100000: data <= 14'h003f; 
        10'b0100100001: data <= 14'h0046; 
        10'b0100100010: data <= 14'h0043; 
        10'b0100100011: data <= 14'h0051; 
        10'b0100100100: data <= 14'h0043; 
        10'b0100100101: data <= 14'h0034; 
        10'b0100100110: data <= 14'h3ff5; 
        10'b0100100111: data <= 14'h3fd6; 
        10'b0100101000: data <= 14'h3fba; 
        10'b0100101001: data <= 14'h3fbc; 
        10'b0100101010: data <= 14'h3fba; 
        10'b0100101011: data <= 14'h3fb0; 
        10'b0100101100: data <= 14'h3fc9; 
        10'b0100101101: data <= 14'h3fef; 
        10'b0100101110: data <= 14'h0009; 
        10'b0100101111: data <= 14'h0034; 
        10'b0100110000: data <= 14'h0067; 
        10'b0100110001: data <= 14'h004d; 
        10'b0100110010: data <= 14'h001a; 
        10'b0100110011: data <= 14'h3ff7; 
        10'b0100110100: data <= 14'h3ff4; 
        10'b0100110101: data <= 14'h0000; 
        10'b0100110110: data <= 14'h3ff6; 
        10'b0100110111: data <= 14'h3ffa; 
        10'b0100111000: data <= 14'h3ff6; 
        10'b0100111001: data <= 14'h3fff; 
        10'b0100111010: data <= 14'h0022; 
        10'b0100111011: data <= 14'h002a; 
        10'b0100111100: data <= 14'h003d; 
        10'b0100111101: data <= 14'h0038; 
        10'b0100111110: data <= 14'h0029; 
        10'b0100111111: data <= 14'h002d; 
        10'b0101000000: data <= 14'h004b; 
        10'b0101000001: data <= 14'h0046; 
        10'b0101000010: data <= 14'h0001; 
        10'b0101000011: data <= 14'h3fd4; 
        10'b0101000100: data <= 14'h3fca; 
        10'b0101000101: data <= 14'h3fc6; 
        10'b0101000110: data <= 14'h3fb2; 
        10'b0101000111: data <= 14'h3f94; 
        10'b0101001000: data <= 14'h3f63; 
        10'b0101001001: data <= 14'h3f70; 
        10'b0101001010: data <= 14'h3f8a; 
        10'b0101001011: data <= 14'h3faa; 
        10'b0101001100: data <= 14'h3fe1; 
        10'b0101001101: data <= 14'h0003; 
        10'b0101001110: data <= 14'h0009; 
        10'b0101001111: data <= 14'h3ffb; 
        10'b0101010000: data <= 14'h3ffb; 
        10'b0101010001: data <= 14'h3ffc; 
        10'b0101010010: data <= 14'h3ffa; 
        10'b0101010011: data <= 14'h3ff7; 
        10'b0101010100: data <= 14'h3ff9; 
        10'b0101010101: data <= 14'h0011; 
        10'b0101010110: data <= 14'h0027; 
        10'b0101010111: data <= 14'h0023; 
        10'b0101011000: data <= 14'h001a; 
        10'b0101011001: data <= 14'h000f; 
        10'b0101011010: data <= 14'h002c; 
        10'b0101011011: data <= 14'h005b; 
        10'b0101011100: data <= 14'h0055; 
        10'b0101011101: data <= 14'h0057; 
        10'b0101011110: data <= 14'h0009; 
        10'b0101011111: data <= 14'h3fd4; 
        10'b0101100000: data <= 14'h3fae; 
        10'b0101100001: data <= 14'h3fbe; 
        10'b0101100010: data <= 14'h3fd3; 
        10'b0101100011: data <= 14'h3fc0; 
        10'b0101100100: data <= 14'h3fb7; 
        10'b0101100101: data <= 14'h3f86; 
        10'b0101100110: data <= 14'h3f75; 
        10'b0101100111: data <= 14'h3f87; 
        10'b0101101000: data <= 14'h3faf; 
        10'b0101101001: data <= 14'h3fe9; 
        10'b0101101010: data <= 14'h0001; 
        10'b0101101011: data <= 14'h0000; 
        10'b0101101100: data <= 14'h3ffb; 
        10'b0101101101: data <= 14'h3ff5; 
        10'b0101101110: data <= 14'h3ff4; 
        10'b0101101111: data <= 14'h3ff8; 
        10'b0101110000: data <= 14'h3ffd; 
        10'b0101110001: data <= 14'h0009; 
        10'b0101110010: data <= 14'h001a; 
        10'b0101110011: data <= 14'h0013; 
        10'b0101110100: data <= 14'h0016; 
        10'b0101110101: data <= 14'h0013; 
        10'b0101110110: data <= 14'h003d; 
        10'b0101110111: data <= 14'h0044; 
        10'b0101111000: data <= 14'h0033; 
        10'b0101111001: data <= 14'h002f; 
        10'b0101111010: data <= 14'h3ff7; 
        10'b0101111011: data <= 14'h3fcc; 
        10'b0101111100: data <= 14'h3fab; 
        10'b0101111101: data <= 14'h3fd3; 
        10'b0101111110: data <= 14'h3ff0; 
        10'b0101111111: data <= 14'h3fee; 
        10'b0110000000: data <= 14'h3ff7; 
        10'b0110000001: data <= 14'h3fdd; 
        10'b0110000010: data <= 14'h3fc2; 
        10'b0110000011: data <= 14'h3fa5; 
        10'b0110000100: data <= 14'h3fbb; 
        10'b0110000101: data <= 14'h3ff4; 
        10'b0110000110: data <= 14'h3ff3; 
        10'b0110000111: data <= 14'h3ffe; 
        10'b0110001000: data <= 14'h3ffb; 
        10'b0110001001: data <= 14'h3ff4; 
        10'b0110001010: data <= 14'h3ffa; 
        10'b0110001011: data <= 14'h3ff1; 
        10'b0110001100: data <= 14'h3ffb; 
        10'b0110001101: data <= 14'h3ffa; 
        10'b0110001110: data <= 14'h0000; 
        10'b0110001111: data <= 14'h3ffd; 
        10'b0110010000: data <= 14'h001c; 
        10'b0110010001: data <= 14'h002c; 
        10'b0110010010: data <= 14'h0035; 
        10'b0110010011: data <= 14'h000a; 
        10'b0110010100: data <= 14'h0012; 
        10'b0110010101: data <= 14'h3ffd; 
        10'b0110010110: data <= 14'h3fda; 
        10'b0110010111: data <= 14'h3fd4; 
        10'b0110011000: data <= 14'h3fc3; 
        10'b0110011001: data <= 14'h3fca; 
        10'b0110011010: data <= 14'h3fce; 
        10'b0110011011: data <= 14'h3fe8; 
        10'b0110011100: data <= 14'h3feb; 
        10'b0110011101: data <= 14'h3fed; 
        10'b0110011110: data <= 14'h3ff4; 
        10'b0110011111: data <= 14'h3fce; 
        10'b0110100000: data <= 14'h3fde; 
        10'b0110100001: data <= 14'h3fef; 
        10'b0110100010: data <= 14'h3ffa; 
        10'b0110100011: data <= 14'h3ff1; 
        10'b0110100100: data <= 14'h3ff3; 
        10'b0110100101: data <= 14'h0002; 
        10'b0110100110: data <= 14'h3ff2; 
        10'b0110100111: data <= 14'h3ffa; 
        10'b0110101000: data <= 14'h3feb; 
        10'b0110101001: data <= 14'h3fe0; 
        10'b0110101010: data <= 14'h3fd3; 
        10'b0110101011: data <= 14'h3fe2; 
        10'b0110101100: data <= 14'h000b; 
        10'b0110101101: data <= 14'h0032; 
        10'b0110101110: data <= 14'h0018; 
        10'b0110101111: data <= 14'h0016; 
        10'b0110110000: data <= 14'h0013; 
        10'b0110110001: data <= 14'h3fef; 
        10'b0110110010: data <= 14'h3fc8; 
        10'b0110110011: data <= 14'h3fbf; 
        10'b0110110100: data <= 14'h3fc5; 
        10'b0110110101: data <= 14'h3fc4; 
        10'b0110110110: data <= 14'h3fd6; 
        10'b0110110111: data <= 14'h3ffe; 
        10'b0110111000: data <= 14'h3ff2; 
        10'b0110111001: data <= 14'h3ff4; 
        10'b0110111010: data <= 14'h3ff1; 
        10'b0110111011: data <= 14'h3fef; 
        10'b0110111100: data <= 14'h3ff4; 
        10'b0110111101: data <= 14'h0000; 
        10'b0110111110: data <= 14'h0002; 
        10'b0110111111: data <= 14'h3ff7; 
        10'b0111000000: data <= 14'h3ff8; 
        10'b0111000001: data <= 14'h3ffb; 
        10'b0111000010: data <= 14'h3ffd; 
        10'b0111000011: data <= 14'h3ff2; 
        10'b0111000100: data <= 14'h3ff8; 
        10'b0111000101: data <= 14'h3fdb; 
        10'b0111000110: data <= 14'h3fb7; 
        10'b0111000111: data <= 14'h3fa9; 
        10'b0111001000: data <= 14'h3fc5; 
        10'b0111001001: data <= 14'h3fe0; 
        10'b0111001010: data <= 14'h3ff3; 
        10'b0111001011: data <= 14'h3fed; 
        10'b0111001100: data <= 14'h3ff4; 
        10'b0111001101: data <= 14'h3fd8; 
        10'b0111001110: data <= 14'h3fb3; 
        10'b0111001111: data <= 14'h3fc1; 
        10'b0111010000: data <= 14'h3fd3; 
        10'b0111010001: data <= 14'h3ff0; 
        10'b0111010010: data <= 14'h3ff1; 
        10'b0111010011: data <= 14'h0002; 
        10'b0111010100: data <= 14'h000d; 
        10'b0111010101: data <= 14'h0002; 
        10'b0111010110: data <= 14'h000e; 
        10'b0111010111: data <= 14'h0003; 
        10'b0111011000: data <= 14'h0002; 
        10'b0111011001: data <= 14'h0002; 
        10'b0111011010: data <= 14'h3ff7; 
        10'b0111011011: data <= 14'h3ff8; 
        10'b0111011100: data <= 14'h3ff6; 
        10'b0111011101: data <= 14'h3fff; 
        10'b0111011110: data <= 14'h0000; 
        10'b0111011111: data <= 14'h0001; 
        10'b0111100000: data <= 14'h3ff7; 
        10'b0111100001: data <= 14'h0003; 
        10'b0111100010: data <= 14'h0005; 
        10'b0111100011: data <= 14'h3fc7; 
        10'b0111100100: data <= 14'h3f98; 
        10'b0111100101: data <= 14'h3f9f; 
        10'b0111100110: data <= 14'h3fba; 
        10'b0111100111: data <= 14'h3fd6; 
        10'b0111101000: data <= 14'h3fbf; 
        10'b0111101001: data <= 14'h3fac; 
        10'b0111101010: data <= 14'h3fae; 
        10'b0111101011: data <= 14'h3fdb; 
        10'b0111101100: data <= 14'h3ff0; 
        10'b0111101101: data <= 14'h0019; 
        10'b0111101110: data <= 14'h0026; 
        10'b0111101111: data <= 14'h0019; 
        10'b0111110000: data <= 14'h0019; 
        10'b0111110001: data <= 14'h0007; 
        10'b0111110010: data <= 14'h0001; 
        10'b0111110011: data <= 14'h000e; 
        10'b0111110100: data <= 14'h000e; 
        10'b0111110101: data <= 14'h3ff4; 
        10'b0111110110: data <= 14'h0000; 
        10'b0111110111: data <= 14'h0000; 
        10'b0111111000: data <= 14'h0001; 
        10'b0111111001: data <= 14'h3ff6; 
        10'b0111111010: data <= 14'h3ffa; 
        10'b0111111011: data <= 14'h3ff8; 
        10'b0111111100: data <= 14'h0015; 
        10'b0111111101: data <= 14'h001b; 
        10'b0111111110: data <= 14'h0040; 
        10'b0111111111: data <= 14'h000b; 
        10'b1000000000: data <= 14'h3fc2; 
        10'b1000000001: data <= 14'h3fa6; 
        10'b1000000010: data <= 14'h3f89; 
        10'b1000000011: data <= 14'h3f96; 
        10'b1000000100: data <= 14'h3fb4; 
        10'b1000000101: data <= 14'h3fd5; 
        10'b1000000110: data <= 14'h3fea; 
        10'b1000000111: data <= 14'h3ff7; 
        10'b1000001000: data <= 14'h3ffe; 
        10'b1000001001: data <= 14'h001d; 
        10'b1000001010: data <= 14'h000f; 
        10'b1000001011: data <= 14'h001a; 
        10'b1000001100: data <= 14'h0011; 
        10'b1000001101: data <= 14'h0019; 
        10'b1000001110: data <= 14'h0015; 
        10'b1000001111: data <= 14'h001d; 
        10'b1000010000: data <= 14'h000f; 
        10'b1000010001: data <= 14'h0001; 
        10'b1000010010: data <= 14'h3ff5; 
        10'b1000010011: data <= 14'h3ffc; 
        10'b1000010100: data <= 14'h0000; 
        10'b1000010101: data <= 14'h3ff6; 
        10'b1000010110: data <= 14'h3ffb; 
        10'b1000010111: data <= 14'h0002; 
        10'b1000011000: data <= 14'h001f; 
        10'b1000011001: data <= 14'h0035; 
        10'b1000011010: data <= 14'h0048; 
        10'b1000011011: data <= 14'h0030; 
        10'b1000011100: data <= 14'h001f; 
        10'b1000011101: data <= 14'h000a; 
        10'b1000011110: data <= 14'h3fe9; 
        10'b1000011111: data <= 14'h3fe8; 
        10'b1000100000: data <= 14'h0002; 
        10'b1000100001: data <= 14'h001d; 
        10'b1000100010: data <= 14'h000b; 
        10'b1000100011: data <= 14'h0010; 
        10'b1000100100: data <= 14'h0010; 
        10'b1000100101: data <= 14'h3ffb; 
        10'b1000100110: data <= 14'h000b; 
        10'b1000100111: data <= 14'h000b; 
        10'b1000101000: data <= 14'h0002; 
        10'b1000101001: data <= 14'h0013; 
        10'b1000101010: data <= 14'h0020; 
        10'b1000101011: data <= 14'h0018; 
        10'b1000101100: data <= 14'h0002; 
        10'b1000101101: data <= 14'h0000; 
        10'b1000101110: data <= 14'h0000; 
        10'b1000101111: data <= 14'h3ff3; 
        10'b1000110000: data <= 14'h3fff; 
        10'b1000110001: data <= 14'h3ff1; 
        10'b1000110010: data <= 14'h3ff9; 
        10'b1000110011: data <= 14'h3ff5; 
        10'b1000110100: data <= 14'h0004; 
        10'b1000110101: data <= 14'h0023; 
        10'b1000110110: data <= 14'h0029; 
        10'b1000110111: data <= 14'h0032; 
        10'b1000111000: data <= 14'h0045; 
        10'b1000111001: data <= 14'h003b; 
        10'b1000111010: data <= 14'h0033; 
        10'b1000111011: data <= 14'h004b; 
        10'b1000111100: data <= 14'h002f; 
        10'b1000111101: data <= 14'h0023; 
        10'b1000111110: data <= 14'h3ff6; 
        10'b1000111111: data <= 14'h3ff7; 
        10'b1001000000: data <= 14'h001a; 
        10'b1001000001: data <= 14'h000d; 
        10'b1001000010: data <= 14'h0016; 
        10'b1001000011: data <= 14'h001d; 
        10'b1001000100: data <= 14'h0019; 
        10'b1001000101: data <= 14'h0014; 
        10'b1001000110: data <= 14'h002f; 
        10'b1001000111: data <= 14'h0023; 
        10'b1001001000: data <= 14'h3ffb; 
        10'b1001001001: data <= 14'h3ff1; 
        10'b1001001010: data <= 14'h3ffb; 
        10'b1001001011: data <= 14'h3ff7; 
        10'b1001001100: data <= 14'h3ff5; 
        10'b1001001101: data <= 14'h0000; 
        10'b1001001110: data <= 14'h3ff1; 
        10'b1001001111: data <= 14'h3ffa; 
        10'b1001010000: data <= 14'h000e; 
        10'b1001010001: data <= 14'h3ffc; 
        10'b1001010010: data <= 14'h0011; 
        10'b1001010011: data <= 14'h002d; 
        10'b1001010100: data <= 14'h0041; 
        10'b1001010101: data <= 14'h002b; 
        10'b1001010110: data <= 14'h0024; 
        10'b1001010111: data <= 14'h0014; 
        10'b1001011000: data <= 14'h0019; 
        10'b1001011001: data <= 14'h0010; 
        10'b1001011010: data <= 14'h0010; 
        10'b1001011011: data <= 14'h0014; 
        10'b1001011100: data <= 14'h0005; 
        10'b1001011101: data <= 14'h0010; 
        10'b1001011110: data <= 14'h0008; 
        10'b1001011111: data <= 14'h001a; 
        10'b1001100000: data <= 14'h0019; 
        10'b1001100001: data <= 14'h002b; 
        10'b1001100010: data <= 14'h0034; 
        10'b1001100011: data <= 14'h000b; 
        10'b1001100100: data <= 14'h0000; 
        10'b1001100101: data <= 14'h3ff4; 
        10'b1001100110: data <= 14'h3ff7; 
        10'b1001100111: data <= 14'h3ff7; 
        10'b1001101000: data <= 14'h3ffd; 
        10'b1001101001: data <= 14'h3ff2; 
        10'b1001101010: data <= 14'h3ff9; 
        10'b1001101011: data <= 14'h3ff7; 
        10'b1001101100: data <= 14'h0005; 
        10'b1001101101: data <= 14'h3ff9; 
        10'b1001101110: data <= 14'h3ff1; 
        10'b1001101111: data <= 14'h3ffd; 
        10'b1001110000: data <= 14'h0019; 
        10'b1001110001: data <= 14'h0025; 
        10'b1001110010: data <= 14'h0006; 
        10'b1001110011: data <= 14'h0021; 
        10'b1001110100: data <= 14'h0035; 
        10'b1001110101: data <= 14'h0042; 
        10'b1001110110: data <= 14'h0021; 
        10'b1001110111: data <= 14'h0005; 
        10'b1001111000: data <= 14'h0004; 
        10'b1001111001: data <= 14'h0008; 
        10'b1001111010: data <= 14'h0011; 
        10'b1001111011: data <= 14'h0011; 
        10'b1001111100: data <= 14'h001d; 
        10'b1001111101: data <= 14'h001b; 
        10'b1001111110: data <= 14'h001c; 
        10'b1001111111: data <= 14'h000a; 
        10'b1010000000: data <= 14'h3fff; 
        10'b1010000001: data <= 14'h0002; 
        10'b1010000010: data <= 14'h3ffb; 
        10'b1010000011: data <= 14'h3ffc; 
        10'b1010000100: data <= 14'h3ff4; 
        10'b1010000101: data <= 14'h3ffa; 
        10'b1010000110: data <= 14'h3ffd; 
        10'b1010000111: data <= 14'h3ffb; 
        10'b1010001000: data <= 14'h3ff5; 
        10'b1010001001: data <= 14'h3ff9; 
        10'b1010001010: data <= 14'h3fea; 
        10'b1010001011: data <= 14'h3ff6; 
        10'b1010001100: data <= 14'h0014; 
        10'b1010001101: data <= 14'h0014; 
        10'b1010001110: data <= 14'h0014; 
        10'b1010001111: data <= 14'h0023; 
        10'b1010010000: data <= 14'h0022; 
        10'b1010010001: data <= 14'h0017; 
        10'b1010010010: data <= 14'h001a; 
        10'b1010010011: data <= 14'h0018; 
        10'b1010010100: data <= 14'h0018; 
        10'b1010010101: data <= 14'h000b; 
        10'b1010010110: data <= 14'h3ff3; 
        10'b1010010111: data <= 14'h3ffe; 
        10'b1010011000: data <= 14'h000c; 
        10'b1010011001: data <= 14'h0005; 
        10'b1010011010: data <= 14'h0010; 
        10'b1010011011: data <= 14'h3ff6; 
        10'b1010011100: data <= 14'h0003; 
        10'b1010011101: data <= 14'h3ff8; 
        10'b1010011110: data <= 14'h3ff8; 
        10'b1010011111: data <= 14'h0002; 
        10'b1010100000: data <= 14'h3fff; 
        10'b1010100001: data <= 14'h3ff8; 
        10'b1010100010: data <= 14'h3ff7; 
        10'b1010100011: data <= 14'h0003; 
        10'b1010100100: data <= 14'h3ff1; 
        10'b1010100101: data <= 14'h3ff0; 
        10'b1010100110: data <= 14'h3ffa; 
        10'b1010100111: data <= 14'h3ffd; 
        10'b1010101000: data <= 14'h3fff; 
        10'b1010101001: data <= 14'h001a; 
        10'b1010101010: data <= 14'h0022; 
        10'b1010101011: data <= 14'h001a; 
        10'b1010101100: data <= 14'h0011; 
        10'b1010101101: data <= 14'h0018; 
        10'b1010101110: data <= 14'h002b; 
        10'b1010101111: data <= 14'h0024; 
        10'b1010110000: data <= 14'h0015; 
        10'b1010110001: data <= 14'h000a; 
        10'b1010110010: data <= 14'h0014; 
        10'b1010110011: data <= 14'h000d; 
        10'b1010110100: data <= 14'h3fff; 
        10'b1010110101: data <= 14'h3ffe; 
        10'b1010110110: data <= 14'h3ffb; 
        10'b1010110111: data <= 14'h0001; 
        10'b1010111000: data <= 14'h3ff6; 
        10'b1010111001: data <= 14'h3ffc; 
        10'b1010111010: data <= 14'h0002; 
        10'b1010111011: data <= 14'h3ff3; 
        10'b1010111100: data <= 14'h3ffa; 
        10'b1010111101: data <= 14'h0001; 
        10'b1010111110: data <= 14'h0002; 
        10'b1010111111: data <= 14'h3ff3; 
        10'b1011000000: data <= 14'h0000; 
        10'b1011000001: data <= 14'h3ffc; 
        10'b1011000010: data <= 14'h3ff0; 
        10'b1011000011: data <= 14'h3ffa; 
        10'b1011000100: data <= 14'h3ff2; 
        10'b1011000101: data <= 14'h0008; 
        10'b1011000110: data <= 14'h0006; 
        10'b1011000111: data <= 14'h0012; 
        10'b1011001000: data <= 14'h0012; 
        10'b1011001001: data <= 14'h001f; 
        10'b1011001010: data <= 14'h0002; 
        10'b1011001011: data <= 14'h0009; 
        10'b1011001100: data <= 14'h0008; 
        10'b1011001101: data <= 14'h000f; 
        10'b1011001110: data <= 14'h3ff6; 
        10'b1011001111: data <= 14'h0000; 
        10'b1011010000: data <= 14'h3fef; 
        10'b1011010001: data <= 14'h0001; 
        10'b1011010010: data <= 14'h3ffa; 
        10'b1011010011: data <= 14'h3ff5; 
        10'b1011010100: data <= 14'h3fff; 
        10'b1011010101: data <= 14'h0001; 
        10'b1011010110: data <= 14'h3ff2; 
        10'b1011010111: data <= 14'h3ff8; 
        10'b1011011000: data <= 14'h3ffc; 
        10'b1011011001: data <= 14'h3ffb; 
        10'b1011011010: data <= 14'h3ff5; 
        10'b1011011011: data <= 14'h3ff8; 
        10'b1011011100: data <= 14'h3ff7; 
        10'b1011011101: data <= 14'h3ff9; 
        10'b1011011110: data <= 14'h3ffd; 
        10'b1011011111: data <= 14'h3ff6; 
        10'b1011100000: data <= 14'h3ff2; 
        10'b1011100001: data <= 14'h3ff9; 
        10'b1011100010: data <= 14'h3ff7; 
        10'b1011100011: data <= 14'h3ffe; 
        10'b1011100100: data <= 14'h0000; 
        10'b1011100101: data <= 14'h3ffc; 
        10'b1011100110: data <= 14'h3ff6; 
        10'b1011100111: data <= 14'h3ffb; 
        10'b1011101000: data <= 14'h3ffe; 
        10'b1011101001: data <= 14'h3ff6; 
        10'b1011101010: data <= 14'h3fec; 
        10'b1011101011: data <= 14'h3ff0; 
        10'b1011101100: data <= 14'h3ffd; 
        10'b1011101101: data <= 14'h3ffc; 
        10'b1011101110: data <= 14'h3ff7; 
        10'b1011101111: data <= 14'h3ffd; 
        10'b1011110000: data <= 14'h3ff9; 
        10'b1011110001: data <= 14'h3ffb; 
        10'b1011110010: data <= 14'h3ff7; 
        10'b1011110011: data <= 14'h3ff2; 
        10'b1011110100: data <= 14'h3ffd; 
        10'b1011110101: data <= 14'h3ffe; 
        10'b1011110110: data <= 14'h3fff; 
        10'b1011110111: data <= 14'h3ffc; 
        10'b1011111000: data <= 14'h3ff4; 
        10'b1011111001: data <= 14'h3fff; 
        10'b1011111010: data <= 14'h3ff8; 
        10'b1011111011: data <= 14'h3ff7; 
        10'b1011111100: data <= 14'h0003; 
        10'b1011111101: data <= 14'h3ff7; 
        10'b1011111110: data <= 14'h3ff6; 
        10'b1011111111: data <= 14'h3fff; 
        10'b1100000000: data <= 14'h3ffb; 
        10'b1100000001: data <= 14'h3ff1; 
        10'b1100000010: data <= 14'h0000; 
        10'b1100000011: data <= 14'h3ffb; 
        10'b1100000100: data <= 14'h3ff2; 
        10'b1100000101: data <= 14'h3ff1; 
        10'b1100000110: data <= 14'h3ff5; 
        10'b1100000111: data <= 14'h3ff1; 
        10'b1100001000: data <= 14'h0000; 
        10'b1100001001: data <= 14'h3ff8; 
        10'b1100001010: data <= 14'h0003; 
        10'b1100001011: data <= 14'h3ff3; 
        10'b1100001100: data <= 14'h3ffc; 
        10'b1100001101: data <= 14'h3ff9; 
        10'b1100001110: data <= 14'h3ff4; 
        10'b1100001111: data <= 14'h3ffe; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 9) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 15'h7fee; 
        10'b0000000001: data <= 15'h7ffd; 
        10'b0000000010: data <= 15'h7ffd; 
        10'b0000000011: data <= 15'h7fe8; 
        10'b0000000100: data <= 15'h7ff5; 
        10'b0000000101: data <= 15'h7ff2; 
        10'b0000000110: data <= 15'h0000; 
        10'b0000000111: data <= 15'h7ff1; 
        10'b0000001000: data <= 15'h7ffa; 
        10'b0000001001: data <= 15'h0005; 
        10'b0000001010: data <= 15'h7ffa; 
        10'b0000001011: data <= 15'h7ff9; 
        10'b0000001100: data <= 15'h7fee; 
        10'b0000001101: data <= 15'h7fff; 
        10'b0000001110: data <= 15'h7fe8; 
        10'b0000001111: data <= 15'h7fec; 
        10'b0000010000: data <= 15'h7fe5; 
        10'b0000010001: data <= 15'h7fea; 
        10'b0000010010: data <= 15'h7ffd; 
        10'b0000010011: data <= 15'h7ffa; 
        10'b0000010100: data <= 15'h7fe4; 
        10'b0000010101: data <= 15'h7ff5; 
        10'b0000010110: data <= 15'h7ff8; 
        10'b0000010111: data <= 15'h7ff2; 
        10'b0000011000: data <= 15'h7fe6; 
        10'b0000011001: data <= 15'h7ff6; 
        10'b0000011010: data <= 15'h7ff8; 
        10'b0000011011: data <= 15'h7fef; 
        10'b0000011100: data <= 15'h7ffe; 
        10'b0000011101: data <= 15'h7fe3; 
        10'b0000011110: data <= 15'h0000; 
        10'b0000011111: data <= 15'h7fe7; 
        10'b0000100000: data <= 15'h7fff; 
        10'b0000100001: data <= 15'h7ff0; 
        10'b0000100010: data <= 15'h7ff8; 
        10'b0000100011: data <= 15'h7fef; 
        10'b0000100100: data <= 15'h7feb; 
        10'b0000100101: data <= 15'h7ff8; 
        10'b0000100110: data <= 15'h0003; 
        10'b0000100111: data <= 15'h7fe8; 
        10'b0000101000: data <= 15'h7fef; 
        10'b0000101001: data <= 15'h7fea; 
        10'b0000101010: data <= 15'h7fe4; 
        10'b0000101011: data <= 15'h7ffb; 
        10'b0000101100: data <= 15'h7fed; 
        10'b0000101101: data <= 15'h7fea; 
        10'b0000101110: data <= 15'h7fee; 
        10'b0000101111: data <= 15'h7fec; 
        10'b0000110000: data <= 15'h7ffa; 
        10'b0000110001: data <= 15'h7fe7; 
        10'b0000110010: data <= 15'h0000; 
        10'b0000110011: data <= 15'h7fe8; 
        10'b0000110100: data <= 15'h0000; 
        10'b0000110101: data <= 15'h7ffe; 
        10'b0000110110: data <= 15'h7fe9; 
        10'b0000110111: data <= 15'h7ff3; 
        10'b0000111000: data <= 15'h7ff4; 
        10'b0000111001: data <= 15'h7ffb; 
        10'b0000111010: data <= 15'h7fef; 
        10'b0000111011: data <= 15'h7fe4; 
        10'b0000111100: data <= 15'h7fe9; 
        10'b0000111101: data <= 15'h7ff6; 
        10'b0000111110: data <= 15'h7fff; 
        10'b0000111111: data <= 15'h7ff8; 
        10'b0001000000: data <= 15'h7fec; 
        10'b0001000001: data <= 15'h7ff1; 
        10'b0001000010: data <= 15'h0004; 
        10'b0001000011: data <= 15'h7fe2; 
        10'b0001000100: data <= 15'h7fff; 
        10'b0001000101: data <= 15'h7feb; 
        10'b0001000110: data <= 15'h7fe5; 
        10'b0001000111: data <= 15'h7fea; 
        10'b0001001000: data <= 15'h7fee; 
        10'b0001001001: data <= 15'h7ff6; 
        10'b0001001010: data <= 15'h7ff1; 
        10'b0001001011: data <= 15'h7ff1; 
        10'b0001001100: data <= 15'h0007; 
        10'b0001001101: data <= 15'h0001; 
        10'b0001001110: data <= 15'h0003; 
        10'b0001001111: data <= 15'h7feb; 
        10'b0001010000: data <= 15'h7fe4; 
        10'b0001010001: data <= 15'h7ff2; 
        10'b0001010010: data <= 15'h7ffe; 
        10'b0001010011: data <= 15'h7ff8; 
        10'b0001010100: data <= 15'h7ffb; 
        10'b0001010101: data <= 15'h7ff8; 
        10'b0001010110: data <= 15'h7fe9; 
        10'b0001010111: data <= 15'h7fff; 
        10'b0001011000: data <= 15'h7fe7; 
        10'b0001011001: data <= 15'h7ff0; 
        10'b0001011010: data <= 15'h7fe2; 
        10'b0001011011: data <= 15'h7fed; 
        10'b0001011100: data <= 15'h7fe4; 
        10'b0001011101: data <= 15'h7fec; 
        10'b0001011110: data <= 15'h7fd0; 
        10'b0001011111: data <= 15'h7fc3; 
        10'b0001100000: data <= 15'h7fdd; 
        10'b0001100001: data <= 15'h7fdf; 
        10'b0001100010: data <= 15'h7fd8; 
        10'b0001100011: data <= 15'h7ff3; 
        10'b0001100100: data <= 15'h7ffa; 
        10'b0001100101: data <= 15'h7fe0; 
        10'b0001100110: data <= 15'h7fed; 
        10'b0001100111: data <= 15'h7ffa; 
        10'b0001101000: data <= 15'h7ffc; 
        10'b0001101001: data <= 15'h7ff3; 
        10'b0001101010: data <= 15'h7fe0; 
        10'b0001101011: data <= 15'h7fea; 
        10'b0001101100: data <= 15'h7fd9; 
        10'b0001101101: data <= 15'h0004; 
        10'b0001101110: data <= 15'h0003; 
        10'b0001101111: data <= 15'h7fe7; 
        10'b0001110000: data <= 15'h7fe5; 
        10'b0001110001: data <= 15'h7fef; 
        10'b0001110010: data <= 15'h0003; 
        10'b0001110011: data <= 15'h0001; 
        10'b0001110100: data <= 15'h0004; 
        10'b0001110101: data <= 15'h7fed; 
        10'b0001110110: data <= 15'h7feb; 
        10'b0001110111: data <= 15'h7fd5; 
        10'b0001111000: data <= 15'h7fb7; 
        10'b0001111001: data <= 15'h7f9f; 
        10'b0001111010: data <= 15'h7f73; 
        10'b0001111011: data <= 15'h7fa6; 
        10'b0001111100: data <= 15'h7fa5; 
        10'b0001111101: data <= 15'h7f86; 
        10'b0001111110: data <= 15'h7fbd; 
        10'b0001111111: data <= 15'h0000; 
        10'b0010000000: data <= 15'h7ff8; 
        10'b0010000001: data <= 15'h0017; 
        10'b0010000010: data <= 15'h7ff9; 
        10'b0010000011: data <= 15'h7fdd; 
        10'b0010000100: data <= 15'h7fd3; 
        10'b0010000101: data <= 15'h7fe8; 
        10'b0010000110: data <= 15'h7fec; 
        10'b0010000111: data <= 15'h7ff2; 
        10'b0010001000: data <= 15'h7fef; 
        10'b0010001001: data <= 15'h0006; 
        10'b0010001010: data <= 15'h0004; 
        10'b0010001011: data <= 15'h7ff3; 
        10'b0010001100: data <= 15'h7ff6; 
        10'b0010001101: data <= 15'h0006; 
        10'b0010001110: data <= 15'h7fea; 
        10'b0010001111: data <= 15'h7fe7; 
        10'b0010010000: data <= 15'h7fed; 
        10'b0010010001: data <= 15'h7fd4; 
        10'b0010010010: data <= 15'h7fbd; 
        10'b0010010011: data <= 15'h7fc0; 
        10'b0010010100: data <= 15'h7fd6; 
        10'b0010010101: data <= 15'h7ff8; 
        10'b0010010110: data <= 15'h000e; 
        10'b0010010111: data <= 15'h000f; 
        10'b0010011000: data <= 15'h7fe9; 
        10'b0010011001: data <= 15'h7fdf; 
        10'b0010011010: data <= 15'h7fec; 
        10'b0010011011: data <= 15'h7ff7; 
        10'b0010011100: data <= 15'h0021; 
        10'b0010011101: data <= 15'h0021; 
        10'b0010011110: data <= 15'h003f; 
        10'b0010011111: data <= 15'h0027; 
        10'b0010100000: data <= 15'h0026; 
        10'b0010100001: data <= 15'h0031; 
        10'b0010100010: data <= 15'h005b; 
        10'b0010100011: data <= 15'h004d; 
        10'b0010100100: data <= 15'h0036; 
        10'b0010100101: data <= 15'h001e; 
        10'b0010100110: data <= 15'h0013; 
        10'b0010100111: data <= 15'h0007; 
        10'b0010101000: data <= 15'h7fe8; 
        10'b0010101001: data <= 15'h7fe6; 
        10'b0010101010: data <= 15'h0003; 
        10'b0010101011: data <= 15'h7fe7; 
        10'b0010101100: data <= 15'h7fdf; 
        10'b0010101101: data <= 15'h7fb2; 
        10'b0010101110: data <= 15'h7fdd; 
        10'b0010101111: data <= 15'h7ffc; 
        10'b0010110000: data <= 15'h7ffd; 
        10'b0010110001: data <= 15'h0020; 
        10'b0010110010: data <= 15'h0042; 
        10'b0010110011: data <= 15'h0037; 
        10'b0010110100: data <= 15'h0009; 
        10'b0010110101: data <= 15'h0014; 
        10'b0010110110: data <= 15'h7ff7; 
        10'b0010110111: data <= 15'h7fe1; 
        10'b0010111000: data <= 15'h7fed; 
        10'b0010111001: data <= 15'h7ff0; 
        10'b0010111010: data <= 15'h0001; 
        10'b0010111011: data <= 15'h003e; 
        10'b0010111100: data <= 15'h0024; 
        10'b0010111101: data <= 15'h0028; 
        10'b0010111110: data <= 15'h007c; 
        10'b0010111111: data <= 15'h0095; 
        10'b0011000000: data <= 15'h00a7; 
        10'b0011000001: data <= 15'h0058; 
        10'b0011000010: data <= 15'h002c; 
        10'b0011000011: data <= 15'h000b; 
        10'b0011000100: data <= 15'h7ff2; 
        10'b0011000101: data <= 15'h7ff9; 
        10'b0011000110: data <= 15'h7ff5; 
        10'b0011000111: data <= 15'h7fe0; 
        10'b0011001000: data <= 15'h7fa6; 
        10'b0011001001: data <= 15'h7f96; 
        10'b0011001010: data <= 15'h7fbf; 
        10'b0011001011: data <= 15'h0008; 
        10'b0011001100: data <= 15'h002a; 
        10'b0011001101: data <= 15'h0053; 
        10'b0011001110: data <= 15'h0051; 
        10'b0011001111: data <= 15'h0047; 
        10'b0011010000: data <= 15'h0014; 
        10'b0011010001: data <= 15'h7ff9; 
        10'b0011010010: data <= 15'h7fe9; 
        10'b0011010011: data <= 15'h0002; 
        10'b0011010100: data <= 15'h0023; 
        10'b0011010101: data <= 15'h0020; 
        10'b0011010110: data <= 15'h0028; 
        10'b0011010111: data <= 15'h005a; 
        10'b0011011000: data <= 15'h004d; 
        10'b0011011001: data <= 15'h005d; 
        10'b0011011010: data <= 15'h0082; 
        10'b0011011011: data <= 15'h00ae; 
        10'b0011011100: data <= 15'h00d4; 
        10'b0011011101: data <= 15'h0099; 
        10'b0011011110: data <= 15'h0018; 
        10'b0011011111: data <= 15'h7ffc; 
        10'b0011100000: data <= 15'h7ffa; 
        10'b0011100001: data <= 15'h0006; 
        10'b0011100010: data <= 15'h0000; 
        10'b0011100011: data <= 15'h7fd4; 
        10'b0011100100: data <= 15'h7f7e; 
        10'b0011100101: data <= 15'h7f91; 
        10'b0011100110: data <= 15'h7faf; 
        10'b0011100111: data <= 15'h0005; 
        10'b0011101000: data <= 15'h003f; 
        10'b0011101001: data <= 15'h0013; 
        10'b0011101010: data <= 15'h0022; 
        10'b0011101011: data <= 15'h0042; 
        10'b0011101100: data <= 15'h0028; 
        10'b0011101101: data <= 15'h7fd3; 
        10'b0011101110: data <= 15'h7f9d; 
        10'b0011101111: data <= 15'h7fc4; 
        10'b0011110000: data <= 15'h7fdb; 
        10'b0011110001: data <= 15'h0004; 
        10'b0011110010: data <= 15'h000a; 
        10'b0011110011: data <= 15'h004b; 
        10'b0011110100: data <= 15'h004f; 
        10'b0011110101: data <= 15'h0070; 
        10'b0011110110: data <= 15'h00b1; 
        10'b0011110111: data <= 15'h00e8; 
        10'b0011111000: data <= 15'h0136; 
        10'b0011111001: data <= 15'h00c8; 
        10'b0011111010: data <= 15'h0024; 
        10'b0011111011: data <= 15'h7ffc; 
        10'b0011111100: data <= 15'h7fe6; 
        10'b0011111101: data <= 15'h7ff1; 
        10'b0011111110: data <= 15'h7fe4; 
        10'b0011111111: data <= 15'h7fc3; 
        10'b0100000000: data <= 15'h7fba; 
        10'b0100000001: data <= 15'h7fbf; 
        10'b0100000010: data <= 15'h0008; 
        10'b0100000011: data <= 15'h7ffb; 
        10'b0100000100: data <= 15'h0036; 
        10'b0100000101: data <= 15'h002f; 
        10'b0100000110: data <= 15'h0033; 
        10'b0100000111: data <= 15'h0088; 
        10'b0100001000: data <= 15'h0057; 
        10'b0100001001: data <= 15'h7fdc; 
        10'b0100001010: data <= 15'h7f89; 
        10'b0100001011: data <= 15'h7f55; 
        10'b0100001100: data <= 15'h7f60; 
        10'b0100001101: data <= 15'h7fa3; 
        10'b0100001110: data <= 15'h7feb; 
        10'b0100001111: data <= 15'h7fff; 
        10'b0100010000: data <= 15'h0049; 
        10'b0100010001: data <= 15'h009b; 
        10'b0100010010: data <= 15'h00e0; 
        10'b0100010011: data <= 15'h0133; 
        10'b0100010100: data <= 15'h0182; 
        10'b0100010101: data <= 15'h00fe; 
        10'b0100010110: data <= 15'h002d; 
        10'b0100010111: data <= 15'h7fee; 
        10'b0100011000: data <= 15'h7ffa; 
        10'b0100011001: data <= 15'h7fee; 
        10'b0100011010: data <= 15'h7fe8; 
        10'b0100011011: data <= 15'h7fed; 
        10'b0100011100: data <= 15'h7fec; 
        10'b0100011101: data <= 15'h7ff3; 
        10'b0100011110: data <= 15'h002b; 
        10'b0100011111: data <= 15'h0051; 
        10'b0100100000: data <= 15'h007e; 
        10'b0100100001: data <= 15'h008b; 
        10'b0100100010: data <= 15'h0085; 
        10'b0100100011: data <= 15'h00a1; 
        10'b0100100100: data <= 15'h0086; 
        10'b0100100101: data <= 15'h0067; 
        10'b0100100110: data <= 15'h7fea; 
        10'b0100100111: data <= 15'h7fac; 
        10'b0100101000: data <= 15'h7f73; 
        10'b0100101001: data <= 15'h7f78; 
        10'b0100101010: data <= 15'h7f73; 
        10'b0100101011: data <= 15'h7f5f; 
        10'b0100101100: data <= 15'h7f92; 
        10'b0100101101: data <= 15'h7fde; 
        10'b0100101110: data <= 15'h0013; 
        10'b0100101111: data <= 15'h0067; 
        10'b0100110000: data <= 15'h00ce; 
        10'b0100110001: data <= 15'h009b; 
        10'b0100110010: data <= 15'h0035; 
        10'b0100110011: data <= 15'h7fee; 
        10'b0100110100: data <= 15'h7fe8; 
        10'b0100110101: data <= 15'h0000; 
        10'b0100110110: data <= 15'h7fec; 
        10'b0100110111: data <= 15'h7ff3; 
        10'b0100111000: data <= 15'h7fec; 
        10'b0100111001: data <= 15'h7ffd; 
        10'b0100111010: data <= 15'h0045; 
        10'b0100111011: data <= 15'h0054; 
        10'b0100111100: data <= 15'h0079; 
        10'b0100111101: data <= 15'h0070; 
        10'b0100111110: data <= 15'h0052; 
        10'b0100111111: data <= 15'h005a; 
        10'b0101000000: data <= 15'h0096; 
        10'b0101000001: data <= 15'h008c; 
        10'b0101000010: data <= 15'h0002; 
        10'b0101000011: data <= 15'h7fa9; 
        10'b0101000100: data <= 15'h7f94; 
        10'b0101000101: data <= 15'h7f8c; 
        10'b0101000110: data <= 15'h7f65; 
        10'b0101000111: data <= 15'h7f27; 
        10'b0101001000: data <= 15'h7ec6; 
        10'b0101001001: data <= 15'h7edf; 
        10'b0101001010: data <= 15'h7f13; 
        10'b0101001011: data <= 15'h7f54; 
        10'b0101001100: data <= 15'h7fc3; 
        10'b0101001101: data <= 15'h0007; 
        10'b0101001110: data <= 15'h0011; 
        10'b0101001111: data <= 15'h7ff6; 
        10'b0101010000: data <= 15'h7ff5; 
        10'b0101010001: data <= 15'h7ff7; 
        10'b0101010010: data <= 15'h7ff3; 
        10'b0101010011: data <= 15'h7fee; 
        10'b0101010100: data <= 15'h7ff2; 
        10'b0101010101: data <= 15'h0023; 
        10'b0101010110: data <= 15'h004f; 
        10'b0101010111: data <= 15'h0046; 
        10'b0101011000: data <= 15'h0034; 
        10'b0101011001: data <= 15'h001e; 
        10'b0101011010: data <= 15'h0057; 
        10'b0101011011: data <= 15'h00b5; 
        10'b0101011100: data <= 15'h00a9; 
        10'b0101011101: data <= 15'h00ad; 
        10'b0101011110: data <= 15'h0012; 
        10'b0101011111: data <= 15'h7fa8; 
        10'b0101100000: data <= 15'h7f5c; 
        10'b0101100001: data <= 15'h7f7c; 
        10'b0101100010: data <= 15'h7fa6; 
        10'b0101100011: data <= 15'h7f7f; 
        10'b0101100100: data <= 15'h7f6d; 
        10'b0101100101: data <= 15'h7f0c; 
        10'b0101100110: data <= 15'h7eea; 
        10'b0101100111: data <= 15'h7f0e; 
        10'b0101101000: data <= 15'h7f5e; 
        10'b0101101001: data <= 15'h7fd2; 
        10'b0101101010: data <= 15'h0002; 
        10'b0101101011: data <= 15'h0000; 
        10'b0101101100: data <= 15'h7ff6; 
        10'b0101101101: data <= 15'h7fe9; 
        10'b0101101110: data <= 15'h7fe8; 
        10'b0101101111: data <= 15'h7fef; 
        10'b0101110000: data <= 15'h7ffb; 
        10'b0101110001: data <= 15'h0012; 
        10'b0101110010: data <= 15'h0035; 
        10'b0101110011: data <= 15'h0027; 
        10'b0101110100: data <= 15'h002d; 
        10'b0101110101: data <= 15'h0025; 
        10'b0101110110: data <= 15'h007a; 
        10'b0101110111: data <= 15'h0088; 
        10'b0101111000: data <= 15'h0065; 
        10'b0101111001: data <= 15'h005f; 
        10'b0101111010: data <= 15'h7fed; 
        10'b0101111011: data <= 15'h7f97; 
        10'b0101111100: data <= 15'h7f56; 
        10'b0101111101: data <= 15'h7fa6; 
        10'b0101111110: data <= 15'h7fe0; 
        10'b0101111111: data <= 15'h7fdb; 
        10'b0110000000: data <= 15'h7fee; 
        10'b0110000001: data <= 15'h7fbb; 
        10'b0110000010: data <= 15'h7f83; 
        10'b0110000011: data <= 15'h7f49; 
        10'b0110000100: data <= 15'h7f77; 
        10'b0110000101: data <= 15'h7fe8; 
        10'b0110000110: data <= 15'h7fe6; 
        10'b0110000111: data <= 15'h7ffc; 
        10'b0110001000: data <= 15'h7ff7; 
        10'b0110001001: data <= 15'h7fe7; 
        10'b0110001010: data <= 15'h7ff4; 
        10'b0110001011: data <= 15'h7fe1; 
        10'b0110001100: data <= 15'h7ff6; 
        10'b0110001101: data <= 15'h7ff5; 
        10'b0110001110: data <= 15'h7fff; 
        10'b0110001111: data <= 15'h7ffa; 
        10'b0110010000: data <= 15'h0038; 
        10'b0110010001: data <= 15'h0059; 
        10'b0110010010: data <= 15'h006a; 
        10'b0110010011: data <= 15'h0014; 
        10'b0110010100: data <= 15'h0024; 
        10'b0110010101: data <= 15'h7ff9; 
        10'b0110010110: data <= 15'h7fb4; 
        10'b0110010111: data <= 15'h7fa8; 
        10'b0110011000: data <= 15'h7f86; 
        10'b0110011001: data <= 15'h7f95; 
        10'b0110011010: data <= 15'h7f9b; 
        10'b0110011011: data <= 15'h7fcf; 
        10'b0110011100: data <= 15'h7fd6; 
        10'b0110011101: data <= 15'h7fda; 
        10'b0110011110: data <= 15'h7fe9; 
        10'b0110011111: data <= 15'h7f9c; 
        10'b0110100000: data <= 15'h7fbd; 
        10'b0110100001: data <= 15'h7fde; 
        10'b0110100010: data <= 15'h7ff4; 
        10'b0110100011: data <= 15'h7fe2; 
        10'b0110100100: data <= 15'h7fe5; 
        10'b0110100101: data <= 15'h0004; 
        10'b0110100110: data <= 15'h7fe3; 
        10'b0110100111: data <= 15'h7ff4; 
        10'b0110101000: data <= 15'h7fd5; 
        10'b0110101001: data <= 15'h7fc0; 
        10'b0110101010: data <= 15'h7fa6; 
        10'b0110101011: data <= 15'h7fc4; 
        10'b0110101100: data <= 15'h0016; 
        10'b0110101101: data <= 15'h0064; 
        10'b0110101110: data <= 15'h002f; 
        10'b0110101111: data <= 15'h002c; 
        10'b0110110000: data <= 15'h0026; 
        10'b0110110001: data <= 15'h7fde; 
        10'b0110110010: data <= 15'h7f8f; 
        10'b0110110011: data <= 15'h7f7e; 
        10'b0110110100: data <= 15'h7f8b; 
        10'b0110110101: data <= 15'h7f88; 
        10'b0110110110: data <= 15'h7fab; 
        10'b0110110111: data <= 15'h7ffc; 
        10'b0110111000: data <= 15'h7fe3; 
        10'b0110111001: data <= 15'h7fe8; 
        10'b0110111010: data <= 15'h7fe3; 
        10'b0110111011: data <= 15'h7fdf; 
        10'b0110111100: data <= 15'h7fe9; 
        10'b0110111101: data <= 15'h7fff; 
        10'b0110111110: data <= 15'h0005; 
        10'b0110111111: data <= 15'h7fee; 
        10'b0111000000: data <= 15'h7ff0; 
        10'b0111000001: data <= 15'h7ff6; 
        10'b0111000010: data <= 15'h7ff9; 
        10'b0111000011: data <= 15'h7fe3; 
        10'b0111000100: data <= 15'h7fef; 
        10'b0111000101: data <= 15'h7fb7; 
        10'b0111000110: data <= 15'h7f6d; 
        10'b0111000111: data <= 15'h7f52; 
        10'b0111001000: data <= 15'h7f8b; 
        10'b0111001001: data <= 15'h7fbf; 
        10'b0111001010: data <= 15'h7fe6; 
        10'b0111001011: data <= 15'h7fdb; 
        10'b0111001100: data <= 15'h7fe8; 
        10'b0111001101: data <= 15'h7fb0; 
        10'b0111001110: data <= 15'h7f66; 
        10'b0111001111: data <= 15'h7f83; 
        10'b0111010000: data <= 15'h7fa5; 
        10'b0111010001: data <= 15'h7fdf; 
        10'b0111010010: data <= 15'h7fe1; 
        10'b0111010011: data <= 15'h0005; 
        10'b0111010100: data <= 15'h0019; 
        10'b0111010101: data <= 15'h0004; 
        10'b0111010110: data <= 15'h001c; 
        10'b0111010111: data <= 15'h0006; 
        10'b0111011000: data <= 15'h0004; 
        10'b0111011001: data <= 15'h0004; 
        10'b0111011010: data <= 15'h7fef; 
        10'b0111011011: data <= 15'h7ff0; 
        10'b0111011100: data <= 15'h7fed; 
        10'b0111011101: data <= 15'h7fff; 
        10'b0111011110: data <= 15'h0000; 
        10'b0111011111: data <= 15'h0002; 
        10'b0111100000: data <= 15'h7fed; 
        10'b0111100001: data <= 15'h0005; 
        10'b0111100010: data <= 15'h000b; 
        10'b0111100011: data <= 15'h7f8d; 
        10'b0111100100: data <= 15'h7f31; 
        10'b0111100101: data <= 15'h7f3e; 
        10'b0111100110: data <= 15'h7f75; 
        10'b0111100111: data <= 15'h7fac; 
        10'b0111101000: data <= 15'h7f7d; 
        10'b0111101001: data <= 15'h7f57; 
        10'b0111101010: data <= 15'h7f5c; 
        10'b0111101011: data <= 15'h7fb5; 
        10'b0111101100: data <= 15'h7fdf; 
        10'b0111101101: data <= 15'h0032; 
        10'b0111101110: data <= 15'h004c; 
        10'b0111101111: data <= 15'h0032; 
        10'b0111110000: data <= 15'h0032; 
        10'b0111110001: data <= 15'h000f; 
        10'b0111110010: data <= 15'h0002; 
        10'b0111110011: data <= 15'h001c; 
        10'b0111110100: data <= 15'h001c; 
        10'b0111110101: data <= 15'h7fe8; 
        10'b0111110110: data <= 15'h7fff; 
        10'b0111110111: data <= 15'h0001; 
        10'b0111111000: data <= 15'h0003; 
        10'b0111111001: data <= 15'h7fec; 
        10'b0111111010: data <= 15'h7ff3; 
        10'b0111111011: data <= 15'h7ff0; 
        10'b0111111100: data <= 15'h0029; 
        10'b0111111101: data <= 15'h0036; 
        10'b0111111110: data <= 15'h0081; 
        10'b0111111111: data <= 15'h0017; 
        10'b1000000000: data <= 15'h7f84; 
        10'b1000000001: data <= 15'h7f4b; 
        10'b1000000010: data <= 15'h7f12; 
        10'b1000000011: data <= 15'h7f2c; 
        10'b1000000100: data <= 15'h7f68; 
        10'b1000000101: data <= 15'h7fa9; 
        10'b1000000110: data <= 15'h7fd5; 
        10'b1000000111: data <= 15'h7fee; 
        10'b1000001000: data <= 15'h7ffd; 
        10'b1000001001: data <= 15'h003a; 
        10'b1000001010: data <= 15'h001d; 
        10'b1000001011: data <= 15'h0034; 
        10'b1000001100: data <= 15'h0023; 
        10'b1000001101: data <= 15'h0033; 
        10'b1000001110: data <= 15'h002a; 
        10'b1000001111: data <= 15'h003a; 
        10'b1000010000: data <= 15'h001e; 
        10'b1000010001: data <= 15'h0002; 
        10'b1000010010: data <= 15'h7fea; 
        10'b1000010011: data <= 15'h7ff9; 
        10'b1000010100: data <= 15'h0000; 
        10'b1000010101: data <= 15'h7fec; 
        10'b1000010110: data <= 15'h7ff5; 
        10'b1000010111: data <= 15'h0004; 
        10'b1000011000: data <= 15'h003e; 
        10'b1000011001: data <= 15'h006a; 
        10'b1000011010: data <= 15'h008f; 
        10'b1000011011: data <= 15'h0060; 
        10'b1000011100: data <= 15'h003d; 
        10'b1000011101: data <= 15'h0014; 
        10'b1000011110: data <= 15'h7fd2; 
        10'b1000011111: data <= 15'h7fcf; 
        10'b1000100000: data <= 15'h0004; 
        10'b1000100001: data <= 15'h003a; 
        10'b1000100010: data <= 15'h0016; 
        10'b1000100011: data <= 15'h001f; 
        10'b1000100100: data <= 15'h001f; 
        10'b1000100101: data <= 15'h7ff6; 
        10'b1000100110: data <= 15'h0017; 
        10'b1000100111: data <= 15'h0016; 
        10'b1000101000: data <= 15'h0005; 
        10'b1000101001: data <= 15'h0026; 
        10'b1000101010: data <= 15'h0041; 
        10'b1000101011: data <= 15'h002f; 
        10'b1000101100: data <= 15'h0004; 
        10'b1000101101: data <= 15'h7fff; 
        10'b1000101110: data <= 15'h0000; 
        10'b1000101111: data <= 15'h7fe6; 
        10'b1000110000: data <= 15'h7fff; 
        10'b1000110001: data <= 15'h7fe2; 
        10'b1000110010: data <= 15'h7ff2; 
        10'b1000110011: data <= 15'h7fea; 
        10'b1000110100: data <= 15'h0008; 
        10'b1000110101: data <= 15'h0046; 
        10'b1000110110: data <= 15'h0051; 
        10'b1000110111: data <= 15'h0063; 
        10'b1000111000: data <= 15'h008b; 
        10'b1000111001: data <= 15'h0075; 
        10'b1000111010: data <= 15'h0067; 
        10'b1000111011: data <= 15'h0096; 
        10'b1000111100: data <= 15'h005d; 
        10'b1000111101: data <= 15'h0046; 
        10'b1000111110: data <= 15'h7fec; 
        10'b1000111111: data <= 15'h7fee; 
        10'b1001000000: data <= 15'h0034; 
        10'b1001000001: data <= 15'h001a; 
        10'b1001000010: data <= 15'h002b; 
        10'b1001000011: data <= 15'h0039; 
        10'b1001000100: data <= 15'h0032; 
        10'b1001000101: data <= 15'h0027; 
        10'b1001000110: data <= 15'h005e; 
        10'b1001000111: data <= 15'h0046; 
        10'b1001001000: data <= 15'h7ff7; 
        10'b1001001001: data <= 15'h7fe3; 
        10'b1001001010: data <= 15'h7ff6; 
        10'b1001001011: data <= 15'h7fed; 
        10'b1001001100: data <= 15'h7feb; 
        10'b1001001101: data <= 15'h0001; 
        10'b1001001110: data <= 15'h7fe1; 
        10'b1001001111: data <= 15'h7ff4; 
        10'b1001010000: data <= 15'h001c; 
        10'b1001010001: data <= 15'h7ff7; 
        10'b1001010010: data <= 15'h0021; 
        10'b1001010011: data <= 15'h005b; 
        10'b1001010100: data <= 15'h0083; 
        10'b1001010101: data <= 15'h0056; 
        10'b1001010110: data <= 15'h0049; 
        10'b1001010111: data <= 15'h0027; 
        10'b1001011000: data <= 15'h0033; 
        10'b1001011001: data <= 15'h001f; 
        10'b1001011010: data <= 15'h0021; 
        10'b1001011011: data <= 15'h0028; 
        10'b1001011100: data <= 15'h000a; 
        10'b1001011101: data <= 15'h0020; 
        10'b1001011110: data <= 15'h0010; 
        10'b1001011111: data <= 15'h0034; 
        10'b1001100000: data <= 15'h0033; 
        10'b1001100001: data <= 15'h0055; 
        10'b1001100010: data <= 15'h0069; 
        10'b1001100011: data <= 15'h0017; 
        10'b1001100100: data <= 15'h0001; 
        10'b1001100101: data <= 15'h7fe7; 
        10'b1001100110: data <= 15'h7fee; 
        10'b1001100111: data <= 15'h7fee; 
        10'b1001101000: data <= 15'h7ffa; 
        10'b1001101001: data <= 15'h7fe4; 
        10'b1001101010: data <= 15'h7ff1; 
        10'b1001101011: data <= 15'h7fee; 
        10'b1001101100: data <= 15'h000a; 
        10'b1001101101: data <= 15'h7ff2; 
        10'b1001101110: data <= 15'h7fe1; 
        10'b1001101111: data <= 15'h7ffb; 
        10'b1001110000: data <= 15'h0033; 
        10'b1001110001: data <= 15'h004a; 
        10'b1001110010: data <= 15'h000d; 
        10'b1001110011: data <= 15'h0042; 
        10'b1001110100: data <= 15'h006a; 
        10'b1001110101: data <= 15'h0083; 
        10'b1001110110: data <= 15'h0043; 
        10'b1001110111: data <= 15'h000a; 
        10'b1001111000: data <= 15'h0007; 
        10'b1001111001: data <= 15'h0010; 
        10'b1001111010: data <= 15'h0022; 
        10'b1001111011: data <= 15'h0022; 
        10'b1001111100: data <= 15'h003b; 
        10'b1001111101: data <= 15'h0035; 
        10'b1001111110: data <= 15'h0037; 
        10'b1001111111: data <= 15'h0013; 
        10'b1010000000: data <= 15'h7ffd; 
        10'b1010000001: data <= 15'h0003; 
        10'b1010000010: data <= 15'h7ff5; 
        10'b1010000011: data <= 15'h7ff9; 
        10'b1010000100: data <= 15'h7fe9; 
        10'b1010000101: data <= 15'h7ff5; 
        10'b1010000110: data <= 15'h7ff9; 
        10'b1010000111: data <= 15'h7ff7; 
        10'b1010001000: data <= 15'h7fea; 
        10'b1010001001: data <= 15'h7ff1; 
        10'b1010001010: data <= 15'h7fd4; 
        10'b1010001011: data <= 15'h7fec; 
        10'b1010001100: data <= 15'h0028; 
        10'b1010001101: data <= 15'h0027; 
        10'b1010001110: data <= 15'h0027; 
        10'b1010001111: data <= 15'h0046; 
        10'b1010010000: data <= 15'h0043; 
        10'b1010010001: data <= 15'h002e; 
        10'b1010010010: data <= 15'h0035; 
        10'b1010010011: data <= 15'h0030; 
        10'b1010010100: data <= 15'h002f; 
        10'b1010010101: data <= 15'h0016; 
        10'b1010010110: data <= 15'h7fe7; 
        10'b1010010111: data <= 15'h7ffc; 
        10'b1010011000: data <= 15'h0017; 
        10'b1010011001: data <= 15'h0009; 
        10'b1010011010: data <= 15'h001f; 
        10'b1010011011: data <= 15'h7fed; 
        10'b1010011100: data <= 15'h0005; 
        10'b1010011101: data <= 15'h7ff0; 
        10'b1010011110: data <= 15'h7ff0; 
        10'b1010011111: data <= 15'h0005; 
        10'b1010100000: data <= 15'h7ffe; 
        10'b1010100001: data <= 15'h7ff1; 
        10'b1010100010: data <= 15'h7fee; 
        10'b1010100011: data <= 15'h0005; 
        10'b1010100100: data <= 15'h7fe2; 
        10'b1010100101: data <= 15'h7fe0; 
        10'b1010100110: data <= 15'h7ff4; 
        10'b1010100111: data <= 15'h7ffa; 
        10'b1010101000: data <= 15'h7ffe; 
        10'b1010101001: data <= 15'h0034; 
        10'b1010101010: data <= 15'h0044; 
        10'b1010101011: data <= 15'h0034; 
        10'b1010101100: data <= 15'h0022; 
        10'b1010101101: data <= 15'h002f; 
        10'b1010101110: data <= 15'h0057; 
        10'b1010101111: data <= 15'h0048; 
        10'b1010110000: data <= 15'h002b; 
        10'b1010110001: data <= 15'h0015; 
        10'b1010110010: data <= 15'h0028; 
        10'b1010110011: data <= 15'h001a; 
        10'b1010110100: data <= 15'h7fff; 
        10'b1010110101: data <= 15'h7ffc; 
        10'b1010110110: data <= 15'h7ff7; 
        10'b1010110111: data <= 15'h0002; 
        10'b1010111000: data <= 15'h7feb; 
        10'b1010111001: data <= 15'h7ff8; 
        10'b1010111010: data <= 15'h0003; 
        10'b1010111011: data <= 15'h7fe6; 
        10'b1010111100: data <= 15'h7ff5; 
        10'b1010111101: data <= 15'h0001; 
        10'b1010111110: data <= 15'h0003; 
        10'b1010111111: data <= 15'h7fe5; 
        10'b1011000000: data <= 15'h0000; 
        10'b1011000001: data <= 15'h7ff8; 
        10'b1011000010: data <= 15'h7fe0; 
        10'b1011000011: data <= 15'h7ff4; 
        10'b1011000100: data <= 15'h7fe3; 
        10'b1011000101: data <= 15'h0011; 
        10'b1011000110: data <= 15'h000d; 
        10'b1011000111: data <= 15'h0023; 
        10'b1011001000: data <= 15'h0023; 
        10'b1011001001: data <= 15'h003d; 
        10'b1011001010: data <= 15'h0003; 
        10'b1011001011: data <= 15'h0012; 
        10'b1011001100: data <= 15'h000f; 
        10'b1011001101: data <= 15'h001e; 
        10'b1011001110: data <= 15'h7fec; 
        10'b1011001111: data <= 15'h7fff; 
        10'b1011010000: data <= 15'h7fde; 
        10'b1011010001: data <= 15'h0003; 
        10'b1011010010: data <= 15'h7ff3; 
        10'b1011010011: data <= 15'h7fe9; 
        10'b1011010100: data <= 15'h7ffd; 
        10'b1011010101: data <= 15'h0002; 
        10'b1011010110: data <= 15'h7fe3; 
        10'b1011010111: data <= 15'h7ff1; 
        10'b1011011000: data <= 15'h7ff7; 
        10'b1011011001: data <= 15'h7ff6; 
        10'b1011011010: data <= 15'h7feb; 
        10'b1011011011: data <= 15'h7ff0; 
        10'b1011011100: data <= 15'h7fee; 
        10'b1011011101: data <= 15'h7ff1; 
        10'b1011011110: data <= 15'h7ffb; 
        10'b1011011111: data <= 15'h7feb; 
        10'b1011100000: data <= 15'h7fe4; 
        10'b1011100001: data <= 15'h7ff2; 
        10'b1011100010: data <= 15'h7fed; 
        10'b1011100011: data <= 15'h7ffc; 
        10'b1011100100: data <= 15'h0001; 
        10'b1011100101: data <= 15'h7ff9; 
        10'b1011100110: data <= 15'h7fec; 
        10'b1011100111: data <= 15'h7ff6; 
        10'b1011101000: data <= 15'h7ffb; 
        10'b1011101001: data <= 15'h7feb; 
        10'b1011101010: data <= 15'h7fd8; 
        10'b1011101011: data <= 15'h7fdf; 
        10'b1011101100: data <= 15'h7ff9; 
        10'b1011101101: data <= 15'h7ff9; 
        10'b1011101110: data <= 15'h7fee; 
        10'b1011101111: data <= 15'h7ffb; 
        10'b1011110000: data <= 15'h7ff2; 
        10'b1011110001: data <= 15'h7ff7; 
        10'b1011110010: data <= 15'h7fef; 
        10'b1011110011: data <= 15'h7fe3; 
        10'b1011110100: data <= 15'h7ffa; 
        10'b1011110101: data <= 15'h7ffc; 
        10'b1011110110: data <= 15'h7ffd; 
        10'b1011110111: data <= 15'h7ff8; 
        10'b1011111000: data <= 15'h7fe8; 
        10'b1011111001: data <= 15'h7ffe; 
        10'b1011111010: data <= 15'h7ff0; 
        10'b1011111011: data <= 15'h7fee; 
        10'b1011111100: data <= 15'h0006; 
        10'b1011111101: data <= 15'h7fef; 
        10'b1011111110: data <= 15'h7fec; 
        10'b1011111111: data <= 15'h7ffe; 
        10'b1100000000: data <= 15'h7ff5; 
        10'b1100000001: data <= 15'h7fe2; 
        10'b1100000010: data <= 15'h0001; 
        10'b1100000011: data <= 15'h7ff7; 
        10'b1100000100: data <= 15'h7fe5; 
        10'b1100000101: data <= 15'h7fe2; 
        10'b1100000110: data <= 15'h7fe9; 
        10'b1100000111: data <= 15'h7fe1; 
        10'b1100001000: data <= 15'h0000; 
        10'b1100001001: data <= 15'h7fef; 
        10'b1100001010: data <= 15'h0006; 
        10'b1100001011: data <= 15'h7fe6; 
        10'b1100001100: data <= 15'h7ff8; 
        10'b1100001101: data <= 15'h7ff3; 
        10'b1100001110: data <= 15'h7fe8; 
        10'b1100001111: data <= 15'h7ffc; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 10) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 16'hffdd; 
        10'b0000000001: data <= 16'hfffb; 
        10'b0000000010: data <= 16'hfffb; 
        10'b0000000011: data <= 16'hffd0; 
        10'b0000000100: data <= 16'hffea; 
        10'b0000000101: data <= 16'hffe4; 
        10'b0000000110: data <= 16'h0000; 
        10'b0000000111: data <= 16'hffe1; 
        10'b0000001000: data <= 16'hfff3; 
        10'b0000001001: data <= 16'h000a; 
        10'b0000001010: data <= 16'hfff3; 
        10'b0000001011: data <= 16'hfff2; 
        10'b0000001100: data <= 16'hffdc; 
        10'b0000001101: data <= 16'hfffe; 
        10'b0000001110: data <= 16'hffcf; 
        10'b0000001111: data <= 16'hffd8; 
        10'b0000010000: data <= 16'hffc9; 
        10'b0000010001: data <= 16'hffd3; 
        10'b0000010010: data <= 16'hfff9; 
        10'b0000010011: data <= 16'hfff4; 
        10'b0000010100: data <= 16'hffc8; 
        10'b0000010101: data <= 16'hffeb; 
        10'b0000010110: data <= 16'hfff1; 
        10'b0000010111: data <= 16'hffe5; 
        10'b0000011000: data <= 16'hffcc; 
        10'b0000011001: data <= 16'hffec; 
        10'b0000011010: data <= 16'hfff1; 
        10'b0000011011: data <= 16'hffde; 
        10'b0000011100: data <= 16'hfffd; 
        10'b0000011101: data <= 16'hffc6; 
        10'b0000011110: data <= 16'h0000; 
        10'b0000011111: data <= 16'hffce; 
        10'b0000100000: data <= 16'hfffe; 
        10'b0000100001: data <= 16'hffe0; 
        10'b0000100010: data <= 16'hfff0; 
        10'b0000100011: data <= 16'hffdf; 
        10'b0000100100: data <= 16'hffd6; 
        10'b0000100101: data <= 16'hfff1; 
        10'b0000100110: data <= 16'h0005; 
        10'b0000100111: data <= 16'hffcf; 
        10'b0000101000: data <= 16'hffde; 
        10'b0000101001: data <= 16'hffd5; 
        10'b0000101010: data <= 16'hffc8; 
        10'b0000101011: data <= 16'hfff7; 
        10'b0000101100: data <= 16'hffda; 
        10'b0000101101: data <= 16'hffd4; 
        10'b0000101110: data <= 16'hffdb; 
        10'b0000101111: data <= 16'hffd9; 
        10'b0000110000: data <= 16'hfff4; 
        10'b0000110001: data <= 16'hffcd; 
        10'b0000110010: data <= 16'hffff; 
        10'b0000110011: data <= 16'hffd1; 
        10'b0000110100: data <= 16'h0001; 
        10'b0000110101: data <= 16'hfffc; 
        10'b0000110110: data <= 16'hffd3; 
        10'b0000110111: data <= 16'hffe7; 
        10'b0000111000: data <= 16'hffe8; 
        10'b0000111001: data <= 16'hfff5; 
        10'b0000111010: data <= 16'hffde; 
        10'b0000111011: data <= 16'hffc8; 
        10'b0000111100: data <= 16'hffd2; 
        10'b0000111101: data <= 16'hffed; 
        10'b0000111110: data <= 16'hfffe; 
        10'b0000111111: data <= 16'hfff1; 
        10'b0001000000: data <= 16'hffd8; 
        10'b0001000001: data <= 16'hffe1; 
        10'b0001000010: data <= 16'h0008; 
        10'b0001000011: data <= 16'hffc5; 
        10'b0001000100: data <= 16'hfffd; 
        10'b0001000101: data <= 16'hffd6; 
        10'b0001000110: data <= 16'hffca; 
        10'b0001000111: data <= 16'hffd4; 
        10'b0001001000: data <= 16'hffdd; 
        10'b0001001001: data <= 16'hffeb; 
        10'b0001001010: data <= 16'hffe1; 
        10'b0001001011: data <= 16'hffe2; 
        10'b0001001100: data <= 16'h000e; 
        10'b0001001101: data <= 16'h0001; 
        10'b0001001110: data <= 16'h0006; 
        10'b0001001111: data <= 16'hffd5; 
        10'b0001010000: data <= 16'hffc8; 
        10'b0001010001: data <= 16'hffe4; 
        10'b0001010010: data <= 16'hfffd; 
        10'b0001010011: data <= 16'hfff1; 
        10'b0001010100: data <= 16'hfff6; 
        10'b0001010101: data <= 16'hfff0; 
        10'b0001010110: data <= 16'hffd3; 
        10'b0001010111: data <= 16'hfffd; 
        10'b0001011000: data <= 16'hffce; 
        10'b0001011001: data <= 16'hffdf; 
        10'b0001011010: data <= 16'hffc5; 
        10'b0001011011: data <= 16'hffd9; 
        10'b0001011100: data <= 16'hffc9; 
        10'b0001011101: data <= 16'hffd9; 
        10'b0001011110: data <= 16'hffa0; 
        10'b0001011111: data <= 16'hff86; 
        10'b0001100000: data <= 16'hffba; 
        10'b0001100001: data <= 16'hffbf; 
        10'b0001100010: data <= 16'hffb0; 
        10'b0001100011: data <= 16'hffe5; 
        10'b0001100100: data <= 16'hfff4; 
        10'b0001100101: data <= 16'hffc1; 
        10'b0001100110: data <= 16'hffda; 
        10'b0001100111: data <= 16'hfff4; 
        10'b0001101000: data <= 16'hfff7; 
        10'b0001101001: data <= 16'hffe6; 
        10'b0001101010: data <= 16'hffc0; 
        10'b0001101011: data <= 16'hffd5; 
        10'b0001101100: data <= 16'hffb3; 
        10'b0001101101: data <= 16'h0009; 
        10'b0001101110: data <= 16'h0006; 
        10'b0001101111: data <= 16'hffcd; 
        10'b0001110000: data <= 16'hffca; 
        10'b0001110001: data <= 16'hffdf; 
        10'b0001110010: data <= 16'h0005; 
        10'b0001110011: data <= 16'h0003; 
        10'b0001110100: data <= 16'h0007; 
        10'b0001110101: data <= 16'hffd9; 
        10'b0001110110: data <= 16'hffd6; 
        10'b0001110111: data <= 16'hffaa; 
        10'b0001111000: data <= 16'hff6e; 
        10'b0001111001: data <= 16'hff3e; 
        10'b0001111010: data <= 16'hfee5; 
        10'b0001111011: data <= 16'hff4b; 
        10'b0001111100: data <= 16'hff4a; 
        10'b0001111101: data <= 16'hff0c; 
        10'b0001111110: data <= 16'hff7a; 
        10'b0001111111: data <= 16'hffff; 
        10'b0010000000: data <= 16'hfff0; 
        10'b0010000001: data <= 16'h002e; 
        10'b0010000010: data <= 16'hfff2; 
        10'b0010000011: data <= 16'hffbb; 
        10'b0010000100: data <= 16'hffa5; 
        10'b0010000101: data <= 16'hffd0; 
        10'b0010000110: data <= 16'hffd9; 
        10'b0010000111: data <= 16'hffe4; 
        10'b0010001000: data <= 16'hffde; 
        10'b0010001001: data <= 16'h000d; 
        10'b0010001010: data <= 16'h0007; 
        10'b0010001011: data <= 16'hffe7; 
        10'b0010001100: data <= 16'hffeb; 
        10'b0010001101: data <= 16'h000d; 
        10'b0010001110: data <= 16'hffd4; 
        10'b0010001111: data <= 16'hffce; 
        10'b0010010000: data <= 16'hffdb; 
        10'b0010010001: data <= 16'hffa8; 
        10'b0010010010: data <= 16'hff7b; 
        10'b0010010011: data <= 16'hff7f; 
        10'b0010010100: data <= 16'hffac; 
        10'b0010010101: data <= 16'hfff0; 
        10'b0010010110: data <= 16'h001c; 
        10'b0010010111: data <= 16'h001f; 
        10'b0010011000: data <= 16'hffd2; 
        10'b0010011001: data <= 16'hffbf; 
        10'b0010011010: data <= 16'hffd9; 
        10'b0010011011: data <= 16'hffee; 
        10'b0010011100: data <= 16'h0041; 
        10'b0010011101: data <= 16'h0043; 
        10'b0010011110: data <= 16'h007f; 
        10'b0010011111: data <= 16'h004f; 
        10'b0010100000: data <= 16'h004d; 
        10'b0010100001: data <= 16'h0062; 
        10'b0010100010: data <= 16'h00b5; 
        10'b0010100011: data <= 16'h009a; 
        10'b0010100100: data <= 16'h006c; 
        10'b0010100101: data <= 16'h003c; 
        10'b0010100110: data <= 16'h0025; 
        10'b0010100111: data <= 16'h000e; 
        10'b0010101000: data <= 16'hffd0; 
        10'b0010101001: data <= 16'hffcb; 
        10'b0010101010: data <= 16'h0007; 
        10'b0010101011: data <= 16'hffcd; 
        10'b0010101100: data <= 16'hffbf; 
        10'b0010101101: data <= 16'hff64; 
        10'b0010101110: data <= 16'hffba; 
        10'b0010101111: data <= 16'hfff8; 
        10'b0010110000: data <= 16'hfffa; 
        10'b0010110001: data <= 16'h003f; 
        10'b0010110010: data <= 16'h0083; 
        10'b0010110011: data <= 16'h006d; 
        10'b0010110100: data <= 16'h0013; 
        10'b0010110101: data <= 16'h0028; 
        10'b0010110110: data <= 16'hffee; 
        10'b0010110111: data <= 16'hffc2; 
        10'b0010111000: data <= 16'hffda; 
        10'b0010111001: data <= 16'hffe0; 
        10'b0010111010: data <= 16'h0001; 
        10'b0010111011: data <= 16'h007c; 
        10'b0010111100: data <= 16'h0047; 
        10'b0010111101: data <= 16'h0051; 
        10'b0010111110: data <= 16'h00f7; 
        10'b0010111111: data <= 16'h0129; 
        10'b0011000000: data <= 16'h014f; 
        10'b0011000001: data <= 16'h00b1; 
        10'b0011000010: data <= 16'h0057; 
        10'b0011000011: data <= 16'h0015; 
        10'b0011000100: data <= 16'hffe5; 
        10'b0011000101: data <= 16'hfff1; 
        10'b0011000110: data <= 16'hffeb; 
        10'b0011000111: data <= 16'hffc0; 
        10'b0011001000: data <= 16'hff4b; 
        10'b0011001001: data <= 16'hff2c; 
        10'b0011001010: data <= 16'hff7f; 
        10'b0011001011: data <= 16'h0011; 
        10'b0011001100: data <= 16'h0055; 
        10'b0011001101: data <= 16'h00a6; 
        10'b0011001110: data <= 16'h00a2; 
        10'b0011001111: data <= 16'h008d; 
        10'b0011010000: data <= 16'h0029; 
        10'b0011010001: data <= 16'hfff3; 
        10'b0011010010: data <= 16'hffd3; 
        10'b0011010011: data <= 16'h0003; 
        10'b0011010100: data <= 16'h0046; 
        10'b0011010101: data <= 16'h003f; 
        10'b0011010110: data <= 16'h0050; 
        10'b0011010111: data <= 16'h00b3; 
        10'b0011011000: data <= 16'h009b; 
        10'b0011011001: data <= 16'h00b9; 
        10'b0011011010: data <= 16'h0103; 
        10'b0011011011: data <= 16'h015b; 
        10'b0011011100: data <= 16'h01a8; 
        10'b0011011101: data <= 16'h0132; 
        10'b0011011110: data <= 16'h002f; 
        10'b0011011111: data <= 16'hfff9; 
        10'b0011100000: data <= 16'hfff4; 
        10'b0011100001: data <= 16'h000b; 
        10'b0011100010: data <= 16'hffff; 
        10'b0011100011: data <= 16'hffa9; 
        10'b0011100100: data <= 16'hfefb; 
        10'b0011100101: data <= 16'hff21; 
        10'b0011100110: data <= 16'hff5f; 
        10'b0011100111: data <= 16'h000a; 
        10'b0011101000: data <= 16'h007e; 
        10'b0011101001: data <= 16'h0025; 
        10'b0011101010: data <= 16'h0044; 
        10'b0011101011: data <= 16'h0083; 
        10'b0011101100: data <= 16'h0050; 
        10'b0011101101: data <= 16'hffa6; 
        10'b0011101110: data <= 16'hff3a; 
        10'b0011101111: data <= 16'hff88; 
        10'b0011110000: data <= 16'hffb7; 
        10'b0011110001: data <= 16'h0007; 
        10'b0011110010: data <= 16'h0014; 
        10'b0011110011: data <= 16'h0095; 
        10'b0011110100: data <= 16'h009e; 
        10'b0011110101: data <= 16'h00e1; 
        10'b0011110110: data <= 16'h0163; 
        10'b0011110111: data <= 16'h01d0; 
        10'b0011111000: data <= 16'h026c; 
        10'b0011111001: data <= 16'h0190; 
        10'b0011111010: data <= 16'h0049; 
        10'b0011111011: data <= 16'hfff9; 
        10'b0011111100: data <= 16'hffcd; 
        10'b0011111101: data <= 16'hffe2; 
        10'b0011111110: data <= 16'hffc8; 
        10'b0011111111: data <= 16'hff86; 
        10'b0100000000: data <= 16'hff74; 
        10'b0100000001: data <= 16'hff7f; 
        10'b0100000010: data <= 16'h0010; 
        10'b0100000011: data <= 16'hfff7; 
        10'b0100000100: data <= 16'h006c; 
        10'b0100000101: data <= 16'h005d; 
        10'b0100000110: data <= 16'h0066; 
        10'b0100000111: data <= 16'h010f; 
        10'b0100001000: data <= 16'h00af; 
        10'b0100001001: data <= 16'hffb7; 
        10'b0100001010: data <= 16'hff12; 
        10'b0100001011: data <= 16'hfeaa; 
        10'b0100001100: data <= 16'hfec1; 
        10'b0100001101: data <= 16'hff46; 
        10'b0100001110: data <= 16'hffd5; 
        10'b0100001111: data <= 16'hffff; 
        10'b0100010000: data <= 16'h0091; 
        10'b0100010001: data <= 16'h0136; 
        10'b0100010010: data <= 16'h01c1; 
        10'b0100010011: data <= 16'h0266; 
        10'b0100010100: data <= 16'h0304; 
        10'b0100010101: data <= 16'h01fb; 
        10'b0100010110: data <= 16'h005b; 
        10'b0100010111: data <= 16'hffdc; 
        10'b0100011000: data <= 16'hfff5; 
        10'b0100011001: data <= 16'hffdd; 
        10'b0100011010: data <= 16'hffd0; 
        10'b0100011011: data <= 16'hffd9; 
        10'b0100011100: data <= 16'hffd7; 
        10'b0100011101: data <= 16'hffe6; 
        10'b0100011110: data <= 16'h0057; 
        10'b0100011111: data <= 16'h00a1; 
        10'b0100100000: data <= 16'h00fc; 
        10'b0100100001: data <= 16'h0117; 
        10'b0100100010: data <= 16'h010a; 
        10'b0100100011: data <= 16'h0142; 
        10'b0100100100: data <= 16'h010c; 
        10'b0100100101: data <= 16'h00ce; 
        10'b0100100110: data <= 16'hffd4; 
        10'b0100100111: data <= 16'hff58; 
        10'b0100101000: data <= 16'hfee7; 
        10'b0100101001: data <= 16'hfef0; 
        10'b0100101010: data <= 16'hfee6; 
        10'b0100101011: data <= 16'hfebf; 
        10'b0100101100: data <= 16'hff24; 
        10'b0100101101: data <= 16'hffbc; 
        10'b0100101110: data <= 16'h0025; 
        10'b0100101111: data <= 16'h00ce; 
        10'b0100110000: data <= 16'h019b; 
        10'b0100110001: data <= 16'h0135; 
        10'b0100110010: data <= 16'h0069; 
        10'b0100110011: data <= 16'hffdc; 
        10'b0100110100: data <= 16'hffd0; 
        10'b0100110101: data <= 16'h0000; 
        10'b0100110110: data <= 16'hffd9; 
        10'b0100110111: data <= 16'hffe6; 
        10'b0100111000: data <= 16'hffd8; 
        10'b0100111001: data <= 16'hfffa; 
        10'b0100111010: data <= 16'h008a; 
        10'b0100111011: data <= 16'h00a8; 
        10'b0100111100: data <= 16'h00f3; 
        10'b0100111101: data <= 16'h00e0; 
        10'b0100111110: data <= 16'h00a4; 
        10'b0100111111: data <= 16'h00b5; 
        10'b0101000000: data <= 16'h012b; 
        10'b0101000001: data <= 16'h0118; 
        10'b0101000010: data <= 16'h0004; 
        10'b0101000011: data <= 16'hff52; 
        10'b0101000100: data <= 16'hff28; 
        10'b0101000101: data <= 16'hff17; 
        10'b0101000110: data <= 16'hfeca; 
        10'b0101000111: data <= 16'hfe4f; 
        10'b0101001000: data <= 16'hfd8b; 
        10'b0101001001: data <= 16'hfdbf; 
        10'b0101001010: data <= 16'hfe27; 
        10'b0101001011: data <= 16'hfea7; 
        10'b0101001100: data <= 16'hff85; 
        10'b0101001101: data <= 16'h000d; 
        10'b0101001110: data <= 16'h0023; 
        10'b0101001111: data <= 16'hffeb; 
        10'b0101010000: data <= 16'hffea; 
        10'b0101010001: data <= 16'hffee; 
        10'b0101010010: data <= 16'hffe6; 
        10'b0101010011: data <= 16'hffdc; 
        10'b0101010100: data <= 16'hffe5; 
        10'b0101010101: data <= 16'h0046; 
        10'b0101010110: data <= 16'h009e; 
        10'b0101010111: data <= 16'h008d; 
        10'b0101011000: data <= 16'h0068; 
        10'b0101011001: data <= 16'h003b; 
        10'b0101011010: data <= 16'h00af; 
        10'b0101011011: data <= 16'h016a; 
        10'b0101011100: data <= 16'h0152; 
        10'b0101011101: data <= 16'h015b; 
        10'b0101011110: data <= 16'h0024; 
        10'b0101011111: data <= 16'hff50; 
        10'b0101100000: data <= 16'hfeb9; 
        10'b0101100001: data <= 16'hfef7; 
        10'b0101100010: data <= 16'hff4c; 
        10'b0101100011: data <= 16'hfefe; 
        10'b0101100100: data <= 16'hfeda; 
        10'b0101100101: data <= 16'hfe18; 
        10'b0101100110: data <= 16'hfdd3; 
        10'b0101100111: data <= 16'hfe1c; 
        10'b0101101000: data <= 16'hfebd; 
        10'b0101101001: data <= 16'hffa4; 
        10'b0101101010: data <= 16'h0005; 
        10'b0101101011: data <= 16'h0000; 
        10'b0101101100: data <= 16'hffed; 
        10'b0101101101: data <= 16'hffd2; 
        10'b0101101110: data <= 16'hffcf; 
        10'b0101101111: data <= 16'hffde; 
        10'b0101110000: data <= 16'hfff6; 
        10'b0101110001: data <= 16'h0024; 
        10'b0101110010: data <= 16'h006a; 
        10'b0101110011: data <= 16'h004e; 
        10'b0101110100: data <= 16'h005a; 
        10'b0101110101: data <= 16'h004a; 
        10'b0101110110: data <= 16'h00f4; 
        10'b0101110111: data <= 16'h0110; 
        10'b0101111000: data <= 16'h00cb; 
        10'b0101111001: data <= 16'h00bd; 
        10'b0101111010: data <= 16'hffda; 
        10'b0101111011: data <= 16'hff2f; 
        10'b0101111100: data <= 16'hfeab; 
        10'b0101111101: data <= 16'hff4c; 
        10'b0101111110: data <= 16'hffc0; 
        10'b0101111111: data <= 16'hffb6; 
        10'b0110000000: data <= 16'hffdd; 
        10'b0110000001: data <= 16'hff76; 
        10'b0110000010: data <= 16'hff06; 
        10'b0110000011: data <= 16'hfe93; 
        10'b0110000100: data <= 16'hfeed; 
        10'b0110000101: data <= 16'hffd0; 
        10'b0110000110: data <= 16'hffcc; 
        10'b0110000111: data <= 16'hfff8; 
        10'b0110001000: data <= 16'hffee; 
        10'b0110001001: data <= 16'hffce; 
        10'b0110001010: data <= 16'hffe8; 
        10'b0110001011: data <= 16'hffc3; 
        10'b0110001100: data <= 16'hffeb; 
        10'b0110001101: data <= 16'hffea; 
        10'b0110001110: data <= 16'hffff; 
        10'b0110001111: data <= 16'hfff4; 
        10'b0110010000: data <= 16'h0070; 
        10'b0110010001: data <= 16'h00b1; 
        10'b0110010010: data <= 16'h00d5; 
        10'b0110010011: data <= 16'h0029; 
        10'b0110010100: data <= 16'h0048; 
        10'b0110010101: data <= 16'hfff3; 
        10'b0110010110: data <= 16'hff68; 
        10'b0110010111: data <= 16'hff51; 
        10'b0110011000: data <= 16'hff0d; 
        10'b0110011001: data <= 16'hff29; 
        10'b0110011010: data <= 16'hff37; 
        10'b0110011011: data <= 16'hff9f; 
        10'b0110011100: data <= 16'hffac; 
        10'b0110011101: data <= 16'hffb4; 
        10'b0110011110: data <= 16'hffd2; 
        10'b0110011111: data <= 16'hff37; 
        10'b0110100000: data <= 16'hff79; 
        10'b0110100001: data <= 16'hffbc; 
        10'b0110100010: data <= 16'hffe8; 
        10'b0110100011: data <= 16'hffc4; 
        10'b0110100100: data <= 16'hffca; 
        10'b0110100101: data <= 16'h0008; 
        10'b0110100110: data <= 16'hffc6; 
        10'b0110100111: data <= 16'hffe8; 
        10'b0110101000: data <= 16'hffaa; 
        10'b0110101001: data <= 16'hff7f; 
        10'b0110101010: data <= 16'hff4c; 
        10'b0110101011: data <= 16'hff89; 
        10'b0110101100: data <= 16'h002b; 
        10'b0110101101: data <= 16'h00c8; 
        10'b0110101110: data <= 16'h005f; 
        10'b0110101111: data <= 16'h0057; 
        10'b0110110000: data <= 16'h004b; 
        10'b0110110001: data <= 16'hffbc; 
        10'b0110110010: data <= 16'hff1e; 
        10'b0110110011: data <= 16'hfefc; 
        10'b0110110100: data <= 16'hff16; 
        10'b0110110101: data <= 16'hff10; 
        10'b0110110110: data <= 16'hff57; 
        10'b0110110111: data <= 16'hfff7; 
        10'b0110111000: data <= 16'hffc7; 
        10'b0110111001: data <= 16'hffd0; 
        10'b0110111010: data <= 16'hffc6; 
        10'b0110111011: data <= 16'hffbd; 
        10'b0110111100: data <= 16'hffd1; 
        10'b0110111101: data <= 16'hffff; 
        10'b0110111110: data <= 16'h0009; 
        10'b0110111111: data <= 16'hffdc; 
        10'b0111000000: data <= 16'hffe0; 
        10'b0111000001: data <= 16'hffeb; 
        10'b0111000010: data <= 16'hfff2; 
        10'b0111000011: data <= 16'hffc6; 
        10'b0111000100: data <= 16'hffde; 
        10'b0111000101: data <= 16'hff6d; 
        10'b0111000110: data <= 16'hfeda; 
        10'b0111000111: data <= 16'hfea5; 
        10'b0111001000: data <= 16'hff15; 
        10'b0111001001: data <= 16'hff7e; 
        10'b0111001010: data <= 16'hffcc; 
        10'b0111001011: data <= 16'hffb6; 
        10'b0111001100: data <= 16'hffd0; 
        10'b0111001101: data <= 16'hff60; 
        10'b0111001110: data <= 16'hfecc; 
        10'b0111001111: data <= 16'hff06; 
        10'b0111010000: data <= 16'hff4a; 
        10'b0111010001: data <= 16'hffbe; 
        10'b0111010010: data <= 16'hffc2; 
        10'b0111010011: data <= 16'h000a; 
        10'b0111010100: data <= 16'h0033; 
        10'b0111010101: data <= 16'h0008; 
        10'b0111010110: data <= 16'h0037; 
        10'b0111010111: data <= 16'h000d; 
        10'b0111011000: data <= 16'h0009; 
        10'b0111011001: data <= 16'h0008; 
        10'b0111011010: data <= 16'hffdd; 
        10'b0111011011: data <= 16'hffe0; 
        10'b0111011100: data <= 16'hffda; 
        10'b0111011101: data <= 16'hfffd; 
        10'b0111011110: data <= 16'h0000; 
        10'b0111011111: data <= 16'h0004; 
        10'b0111100000: data <= 16'hffdb; 
        10'b0111100001: data <= 16'h000b; 
        10'b0111100010: data <= 16'h0015; 
        10'b0111100011: data <= 16'hff1b; 
        10'b0111100100: data <= 16'hfe61; 
        10'b0111100101: data <= 16'hfe7c; 
        10'b0111100110: data <= 16'hfeea; 
        10'b0111100111: data <= 16'hff59; 
        10'b0111101000: data <= 16'hfefa; 
        10'b0111101001: data <= 16'hfeae; 
        10'b0111101010: data <= 16'hfeb8; 
        10'b0111101011: data <= 16'hff6b; 
        10'b0111101100: data <= 16'hffbe; 
        10'b0111101101: data <= 16'h0063; 
        10'b0111101110: data <= 16'h0098; 
        10'b0111101111: data <= 16'h0063; 
        10'b0111110000: data <= 16'h0064; 
        10'b0111110001: data <= 16'h001d; 
        10'b0111110010: data <= 16'h0003; 
        10'b0111110011: data <= 16'h0037; 
        10'b0111110100: data <= 16'h0038; 
        10'b0111110101: data <= 16'hffd1; 
        10'b0111110110: data <= 16'hfffe; 
        10'b0111110111: data <= 16'h0001; 
        10'b0111111000: data <= 16'h0006; 
        10'b0111111001: data <= 16'hffd8; 
        10'b0111111010: data <= 16'hffe7; 
        10'b0111111011: data <= 16'hffdf; 
        10'b0111111100: data <= 16'h0052; 
        10'b0111111101: data <= 16'h006c; 
        10'b0111111110: data <= 16'h0102; 
        10'b0111111111: data <= 16'h002d; 
        10'b1000000000: data <= 16'hff08; 
        10'b1000000001: data <= 16'hfe97; 
        10'b1000000010: data <= 16'hfe25; 
        10'b1000000011: data <= 16'hfe58; 
        10'b1000000100: data <= 16'hfed0; 
        10'b1000000101: data <= 16'hff52; 
        10'b1000000110: data <= 16'hffa9; 
        10'b1000000111: data <= 16'hffdc; 
        10'b1000001000: data <= 16'hfff9; 
        10'b1000001001: data <= 16'h0074; 
        10'b1000001010: data <= 16'h003b; 
        10'b1000001011: data <= 16'h0068; 
        10'b1000001100: data <= 16'h0046; 
        10'b1000001101: data <= 16'h0065; 
        10'b1000001110: data <= 16'h0053; 
        10'b1000001111: data <= 16'h0073; 
        10'b1000010000: data <= 16'h003c; 
        10'b1000010001: data <= 16'h0004; 
        10'b1000010010: data <= 16'hffd4; 
        10'b1000010011: data <= 16'hfff2; 
        10'b1000010100: data <= 16'h0000; 
        10'b1000010101: data <= 16'hffd7; 
        10'b1000010110: data <= 16'hffea; 
        10'b1000010111: data <= 16'h0009; 
        10'b1000011000: data <= 16'h007d; 
        10'b1000011001: data <= 16'h00d5; 
        10'b1000011010: data <= 16'h011f; 
        10'b1000011011: data <= 16'h00c1; 
        10'b1000011100: data <= 16'h007a; 
        10'b1000011101: data <= 16'h0028; 
        10'b1000011110: data <= 16'hffa5; 
        10'b1000011111: data <= 16'hff9f; 
        10'b1000100000: data <= 16'h0008; 
        10'b1000100001: data <= 16'h0075; 
        10'b1000100010: data <= 16'h002c; 
        10'b1000100011: data <= 16'h003e; 
        10'b1000100100: data <= 16'h003f; 
        10'b1000100101: data <= 16'hffec; 
        10'b1000100110: data <= 16'h002d; 
        10'b1000100111: data <= 16'h002c; 
        10'b1000101000: data <= 16'h0009; 
        10'b1000101001: data <= 16'h004c; 
        10'b1000101010: data <= 16'h0082; 
        10'b1000101011: data <= 16'h005f; 
        10'b1000101100: data <= 16'h0008; 
        10'b1000101101: data <= 16'hfffe; 
        10'b1000101110: data <= 16'h0000; 
        10'b1000101111: data <= 16'hffcd; 
        10'b1000110000: data <= 16'hfffd; 
        10'b1000110001: data <= 16'hffc4; 
        10'b1000110010: data <= 16'hffe4; 
        10'b1000110011: data <= 16'hffd4; 
        10'b1000110100: data <= 16'h0011; 
        10'b1000110101: data <= 16'h008c; 
        10'b1000110110: data <= 16'h00a3; 
        10'b1000110111: data <= 16'h00c6; 
        10'b1000111000: data <= 16'h0116; 
        10'b1000111001: data <= 16'h00ea; 
        10'b1000111010: data <= 16'h00ce; 
        10'b1000111011: data <= 16'h012c; 
        10'b1000111100: data <= 16'h00bb; 
        10'b1000111101: data <= 16'h008c; 
        10'b1000111110: data <= 16'hffd9; 
        10'b1000111111: data <= 16'hffdc; 
        10'b1001000000: data <= 16'h0067; 
        10'b1001000001: data <= 16'h0035; 
        10'b1001000010: data <= 16'h0056; 
        10'b1001000011: data <= 16'h0072; 
        10'b1001000100: data <= 16'h0064; 
        10'b1001000101: data <= 16'h004f; 
        10'b1001000110: data <= 16'h00bc; 
        10'b1001000111: data <= 16'h008c; 
        10'b1001001000: data <= 16'hffee; 
        10'b1001001001: data <= 16'hffc6; 
        10'b1001001010: data <= 16'hffeb; 
        10'b1001001011: data <= 16'hffdb; 
        10'b1001001100: data <= 16'hffd6; 
        10'b1001001101: data <= 16'h0001; 
        10'b1001001110: data <= 16'hffc2; 
        10'b1001001111: data <= 16'hffe9; 
        10'b1001010000: data <= 16'h0037; 
        10'b1001010001: data <= 16'hffee; 
        10'b1001010010: data <= 16'h0043; 
        10'b1001010011: data <= 16'h00b5; 
        10'b1001010100: data <= 16'h0106; 
        10'b1001010101: data <= 16'h00ab; 
        10'b1001010110: data <= 16'h0091; 
        10'b1001010111: data <= 16'h004e; 
        10'b1001011000: data <= 16'h0065; 
        10'b1001011001: data <= 16'h003f; 
        10'b1001011010: data <= 16'h0041; 
        10'b1001011011: data <= 16'h0050; 
        10'b1001011100: data <= 16'h0015; 
        10'b1001011101: data <= 16'h0040; 
        10'b1001011110: data <= 16'h0021; 
        10'b1001011111: data <= 16'h0068; 
        10'b1001100000: data <= 16'h0066; 
        10'b1001100001: data <= 16'h00ab; 
        10'b1001100010: data <= 16'h00d2; 
        10'b1001100011: data <= 16'h002d; 
        10'b1001100100: data <= 16'h0002; 
        10'b1001100101: data <= 16'hffce; 
        10'b1001100110: data <= 16'hffdc; 
        10'b1001100111: data <= 16'hffdc; 
        10'b1001101000: data <= 16'hfff4; 
        10'b1001101001: data <= 16'hffc7; 
        10'b1001101010: data <= 16'hffe3; 
        10'b1001101011: data <= 16'hffdc; 
        10'b1001101100: data <= 16'h0014; 
        10'b1001101101: data <= 16'hffe4; 
        10'b1001101110: data <= 16'hffc3; 
        10'b1001101111: data <= 16'hfff5; 
        10'b1001110000: data <= 16'h0066; 
        10'b1001110001: data <= 16'h0095; 
        10'b1001110010: data <= 16'h001a; 
        10'b1001110011: data <= 16'h0084; 
        10'b1001110100: data <= 16'h00d5; 
        10'b1001110101: data <= 16'h0107; 
        10'b1001110110: data <= 16'h0086; 
        10'b1001110111: data <= 16'h0014; 
        10'b1001111000: data <= 16'h000f; 
        10'b1001111001: data <= 16'h0021; 
        10'b1001111010: data <= 16'h0045; 
        10'b1001111011: data <= 16'h0044; 
        10'b1001111100: data <= 16'h0075; 
        10'b1001111101: data <= 16'h006a; 
        10'b1001111110: data <= 16'h006f; 
        10'b1001111111: data <= 16'h0027; 
        10'b1010000000: data <= 16'hfffa; 
        10'b1010000001: data <= 16'h0006; 
        10'b1010000010: data <= 16'hffeb; 
        10'b1010000011: data <= 16'hfff2; 
        10'b1010000100: data <= 16'hffd1; 
        10'b1010000101: data <= 16'hffe9; 
        10'b1010000110: data <= 16'hfff3; 
        10'b1010000111: data <= 16'hffee; 
        10'b1010001000: data <= 16'hffd4; 
        10'b1010001001: data <= 16'hffe3; 
        10'b1010001010: data <= 16'hffa7; 
        10'b1010001011: data <= 16'hffd8; 
        10'b1010001100: data <= 16'h0051; 
        10'b1010001101: data <= 16'h004f; 
        10'b1010001110: data <= 16'h004f; 
        10'b1010001111: data <= 16'h008c; 
        10'b1010010000: data <= 16'h0087; 
        10'b1010010001: data <= 16'h005c; 
        10'b1010010010: data <= 16'h006a; 
        10'b1010010011: data <= 16'h0061; 
        10'b1010010100: data <= 16'h005f; 
        10'b1010010101: data <= 16'h002c; 
        10'b1010010110: data <= 16'hffce; 
        10'b1010010111: data <= 16'hfff9; 
        10'b1010011000: data <= 16'h002f; 
        10'b1010011001: data <= 16'h0013; 
        10'b1010011010: data <= 16'h003e; 
        10'b1010011011: data <= 16'hffd9; 
        10'b1010011100: data <= 16'h000a; 
        10'b1010011101: data <= 16'hffe0; 
        10'b1010011110: data <= 16'hffdf; 
        10'b1010011111: data <= 16'h000a; 
        10'b1010100000: data <= 16'hfffc; 
        10'b1010100001: data <= 16'hffe1; 
        10'b1010100010: data <= 16'hffdd; 
        10'b1010100011: data <= 16'h000b; 
        10'b1010100100: data <= 16'hffc3; 
        10'b1010100101: data <= 16'hffbf; 
        10'b1010100110: data <= 16'hffe9; 
        10'b1010100111: data <= 16'hfff4; 
        10'b1010101000: data <= 16'hfffc; 
        10'b1010101001: data <= 16'h0068; 
        10'b1010101010: data <= 16'h0087; 
        10'b1010101011: data <= 16'h0068; 
        10'b1010101100: data <= 16'h0044; 
        10'b1010101101: data <= 16'h005e; 
        10'b1010101110: data <= 16'h00ae; 
        10'b1010101111: data <= 16'h0090; 
        10'b1010110000: data <= 16'h0056; 
        10'b1010110001: data <= 16'h002a; 
        10'b1010110010: data <= 16'h004f; 
        10'b1010110011: data <= 16'h0034; 
        10'b1010110100: data <= 16'hfffd; 
        10'b1010110101: data <= 16'hfff9; 
        10'b1010110110: data <= 16'hffed; 
        10'b1010110111: data <= 16'h0003; 
        10'b1010111000: data <= 16'hffd6; 
        10'b1010111001: data <= 16'hfff1; 
        10'b1010111010: data <= 16'h0006; 
        10'b1010111011: data <= 16'hffcd; 
        10'b1010111100: data <= 16'hffe9; 
        10'b1010111101: data <= 16'h0002; 
        10'b1010111110: data <= 16'h0006; 
        10'b1010111111: data <= 16'hffca; 
        10'b1011000000: data <= 16'h0000; 
        10'b1011000001: data <= 16'hffef; 
        10'b1011000010: data <= 16'hffc0; 
        10'b1011000011: data <= 16'hffe8; 
        10'b1011000100: data <= 16'hffc7; 
        10'b1011000101: data <= 16'h0022; 
        10'b1011000110: data <= 16'h0019; 
        10'b1011000111: data <= 16'h0046; 
        10'b1011001000: data <= 16'h0046; 
        10'b1011001001: data <= 16'h007b; 
        10'b1011001010: data <= 16'h0007; 
        10'b1011001011: data <= 16'h0025; 
        10'b1011001100: data <= 16'h001f; 
        10'b1011001101: data <= 16'h003c; 
        10'b1011001110: data <= 16'hffd8; 
        10'b1011001111: data <= 16'hfffe; 
        10'b1011010000: data <= 16'hffbd; 
        10'b1011010001: data <= 16'h0006; 
        10'b1011010010: data <= 16'hffe7; 
        10'b1011010011: data <= 16'hffd3; 
        10'b1011010100: data <= 16'hfffb; 
        10'b1011010101: data <= 16'h0003; 
        10'b1011010110: data <= 16'hffc7; 
        10'b1011010111: data <= 16'hffe2; 
        10'b1011011000: data <= 16'hffee; 
        10'b1011011001: data <= 16'hffec; 
        10'b1011011010: data <= 16'hffd6; 
        10'b1011011011: data <= 16'hffe0; 
        10'b1011011100: data <= 16'hffdd; 
        10'b1011011101: data <= 16'hffe3; 
        10'b1011011110: data <= 16'hfff6; 
        10'b1011011111: data <= 16'hffd6; 
        10'b1011100000: data <= 16'hffc9; 
        10'b1011100001: data <= 16'hffe3; 
        10'b1011100010: data <= 16'hffda; 
        10'b1011100011: data <= 16'hfff9; 
        10'b1011100100: data <= 16'h0001; 
        10'b1011100101: data <= 16'hfff2; 
        10'b1011100110: data <= 16'hffd8; 
        10'b1011100111: data <= 16'hffec; 
        10'b1011101000: data <= 16'hfff7; 
        10'b1011101001: data <= 16'hffd6; 
        10'b1011101010: data <= 16'hffaf; 
        10'b1011101011: data <= 16'hffbf; 
        10'b1011101100: data <= 16'hfff2; 
        10'b1011101101: data <= 16'hfff2; 
        10'b1011101110: data <= 16'hffdb; 
        10'b1011101111: data <= 16'hfff5; 
        10'b1011110000: data <= 16'hffe4; 
        10'b1011110001: data <= 16'hffed; 
        10'b1011110010: data <= 16'hffde; 
        10'b1011110011: data <= 16'hffc7; 
        10'b1011110100: data <= 16'hfff3; 
        10'b1011110101: data <= 16'hfff8; 
        10'b1011110110: data <= 16'hfffb; 
        10'b1011110111: data <= 16'hfff0; 
        10'b1011111000: data <= 16'hffcf; 
        10'b1011111001: data <= 16'hfffd; 
        10'b1011111010: data <= 16'hffdf; 
        10'b1011111011: data <= 16'hffdc; 
        10'b1011111100: data <= 16'h000c; 
        10'b1011111101: data <= 16'hffde; 
        10'b1011111110: data <= 16'hffd9; 
        10'b1011111111: data <= 16'hfffb; 
        10'b1100000000: data <= 16'hffeb; 
        10'b1100000001: data <= 16'hffc4; 
        10'b1100000010: data <= 16'h0001; 
        10'b1100000011: data <= 16'hffee; 
        10'b1100000100: data <= 16'hffca; 
        10'b1100000101: data <= 16'hffc4; 
        10'b1100000110: data <= 16'hffd3; 
        10'b1100000111: data <= 16'hffc3; 
        10'b1100001000: data <= 16'hffff; 
        10'b1100001001: data <= 16'hffde; 
        10'b1100001010: data <= 16'h000b; 
        10'b1100001011: data <= 16'hffcc; 
        10'b1100001100: data <= 16'hfff0; 
        10'b1100001101: data <= 16'hffe6; 
        10'b1100001110: data <= 16'hffd0; 
        10'b1100001111: data <= 16'hfff8; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 11) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 17'h1ffb9; 
        10'b0000000001: data <= 17'h1fff6; 
        10'b0000000010: data <= 17'h1fff6; 
        10'b0000000011: data <= 17'h1ffa1; 
        10'b0000000100: data <= 17'h1ffd3; 
        10'b0000000101: data <= 17'h1ffc7; 
        10'b0000000110: data <= 17'h00000; 
        10'b0000000111: data <= 17'h1ffc3; 
        10'b0000001000: data <= 17'h1ffe7; 
        10'b0000001001: data <= 17'h00015; 
        10'b0000001010: data <= 17'h1ffe7; 
        10'b0000001011: data <= 17'h1ffe4; 
        10'b0000001100: data <= 17'h1ffb7; 
        10'b0000001101: data <= 17'h1fffc; 
        10'b0000001110: data <= 17'h1ff9f; 
        10'b0000001111: data <= 17'h1ffb0; 
        10'b0000010000: data <= 17'h1ff92; 
        10'b0000010001: data <= 17'h1ffa7; 
        10'b0000010010: data <= 17'h1fff3; 
        10'b0000010011: data <= 17'h1ffe7; 
        10'b0000010100: data <= 17'h1ff91; 
        10'b0000010101: data <= 17'h1ffd6; 
        10'b0000010110: data <= 17'h1ffe1; 
        10'b0000010111: data <= 17'h1ffc9; 
        10'b0000011000: data <= 17'h1ff97; 
        10'b0000011001: data <= 17'h1ffd8; 
        10'b0000011010: data <= 17'h1ffe1; 
        10'b0000011011: data <= 17'h1ffbc; 
        10'b0000011100: data <= 17'h1fff9; 
        10'b0000011101: data <= 17'h1ff8b; 
        10'b0000011110: data <= 17'h1ffff; 
        10'b0000011111: data <= 17'h1ff9c; 
        10'b0000100000: data <= 17'h1fffc; 
        10'b0000100001: data <= 17'h1ffc0; 
        10'b0000100010: data <= 17'h1ffdf; 
        10'b0000100011: data <= 17'h1ffbd; 
        10'b0000100100: data <= 17'h1ffac; 
        10'b0000100101: data <= 17'h1ffe1; 
        10'b0000100110: data <= 17'h0000a; 
        10'b0000100111: data <= 17'h1ff9f; 
        10'b0000101000: data <= 17'h1ffbc; 
        10'b0000101001: data <= 17'h1ffa9; 
        10'b0000101010: data <= 17'h1ff90; 
        10'b0000101011: data <= 17'h1ffed; 
        10'b0000101100: data <= 17'h1ffb4; 
        10'b0000101101: data <= 17'h1ffa7; 
        10'b0000101110: data <= 17'h1ffb6; 
        10'b0000101111: data <= 17'h1ffb1; 
        10'b0000110000: data <= 17'h1ffe7; 
        10'b0000110001: data <= 17'h1ff9a; 
        10'b0000110010: data <= 17'h1fffe; 
        10'b0000110011: data <= 17'h1ffa1; 
        10'b0000110100: data <= 17'h00001; 
        10'b0000110101: data <= 17'h1fff8; 
        10'b0000110110: data <= 17'h1ffa5; 
        10'b0000110111: data <= 17'h1ffce; 
        10'b0000111000: data <= 17'h1ffcf; 
        10'b0000111001: data <= 17'h1ffea; 
        10'b0000111010: data <= 17'h1ffbd; 
        10'b0000111011: data <= 17'h1ff91; 
        10'b0000111100: data <= 17'h1ffa4; 
        10'b0000111101: data <= 17'h1ffd9; 
        10'b0000111110: data <= 17'h1fffc; 
        10'b0000111111: data <= 17'h1ffe2; 
        10'b0001000000: data <= 17'h1ffaf; 
        10'b0001000001: data <= 17'h1ffc2; 
        10'b0001000010: data <= 17'h0000f; 
        10'b0001000011: data <= 17'h1ff8a; 
        10'b0001000100: data <= 17'h1fffa; 
        10'b0001000101: data <= 17'h1ffad; 
        10'b0001000110: data <= 17'h1ff93; 
        10'b0001000111: data <= 17'h1ffa8; 
        10'b0001001000: data <= 17'h1ffb9; 
        10'b0001001001: data <= 17'h1ffd7; 
        10'b0001001010: data <= 17'h1ffc2; 
        10'b0001001011: data <= 17'h1ffc3; 
        10'b0001001100: data <= 17'h0001b; 
        10'b0001001101: data <= 17'h00003; 
        10'b0001001110: data <= 17'h0000b; 
        10'b0001001111: data <= 17'h1ffaa; 
        10'b0001010000: data <= 17'h1ff90; 
        10'b0001010001: data <= 17'h1ffc8; 
        10'b0001010010: data <= 17'h1fff9; 
        10'b0001010011: data <= 17'h1ffe2; 
        10'b0001010100: data <= 17'h1ffeb; 
        10'b0001010101: data <= 17'h1ffe0; 
        10'b0001010110: data <= 17'h1ffa6; 
        10'b0001010111: data <= 17'h1fffa; 
        10'b0001011000: data <= 17'h1ff9c; 
        10'b0001011001: data <= 17'h1ffbe; 
        10'b0001011010: data <= 17'h1ff8a; 
        10'b0001011011: data <= 17'h1ffb3; 
        10'b0001011100: data <= 17'h1ff92; 
        10'b0001011101: data <= 17'h1ffb1; 
        10'b0001011110: data <= 17'h1ff41; 
        10'b0001011111: data <= 17'h1ff0c; 
        10'b0001100000: data <= 17'h1ff74; 
        10'b0001100001: data <= 17'h1ff7d; 
        10'b0001100010: data <= 17'h1ff5f; 
        10'b0001100011: data <= 17'h1ffcb; 
        10'b0001100100: data <= 17'h1ffe9; 
        10'b0001100101: data <= 17'h1ff82; 
        10'b0001100110: data <= 17'h1ffb4; 
        10'b0001100111: data <= 17'h1ffe8; 
        10'b0001101000: data <= 17'h1ffef; 
        10'b0001101001: data <= 17'h1ffcb; 
        10'b0001101010: data <= 17'h1ff80; 
        10'b0001101011: data <= 17'h1ffaa; 
        10'b0001101100: data <= 17'h1ff65; 
        10'b0001101101: data <= 17'h00012; 
        10'b0001101110: data <= 17'h0000b; 
        10'b0001101111: data <= 17'h1ff9b; 
        10'b0001110000: data <= 17'h1ff94; 
        10'b0001110001: data <= 17'h1ffbd; 
        10'b0001110010: data <= 17'h0000b; 
        10'b0001110011: data <= 17'h00006; 
        10'b0001110100: data <= 17'h0000f; 
        10'b0001110101: data <= 17'h1ffb3; 
        10'b0001110110: data <= 17'h1ffad; 
        10'b0001110111: data <= 17'h1ff53; 
        10'b0001111000: data <= 17'h1fedc; 
        10'b0001111001: data <= 17'h1fe7d; 
        10'b0001111010: data <= 17'h1fdcb; 
        10'b0001111011: data <= 17'h1fe97; 
        10'b0001111100: data <= 17'h1fe94; 
        10'b0001111101: data <= 17'h1fe18; 
        10'b0001111110: data <= 17'h1fef3; 
        10'b0001111111: data <= 17'h1ffff; 
        10'b0010000000: data <= 17'h1ffe0; 
        10'b0010000001: data <= 17'h0005b; 
        10'b0010000010: data <= 17'h1ffe4; 
        10'b0010000011: data <= 17'h1ff75; 
        10'b0010000100: data <= 17'h1ff4b; 
        10'b0010000101: data <= 17'h1ffa0; 
        10'b0010000110: data <= 17'h1ffb1; 
        10'b0010000111: data <= 17'h1ffc9; 
        10'b0010001000: data <= 17'h1ffbc; 
        10'b0010001001: data <= 17'h00019; 
        10'b0010001010: data <= 17'h0000e; 
        10'b0010001011: data <= 17'h1ffce; 
        10'b0010001100: data <= 17'h1ffd7; 
        10'b0010001101: data <= 17'h00019; 
        10'b0010001110: data <= 17'h1ffa9; 
        10'b0010001111: data <= 17'h1ff9c; 
        10'b0010010000: data <= 17'h1ffb6; 
        10'b0010010001: data <= 17'h1ff4f; 
        10'b0010010010: data <= 17'h1fef5; 
        10'b0010010011: data <= 17'h1fefe; 
        10'b0010010100: data <= 17'h1ff57; 
        10'b0010010101: data <= 17'h1ffe0; 
        10'b0010010110: data <= 17'h00039; 
        10'b0010010111: data <= 17'h0003d; 
        10'b0010011000: data <= 17'h1ffa5; 
        10'b0010011001: data <= 17'h1ff7d; 
        10'b0010011010: data <= 17'h1ffb1; 
        10'b0010011011: data <= 17'h1ffdb; 
        10'b0010011100: data <= 17'h00083; 
        10'b0010011101: data <= 17'h00086; 
        10'b0010011110: data <= 17'h000fd; 
        10'b0010011111: data <= 17'h0009e; 
        10'b0010100000: data <= 17'h00099; 
        10'b0010100001: data <= 17'h000c4; 
        10'b0010100010: data <= 17'h0016a; 
        10'b0010100011: data <= 17'h00134; 
        10'b0010100100: data <= 17'h000d8; 
        10'b0010100101: data <= 17'h00078; 
        10'b0010100110: data <= 17'h0004a; 
        10'b0010100111: data <= 17'h0001c; 
        10'b0010101000: data <= 17'h1ffa0; 
        10'b0010101001: data <= 17'h1ff97; 
        10'b0010101010: data <= 17'h0000d; 
        10'b0010101011: data <= 17'h1ff9b; 
        10'b0010101100: data <= 17'h1ff7e; 
        10'b0010101101: data <= 17'h1fec9; 
        10'b0010101110: data <= 17'h1ff74; 
        10'b0010101111: data <= 17'h1fff0; 
        10'b0010110000: data <= 17'h1fff5; 
        10'b0010110001: data <= 17'h0007e; 
        10'b0010110010: data <= 17'h00106; 
        10'b0010110011: data <= 17'h000da; 
        10'b0010110100: data <= 17'h00025; 
        10'b0010110101: data <= 17'h00050; 
        10'b0010110110: data <= 17'h1ffdc; 
        10'b0010110111: data <= 17'h1ff84; 
        10'b0010111000: data <= 17'h1ffb5; 
        10'b0010111001: data <= 17'h1ffc1; 
        10'b0010111010: data <= 17'h00003; 
        10'b0010111011: data <= 17'h000f9; 
        10'b0010111100: data <= 17'h0008e; 
        10'b0010111101: data <= 17'h000a2; 
        10'b0010111110: data <= 17'h001ef; 
        10'b0010111111: data <= 17'h00253; 
        10'b0011000000: data <= 17'h0029d; 
        10'b0011000001: data <= 17'h00162; 
        10'b0011000010: data <= 17'h000af; 
        10'b0011000011: data <= 17'h0002b; 
        10'b0011000100: data <= 17'h1ffc9; 
        10'b0011000101: data <= 17'h1ffe2; 
        10'b0011000110: data <= 17'h1ffd5; 
        10'b0011000111: data <= 17'h1ff80; 
        10'b0011001000: data <= 17'h1fe96; 
        10'b0011001001: data <= 17'h1fe57; 
        10'b0011001010: data <= 17'h1fefd; 
        10'b0011001011: data <= 17'h00021; 
        10'b0011001100: data <= 17'h000a9; 
        10'b0011001101: data <= 17'h0014c; 
        10'b0011001110: data <= 17'h00144; 
        10'b0011001111: data <= 17'h0011b; 
        10'b0011010000: data <= 17'h00052; 
        10'b0011010001: data <= 17'h1ffe5; 
        10'b0011010010: data <= 17'h1ffa6; 
        10'b0011010011: data <= 17'h00006; 
        10'b0011010100: data <= 17'h0008c; 
        10'b0011010101: data <= 17'h0007f; 
        10'b0011010110: data <= 17'h000a0; 
        10'b0011010111: data <= 17'h00166; 
        10'b0011011000: data <= 17'h00136; 
        10'b0011011001: data <= 17'h00173; 
        10'b0011011010: data <= 17'h00206; 
        10'b0011011011: data <= 17'h002b7; 
        10'b0011011100: data <= 17'h00350; 
        10'b0011011101: data <= 17'h00265; 
        10'b0011011110: data <= 17'h0005e; 
        10'b0011011111: data <= 17'h1fff1; 
        10'b0011100000: data <= 17'h1ffe8; 
        10'b0011100001: data <= 17'h00016; 
        10'b0011100010: data <= 17'h1fffe; 
        10'b0011100011: data <= 17'h1ff51; 
        10'b0011100100: data <= 17'h1fdf7; 
        10'b0011100101: data <= 17'h1fe42; 
        10'b0011100110: data <= 17'h1febe; 
        10'b0011100111: data <= 17'h00014; 
        10'b0011101000: data <= 17'h000fc; 
        10'b0011101001: data <= 17'h0004a; 
        10'b0011101010: data <= 17'h00087; 
        10'b0011101011: data <= 17'h00107; 
        10'b0011101100: data <= 17'h000a0; 
        10'b0011101101: data <= 17'h1ff4c; 
        10'b0011101110: data <= 17'h1fe74; 
        10'b0011101111: data <= 17'h1ff10; 
        10'b0011110000: data <= 17'h1ff6d; 
        10'b0011110001: data <= 17'h0000e; 
        10'b0011110010: data <= 17'h00028; 
        10'b0011110011: data <= 17'h0012b; 
        10'b0011110100: data <= 17'h0013b; 
        10'b0011110101: data <= 17'h001c1; 
        10'b0011110110: data <= 17'h002c6; 
        10'b0011110111: data <= 17'h003a1; 
        10'b0011111000: data <= 17'h004d7; 
        10'b0011111001: data <= 17'h00321; 
        10'b0011111010: data <= 17'h00092; 
        10'b0011111011: data <= 17'h1fff1; 
        10'b0011111100: data <= 17'h1ff99; 
        10'b0011111101: data <= 17'h1ffc4; 
        10'b0011111110: data <= 17'h1ff90; 
        10'b0011111111: data <= 17'h1ff0d; 
        10'b0100000000: data <= 17'h1fee8; 
        10'b0100000001: data <= 17'h1fefe; 
        10'b0100000010: data <= 17'h0001f; 
        10'b0100000011: data <= 17'h1ffee; 
        10'b0100000100: data <= 17'h000d7; 
        10'b0100000101: data <= 17'h000bb; 
        10'b0100000110: data <= 17'h000cb; 
        10'b0100000111: data <= 17'h0021e; 
        10'b0100001000: data <= 17'h0015e; 
        10'b0100001001: data <= 17'h1ff6f; 
        10'b0100001010: data <= 17'h1fe23; 
        10'b0100001011: data <= 17'h1fd55; 
        10'b0100001100: data <= 17'h1fd82; 
        10'b0100001101: data <= 17'h1fe8c; 
        10'b0100001110: data <= 17'h1ffab; 
        10'b0100001111: data <= 17'h1fffe; 
        10'b0100010000: data <= 17'h00122; 
        10'b0100010001: data <= 17'h0026d; 
        10'b0100010010: data <= 17'h00382; 
        10'b0100010011: data <= 17'h004cc; 
        10'b0100010100: data <= 17'h00608; 
        10'b0100010101: data <= 17'h003f6; 
        10'b0100010110: data <= 17'h000b6; 
        10'b0100010111: data <= 17'h1ffb8; 
        10'b0100011000: data <= 17'h1ffea; 
        10'b0100011001: data <= 17'h1ffb9; 
        10'b0100011010: data <= 17'h1ffa0; 
        10'b0100011011: data <= 17'h1ffb3; 
        10'b0100011100: data <= 17'h1ffaf; 
        10'b0100011101: data <= 17'h1ffcc; 
        10'b0100011110: data <= 17'h000ad; 
        10'b0100011111: data <= 17'h00143; 
        10'b0100100000: data <= 17'h001f8; 
        10'b0100100001: data <= 17'h0022d; 
        10'b0100100010: data <= 17'h00215; 
        10'b0100100011: data <= 17'h00285; 
        10'b0100100100: data <= 17'h00218; 
        10'b0100100101: data <= 17'h0019c; 
        10'b0100100110: data <= 17'h1ffa8; 
        10'b0100100111: data <= 17'h1feaf; 
        10'b0100101000: data <= 17'h1fdce; 
        10'b0100101001: data <= 17'h1fde0; 
        10'b0100101010: data <= 17'h1fdcd; 
        10'b0100101011: data <= 17'h1fd7e; 
        10'b0100101100: data <= 17'h1fe48; 
        10'b0100101101: data <= 17'h1ff77; 
        10'b0100101110: data <= 17'h0004b; 
        10'b0100101111: data <= 17'h0019c; 
        10'b0100110000: data <= 17'h00337; 
        10'b0100110001: data <= 17'h0026a; 
        10'b0100110010: data <= 17'h000d2; 
        10'b0100110011: data <= 17'h1ffb9; 
        10'b0100110100: data <= 17'h1ffa0; 
        10'b0100110101: data <= 17'h00001; 
        10'b0100110110: data <= 17'h1ffb2; 
        10'b0100110111: data <= 17'h1ffcd; 
        10'b0100111000: data <= 17'h1ffb0; 
        10'b0100111001: data <= 17'h1fff5; 
        10'b0100111010: data <= 17'h00113; 
        10'b0100111011: data <= 17'h00150; 
        10'b0100111100: data <= 17'h001e6; 
        10'b0100111101: data <= 17'h001c1; 
        10'b0100111110: data <= 17'h00148; 
        10'b0100111111: data <= 17'h0016a; 
        10'b0101000000: data <= 17'h00257; 
        10'b0101000001: data <= 17'h0022f; 
        10'b0101000010: data <= 17'h00009; 
        10'b0101000011: data <= 17'h1fea4; 
        10'b0101000100: data <= 17'h1fe50; 
        10'b0101000101: data <= 17'h1fe2f; 
        10'b0101000110: data <= 17'h1fd93; 
        10'b0101000111: data <= 17'h1fc9e; 
        10'b0101001000: data <= 17'h1fb17; 
        10'b0101001001: data <= 17'h1fb7e; 
        10'b0101001010: data <= 17'h1fc4e; 
        10'b0101001011: data <= 17'h1fd4e; 
        10'b0101001100: data <= 17'h1ff0b; 
        10'b0101001101: data <= 17'h0001b; 
        10'b0101001110: data <= 17'h00045; 
        10'b0101001111: data <= 17'h1ffd6; 
        10'b0101010000: data <= 17'h1ffd5; 
        10'b0101010001: data <= 17'h1ffdc; 
        10'b0101010010: data <= 17'h1ffcc; 
        10'b0101010011: data <= 17'h1ffb8; 
        10'b0101010100: data <= 17'h1ffc9; 
        10'b0101010101: data <= 17'h0008b; 
        10'b0101010110: data <= 17'h0013c; 
        10'b0101010111: data <= 17'h0011a; 
        10'b0101011000: data <= 17'h000cf; 
        10'b0101011001: data <= 17'h00077; 
        10'b0101011010: data <= 17'h0015e; 
        10'b0101011011: data <= 17'h002d4; 
        10'b0101011100: data <= 17'h002a5; 
        10'b0101011101: data <= 17'h002b6; 
        10'b0101011110: data <= 17'h00048; 
        10'b0101011111: data <= 17'h1fea0; 
        10'b0101100000: data <= 17'h1fd72; 
        10'b0101100001: data <= 17'h1fdee; 
        10'b0101100010: data <= 17'h1fe99; 
        10'b0101100011: data <= 17'h1fdfc; 
        10'b0101100100: data <= 17'h1fdb4; 
        10'b0101100101: data <= 17'h1fc30; 
        10'b0101100110: data <= 17'h1fba7; 
        10'b0101100111: data <= 17'h1fc39; 
        10'b0101101000: data <= 17'h1fd79; 
        10'b0101101001: data <= 17'h1ff48; 
        10'b0101101010: data <= 17'h0000a; 
        10'b0101101011: data <= 17'h1ffff; 
        10'b0101101100: data <= 17'h1ffda; 
        10'b0101101101: data <= 17'h1ffa4; 
        10'b0101101110: data <= 17'h1ff9f; 
        10'b0101101111: data <= 17'h1ffbc; 
        10'b0101110000: data <= 17'h1ffeb; 
        10'b0101110001: data <= 17'h00049; 
        10'b0101110010: data <= 17'h000d4; 
        10'b0101110011: data <= 17'h0009b; 
        10'b0101110100: data <= 17'h000b3; 
        10'b0101110101: data <= 17'h00094; 
        10'b0101110110: data <= 17'h001e7; 
        10'b0101110111: data <= 17'h00220; 
        10'b0101111000: data <= 17'h00195; 
        10'b0101111001: data <= 17'h0017a; 
        10'b0101111010: data <= 17'h1ffb4; 
        10'b0101111011: data <= 17'h1fe5d; 
        10'b0101111100: data <= 17'h1fd56; 
        10'b0101111101: data <= 17'h1fe98; 
        10'b0101111110: data <= 17'h1ff80; 
        10'b0101111111: data <= 17'h1ff6c; 
        10'b0110000000: data <= 17'h1ffba; 
        10'b0110000001: data <= 17'h1feec; 
        10'b0110000010: data <= 17'h1fe0c; 
        10'b0110000011: data <= 17'h1fd26; 
        10'b0110000100: data <= 17'h1fdda; 
        10'b0110000101: data <= 17'h1ffa1; 
        10'b0110000110: data <= 17'h1ff98; 
        10'b0110000111: data <= 17'h1fff1; 
        10'b0110001000: data <= 17'h1ffdb; 
        10'b0110001001: data <= 17'h1ff9d; 
        10'b0110001010: data <= 17'h1ffcf; 
        10'b0110001011: data <= 17'h1ff85; 
        10'b0110001100: data <= 17'h1ffd7; 
        10'b0110001101: data <= 17'h1ffd3; 
        10'b0110001110: data <= 17'h1fffe; 
        10'b0110001111: data <= 17'h1ffe9; 
        10'b0110010000: data <= 17'h000e0; 
        10'b0110010001: data <= 17'h00162; 
        10'b0110010010: data <= 17'h001a9; 
        10'b0110010011: data <= 17'h00051; 
        10'b0110010100: data <= 17'h00090; 
        10'b0110010101: data <= 17'h1ffe5; 
        10'b0110010110: data <= 17'h1fed0; 
        10'b0110010111: data <= 17'h1fea2; 
        10'b0110011000: data <= 17'h1fe1a; 
        10'b0110011001: data <= 17'h1fe52; 
        10'b0110011010: data <= 17'h1fe6d; 
        10'b0110011011: data <= 17'h1ff3e; 
        10'b0110011100: data <= 17'h1ff58; 
        10'b0110011101: data <= 17'h1ff67; 
        10'b0110011110: data <= 17'h1ffa3; 
        10'b0110011111: data <= 17'h1fe6f; 
        10'b0110100000: data <= 17'h1fef2; 
        10'b0110100001: data <= 17'h1ff79; 
        10'b0110100010: data <= 17'h1ffd0; 
        10'b0110100011: data <= 17'h1ff88; 
        10'b0110100100: data <= 17'h1ff95; 
        10'b0110100101: data <= 17'h00010; 
        10'b0110100110: data <= 17'h1ff8c; 
        10'b0110100111: data <= 17'h1ffd1; 
        10'b0110101000: data <= 17'h1ff54; 
        10'b0110101001: data <= 17'h1fefe; 
        10'b0110101010: data <= 17'h1fe97; 
        10'b0110101011: data <= 17'h1ff11; 
        10'b0110101100: data <= 17'h00057; 
        10'b0110101101: data <= 17'h0018f; 
        10'b0110101110: data <= 17'h000be; 
        10'b0110101111: data <= 17'h000af; 
        10'b0110110000: data <= 17'h00097; 
        10'b0110110001: data <= 17'h1ff78; 
        10'b0110110010: data <= 17'h1fe3d; 
        10'b0110110011: data <= 17'h1fdf9; 
        10'b0110110100: data <= 17'h1fe2b; 
        10'b0110110101: data <= 17'h1fe20; 
        10'b0110110110: data <= 17'h1feae; 
        10'b0110110111: data <= 17'h1ffef; 
        10'b0110111000: data <= 17'h1ff8d; 
        10'b0110111001: data <= 17'h1ff9f; 
        10'b0110111010: data <= 17'h1ff8c; 
        10'b0110111011: data <= 17'h1ff7b; 
        10'b0110111100: data <= 17'h1ffa2; 
        10'b0110111101: data <= 17'h1fffd; 
        10'b0110111110: data <= 17'h00013; 
        10'b0110111111: data <= 17'h1ffb8; 
        10'b0111000000: data <= 17'h1ffbf; 
        10'b0111000001: data <= 17'h1ffd6; 
        10'b0111000010: data <= 17'h1ffe4; 
        10'b0111000011: data <= 17'h1ff8d; 
        10'b0111000100: data <= 17'h1ffbd; 
        10'b0111000101: data <= 17'h1fedb; 
        10'b0111000110: data <= 17'h1fdb5; 
        10'b0111000111: data <= 17'h1fd4a; 
        10'b0111001000: data <= 17'h1fe2a; 
        10'b0111001001: data <= 17'h1fefc; 
        10'b0111001010: data <= 17'h1ff99; 
        10'b0111001011: data <= 17'h1ff6c; 
        10'b0111001100: data <= 17'h1ff9f; 
        10'b0111001101: data <= 17'h1fec0; 
        10'b0111001110: data <= 17'h1fd98; 
        10'b0111001111: data <= 17'h1fe0b; 
        10'b0111010000: data <= 17'h1fe94; 
        10'b0111010001: data <= 17'h1ff7d; 
        10'b0111010010: data <= 17'h1ff85; 
        10'b0111010011: data <= 17'h00014; 
        10'b0111010100: data <= 17'h00065; 
        10'b0111010101: data <= 17'h00010; 
        10'b0111010110: data <= 17'h0006e; 
        10'b0111010111: data <= 17'h00019; 
        10'b0111011000: data <= 17'h00011; 
        10'b0111011001: data <= 17'h00010; 
        10'b0111011010: data <= 17'h1ffbb; 
        10'b0111011011: data <= 17'h1ffc0; 
        10'b0111011100: data <= 17'h1ffb3; 
        10'b0111011101: data <= 17'h1fffb; 
        10'b0111011110: data <= 17'h00000; 
        10'b0111011111: data <= 17'h00008; 
        10'b0111100000: data <= 17'h1ffb6; 
        10'b0111100001: data <= 17'h00015; 
        10'b0111100010: data <= 17'h0002b; 
        10'b0111100011: data <= 17'h1fe35; 
        10'b0111100100: data <= 17'h1fcc2; 
        10'b0111100101: data <= 17'h1fcf8; 
        10'b0111100110: data <= 17'h1fdd4; 
        10'b0111100111: data <= 17'h1feb1; 
        10'b0111101000: data <= 17'h1fdf5; 
        10'b0111101001: data <= 17'h1fd5d; 
        10'b0111101010: data <= 17'h1fd70; 
        10'b0111101011: data <= 17'h1fed5; 
        10'b0111101100: data <= 17'h1ff7d; 
        10'b0111101101: data <= 17'h000c6; 
        10'b0111101110: data <= 17'h0012f; 
        10'b0111101111: data <= 17'h000c6; 
        10'b0111110000: data <= 17'h000c8; 
        10'b0111110001: data <= 17'h0003a; 
        10'b0111110010: data <= 17'h00007; 
        10'b0111110011: data <= 17'h0006e; 
        10'b0111110100: data <= 17'h00070; 
        10'b0111110101: data <= 17'h1ffa1; 
        10'b0111110110: data <= 17'h1fffc; 
        10'b0111110111: data <= 17'h00003; 
        10'b0111111000: data <= 17'h0000b; 
        10'b0111111001: data <= 17'h1ffaf; 
        10'b0111111010: data <= 17'h1ffcd; 
        10'b0111111011: data <= 17'h1ffbf; 
        10'b0111111100: data <= 17'h000a4; 
        10'b0111111101: data <= 17'h000d9; 
        10'b0111111110: data <= 17'h00203; 
        10'b0111111111: data <= 17'h0005b; 
        10'b1000000000: data <= 17'h1fe10; 
        10'b1000000001: data <= 17'h1fd2e; 
        10'b1000000010: data <= 17'h1fc4a; 
        10'b1000000011: data <= 17'h1fcaf; 
        10'b1000000100: data <= 17'h1fd9f; 
        10'b1000000101: data <= 17'h1fea4; 
        10'b1000000110: data <= 17'h1ff52; 
        10'b1000000111: data <= 17'h1ffb7; 
        10'b1000001000: data <= 17'h1fff3; 
        10'b1000001001: data <= 17'h000e9; 
        10'b1000001010: data <= 17'h00075; 
        10'b1000001011: data <= 17'h000d0; 
        10'b1000001100: data <= 17'h0008c; 
        10'b1000001101: data <= 17'h000cb; 
        10'b1000001110: data <= 17'h000a7; 
        10'b1000001111: data <= 17'h000e7; 
        10'b1000010000: data <= 17'h00078; 
        10'b1000010001: data <= 17'h00009; 
        10'b1000010010: data <= 17'h1ffa8; 
        10'b1000010011: data <= 17'h1ffe4; 
        10'b1000010100: data <= 17'h00001; 
        10'b1000010101: data <= 17'h1ffaf; 
        10'b1000010110: data <= 17'h1ffd4; 
        10'b1000010111: data <= 17'h00011; 
        10'b1000011000: data <= 17'h000f9; 
        10'b1000011001: data <= 17'h001aa; 
        10'b1000011010: data <= 17'h0023d; 
        10'b1000011011: data <= 17'h00182; 
        10'b1000011100: data <= 17'h000f4; 
        10'b1000011101: data <= 17'h0004f; 
        10'b1000011110: data <= 17'h1ff4a; 
        10'b1000011111: data <= 17'h1ff3d; 
        10'b1000100000: data <= 17'h00010; 
        10'b1000100001: data <= 17'h000ea; 
        10'b1000100010: data <= 17'h00057; 
        10'b1000100011: data <= 17'h0007c; 
        10'b1000100100: data <= 17'h0007e; 
        10'b1000100101: data <= 17'h1ffd8; 
        10'b1000100110: data <= 17'h0005a; 
        10'b1000100111: data <= 17'h00058; 
        10'b1000101000: data <= 17'h00013; 
        10'b1000101001: data <= 17'h00097; 
        10'b1000101010: data <= 17'h00104; 
        10'b1000101011: data <= 17'h000be; 
        10'b1000101100: data <= 17'h00010; 
        10'b1000101101: data <= 17'h1fffd; 
        10'b1000101110: data <= 17'h1ffff; 
        10'b1000101111: data <= 17'h1ff9a; 
        10'b1000110000: data <= 17'h1fffb; 
        10'b1000110001: data <= 17'h1ff89; 
        10'b1000110010: data <= 17'h1ffc7; 
        10'b1000110011: data <= 17'h1ffa7; 
        10'b1000110100: data <= 17'h00021; 
        10'b1000110101: data <= 17'h00118; 
        10'b1000110110: data <= 17'h00145; 
        10'b1000110111: data <= 17'h0018c; 
        10'b1000111000: data <= 17'h0022b; 
        10'b1000111001: data <= 17'h001d5; 
        10'b1000111010: data <= 17'h0019c; 
        10'b1000111011: data <= 17'h00258; 
        10'b1000111100: data <= 17'h00176; 
        10'b1000111101: data <= 17'h00118; 
        10'b1000111110: data <= 17'h1ffb1; 
        10'b1000111111: data <= 17'h1ffb8; 
        10'b1001000000: data <= 17'h000ce; 
        10'b1001000001: data <= 17'h0006a; 
        10'b1001000010: data <= 17'h000ad; 
        10'b1001000011: data <= 17'h000e4; 
        10'b1001000100: data <= 17'h000c8; 
        10'b1001000101: data <= 17'h0009d; 
        10'b1001000110: data <= 17'h00177; 
        10'b1001000111: data <= 17'h00119; 
        10'b1001001000: data <= 17'h1ffdb; 
        10'b1001001001: data <= 17'h1ff8b; 
        10'b1001001010: data <= 17'h1ffd7; 
        10'b1001001011: data <= 17'h1ffb6; 
        10'b1001001100: data <= 17'h1ffab; 
        10'b1001001101: data <= 17'h00003; 
        10'b1001001110: data <= 17'h1ff84; 
        10'b1001001111: data <= 17'h1ffd1; 
        10'b1001010000: data <= 17'h0006e; 
        10'b1001010001: data <= 17'h1ffdd; 
        10'b1001010010: data <= 17'h00086; 
        10'b1001010011: data <= 17'h0016a; 
        10'b1001010100: data <= 17'h0020b; 
        10'b1001010101: data <= 17'h00156; 
        10'b1001010110: data <= 17'h00122; 
        10'b1001010111: data <= 17'h0009c; 
        10'b1001011000: data <= 17'h000ca; 
        10'b1001011001: data <= 17'h0007e; 
        10'b1001011010: data <= 17'h00083; 
        10'b1001011011: data <= 17'h000a0; 
        10'b1001011100: data <= 17'h0002a; 
        10'b1001011101: data <= 17'h00081; 
        10'b1001011110: data <= 17'h00042; 
        10'b1001011111: data <= 17'h000cf; 
        10'b1001100000: data <= 17'h000cc; 
        10'b1001100001: data <= 17'h00155; 
        10'b1001100010: data <= 17'h001a4; 
        10'b1001100011: data <= 17'h0005b; 
        10'b1001100100: data <= 17'h00004; 
        10'b1001100101: data <= 17'h1ff9c; 
        10'b1001100110: data <= 17'h1ffb7; 
        10'b1001100111: data <= 17'h1ffb8; 
        10'b1001101000: data <= 17'h1ffe7; 
        10'b1001101001: data <= 17'h1ff8f; 
        10'b1001101010: data <= 17'h1ffc5; 
        10'b1001101011: data <= 17'h1ffb7; 
        10'b1001101100: data <= 17'h00028; 
        10'b1001101101: data <= 17'h1ffc8; 
        10'b1001101110: data <= 17'h1ff85; 
        10'b1001101111: data <= 17'h1ffea; 
        10'b1001110000: data <= 17'h000cb; 
        10'b1001110001: data <= 17'h00129; 
        10'b1001110010: data <= 17'h00034; 
        10'b1001110011: data <= 17'h00107; 
        10'b1001110100: data <= 17'h001aa; 
        10'b1001110101: data <= 17'h0020e; 
        10'b1001110110: data <= 17'h0010c; 
        10'b1001110111: data <= 17'h00028; 
        10'b1001111000: data <= 17'h0001e; 
        10'b1001111001: data <= 17'h00042; 
        10'b1001111010: data <= 17'h0008a; 
        10'b1001111011: data <= 17'h00089; 
        10'b1001111100: data <= 17'h000eb; 
        10'b1001111101: data <= 17'h000d4; 
        10'b1001111110: data <= 17'h000dd; 
        10'b1001111111: data <= 17'h0004e; 
        10'b1010000000: data <= 17'h1fff5; 
        10'b1010000001: data <= 17'h0000c; 
        10'b1010000010: data <= 17'h1ffd5; 
        10'b1010000011: data <= 17'h1ffe3; 
        10'b1010000100: data <= 17'h1ffa2; 
        10'b1010000101: data <= 17'h1ffd2; 
        10'b1010000110: data <= 17'h1ffe6; 
        10'b1010000111: data <= 17'h1ffdc; 
        10'b1010001000: data <= 17'h1ffa7; 
        10'b1010001001: data <= 17'h1ffc5; 
        10'b1010001010: data <= 17'h1ff4e; 
        10'b1010001011: data <= 17'h1ffaf; 
        10'b1010001100: data <= 17'h000a1; 
        10'b1010001101: data <= 17'h0009e; 
        10'b1010001110: data <= 17'h0009d; 
        10'b1010001111: data <= 17'h00118; 
        10'b1010010000: data <= 17'h0010d; 
        10'b1010010001: data <= 17'h000b8; 
        10'b1010010010: data <= 17'h000d4; 
        10'b1010010011: data <= 17'h000c2; 
        10'b1010010100: data <= 17'h000be; 
        10'b1010010101: data <= 17'h00057; 
        10'b1010010110: data <= 17'h1ff9c; 
        10'b1010010111: data <= 17'h1fff2; 
        10'b1010011000: data <= 17'h0005d; 
        10'b1010011001: data <= 17'h00026; 
        10'b1010011010: data <= 17'h0007d; 
        10'b1010011011: data <= 17'h1ffb2; 
        10'b1010011100: data <= 17'h00015; 
        10'b1010011101: data <= 17'h1ffc0; 
        10'b1010011110: data <= 17'h1ffbf; 
        10'b1010011111: data <= 17'h00013; 
        10'b1010100000: data <= 17'h1fff7; 
        10'b1010100001: data <= 17'h1ffc3; 
        10'b1010100010: data <= 17'h1ffb9; 
        10'b1010100011: data <= 17'h00016; 
        10'b1010100100: data <= 17'h1ff86; 
        10'b1010100101: data <= 17'h1ff7f; 
        10'b1010100110: data <= 17'h1ffd2; 
        10'b1010100111: data <= 17'h1ffe8; 
        10'b1010101000: data <= 17'h1fff9; 
        10'b1010101001: data <= 17'h000d0; 
        10'b1010101010: data <= 17'h0010e; 
        10'b1010101011: data <= 17'h000d0; 
        10'b1010101100: data <= 17'h00087; 
        10'b1010101101: data <= 17'h000bc; 
        10'b1010101110: data <= 17'h0015b; 
        10'b1010101111: data <= 17'h0011f; 
        10'b1010110000: data <= 17'h000ab; 
        10'b1010110001: data <= 17'h00053; 
        10'b1010110010: data <= 17'h0009f; 
        10'b1010110011: data <= 17'h00067; 
        10'b1010110100: data <= 17'h1fffa; 
        10'b1010110101: data <= 17'h1fff1; 
        10'b1010110110: data <= 17'h1ffda; 
        10'b1010110111: data <= 17'h00007; 
        10'b1010111000: data <= 17'h1ffac; 
        10'b1010111001: data <= 17'h1ffe2; 
        10'b1010111010: data <= 17'h0000d; 
        10'b1010111011: data <= 17'h1ff99; 
        10'b1010111100: data <= 17'h1ffd2; 
        10'b1010111101: data <= 17'h00004; 
        10'b1010111110: data <= 17'h0000c; 
        10'b1010111111: data <= 17'h1ff94; 
        10'b1011000000: data <= 17'h1ffff; 
        10'b1011000001: data <= 17'h1ffdf; 
        10'b1011000010: data <= 17'h1ff80; 
        10'b1011000011: data <= 17'h1ffd1; 
        10'b1011000100: data <= 17'h1ff8d; 
        10'b1011000101: data <= 17'h00044; 
        10'b1011000110: data <= 17'h00032; 
        10'b1011000111: data <= 17'h0008d; 
        10'b1011001000: data <= 17'h0008c; 
        10'b1011001001: data <= 17'h000f6; 
        10'b1011001010: data <= 17'h0000d; 
        10'b1011001011: data <= 17'h00049; 
        10'b1011001100: data <= 17'h0003e; 
        10'b1011001101: data <= 17'h00078; 
        10'b1011001110: data <= 17'h1ffaf; 
        10'b1011001111: data <= 17'h1fffc; 
        10'b1011010000: data <= 17'h1ff7a; 
        10'b1011010001: data <= 17'h0000c; 
        10'b1011010010: data <= 17'h1ffce; 
        10'b1011010011: data <= 17'h1ffa6; 
        10'b1011010100: data <= 17'h1fff5; 
        10'b1011010101: data <= 17'h00006; 
        10'b1011010110: data <= 17'h1ff8e; 
        10'b1011010111: data <= 17'h1ffc4; 
        10'b1011011000: data <= 17'h1ffdc; 
        10'b1011011001: data <= 17'h1ffd9; 
        10'b1011011010: data <= 17'h1ffac; 
        10'b1011011011: data <= 17'h1ffc0; 
        10'b1011011100: data <= 17'h1ffb9; 
        10'b1011011101: data <= 17'h1ffc6; 
        10'b1011011110: data <= 17'h1ffeb; 
        10'b1011011111: data <= 17'h1ffad; 
        10'b1011100000: data <= 17'h1ff92; 
        10'b1011100001: data <= 17'h1ffc7; 
        10'b1011100010: data <= 17'h1ffb5; 
        10'b1011100011: data <= 17'h1fff2; 
        10'b1011100100: data <= 17'h00002; 
        10'b1011100101: data <= 17'h1ffe3; 
        10'b1011100110: data <= 17'h1ffb0; 
        10'b1011100111: data <= 17'h1ffd7; 
        10'b1011101000: data <= 17'h1ffee; 
        10'b1011101001: data <= 17'h1ffac; 
        10'b1011101010: data <= 17'h1ff5e; 
        10'b1011101011: data <= 17'h1ff7d; 
        10'b1011101100: data <= 17'h1ffe4; 
        10'b1011101101: data <= 17'h1ffe4; 
        10'b1011101110: data <= 17'h1ffb6; 
        10'b1011101111: data <= 17'h1ffea; 
        10'b1011110000: data <= 17'h1ffc9; 
        10'b1011110001: data <= 17'h1ffda; 
        10'b1011110010: data <= 17'h1ffbc; 
        10'b1011110011: data <= 17'h1ff8e; 
        10'b1011110100: data <= 17'h1ffe7; 
        10'b1011110101: data <= 17'h1fff0; 
        10'b1011110110: data <= 17'h1fff5; 
        10'b1011110111: data <= 17'h1ffe0; 
        10'b1011111000: data <= 17'h1ff9e; 
        10'b1011111001: data <= 17'h1fffa; 
        10'b1011111010: data <= 17'h1ffbe; 
        10'b1011111011: data <= 17'h1ffb8; 
        10'b1011111100: data <= 17'h00018; 
        10'b1011111101: data <= 17'h1ffbb; 
        10'b1011111110: data <= 17'h1ffb2; 
        10'b1011111111: data <= 17'h1fff7; 
        10'b1100000000: data <= 17'h1ffd6; 
        10'b1100000001: data <= 17'h1ff88; 
        10'b1100000010: data <= 17'h00003; 
        10'b1100000011: data <= 17'h1ffdb; 
        10'b1100000100: data <= 17'h1ff93; 
        10'b1100000101: data <= 17'h1ff87; 
        10'b1100000110: data <= 17'h1ffa6; 
        10'b1100000111: data <= 17'h1ff86; 
        10'b1100001000: data <= 17'h1fffe; 
        10'b1100001001: data <= 17'h1ffbd; 
        10'b1100001010: data <= 17'h00016; 
        10'b1100001011: data <= 17'h1ff98; 
        10'b1100001100: data <= 17'h1ffe1; 
        10'b1100001101: data <= 17'h1ffcc; 
        10'b1100001110: data <= 17'h1ffa0; 
        10'b1100001111: data <= 17'h1fff1; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 12) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 18'h3ff72; 
        10'b0000000001: data <= 18'h3ffec; 
        10'b0000000010: data <= 18'h3ffec; 
        10'b0000000011: data <= 18'h3ff41; 
        10'b0000000100: data <= 18'h3ffa6; 
        10'b0000000101: data <= 18'h3ff8e; 
        10'b0000000110: data <= 18'h3ffff; 
        10'b0000000111: data <= 18'h3ff85; 
        10'b0000001000: data <= 18'h3ffcd; 
        10'b0000001001: data <= 18'h00029; 
        10'b0000001010: data <= 18'h3ffcd; 
        10'b0000001011: data <= 18'h3ffc9; 
        10'b0000001100: data <= 18'h3ff6e; 
        10'b0000001101: data <= 18'h3fff7; 
        10'b0000001110: data <= 18'h3ff3e; 
        10'b0000001111: data <= 18'h3ff60; 
        10'b0000010000: data <= 18'h3ff24; 
        10'b0000010001: data <= 18'h3ff4d; 
        10'b0000010010: data <= 18'h3ffe6; 
        10'b0000010011: data <= 18'h3ffcf; 
        10'b0000010100: data <= 18'h3ff22; 
        10'b0000010101: data <= 18'h3ffab; 
        10'b0000010110: data <= 18'h3ffc3; 
        10'b0000010111: data <= 18'h3ff92; 
        10'b0000011000: data <= 18'h3ff2e; 
        10'b0000011001: data <= 18'h3ffb1; 
        10'b0000011010: data <= 18'h3ffc2; 
        10'b0000011011: data <= 18'h3ff78; 
        10'b0000011100: data <= 18'h3fff3; 
        10'b0000011101: data <= 18'h3ff17; 
        10'b0000011110: data <= 18'h3fffe; 
        10'b0000011111: data <= 18'h3ff38; 
        10'b0000100000: data <= 18'h3fff7; 
        10'b0000100001: data <= 18'h3ff80; 
        10'b0000100010: data <= 18'h3ffbe; 
        10'b0000100011: data <= 18'h3ff7a; 
        10'b0000100100: data <= 18'h3ff59; 
        10'b0000100101: data <= 18'h3ffc3; 
        10'b0000100110: data <= 18'h00015; 
        10'b0000100111: data <= 18'h3ff3d; 
        10'b0000101000: data <= 18'h3ff79; 
        10'b0000101001: data <= 18'h3ff52; 
        10'b0000101010: data <= 18'h3ff20; 
        10'b0000101011: data <= 18'h3ffdb; 
        10'b0000101100: data <= 18'h3ff68; 
        10'b0000101101: data <= 18'h3ff4f; 
        10'b0000101110: data <= 18'h3ff6d; 
        10'b0000101111: data <= 18'h3ff63; 
        10'b0000110000: data <= 18'h3ffce; 
        10'b0000110001: data <= 18'h3ff35; 
        10'b0000110010: data <= 18'h3fffd; 
        10'b0000110011: data <= 18'h3ff43; 
        10'b0000110100: data <= 18'h00003; 
        10'b0000110101: data <= 18'h3fff1; 
        10'b0000110110: data <= 18'h3ff4b; 
        10'b0000110111: data <= 18'h3ff9c; 
        10'b0000111000: data <= 18'h3ff9e; 
        10'b0000111001: data <= 18'h3ffd5; 
        10'b0000111010: data <= 18'h3ff79; 
        10'b0000111011: data <= 18'h3ff22; 
        10'b0000111100: data <= 18'h3ff49; 
        10'b0000111101: data <= 18'h3ffb2; 
        10'b0000111110: data <= 18'h3fff8; 
        10'b0000111111: data <= 18'h3ffc4; 
        10'b0001000000: data <= 18'h3ff5f; 
        10'b0001000001: data <= 18'h3ff85; 
        10'b0001000010: data <= 18'h0001f; 
        10'b0001000011: data <= 18'h3ff13; 
        10'b0001000100: data <= 18'h3fff5; 
        10'b0001000101: data <= 18'h3ff59; 
        10'b0001000110: data <= 18'h3ff27; 
        10'b0001000111: data <= 18'h3ff4f; 
        10'b0001001000: data <= 18'h3ff72; 
        10'b0001001001: data <= 18'h3ffae; 
        10'b0001001010: data <= 18'h3ff85; 
        10'b0001001011: data <= 18'h3ff87; 
        10'b0001001100: data <= 18'h00036; 
        10'b0001001101: data <= 18'h00006; 
        10'b0001001110: data <= 18'h00017; 
        10'b0001001111: data <= 18'h3ff54; 
        10'b0001010000: data <= 18'h3ff21; 
        10'b0001010001: data <= 18'h3ff91; 
        10'b0001010010: data <= 18'h3fff2; 
        10'b0001010011: data <= 18'h3ffc3; 
        10'b0001010100: data <= 18'h3ffd6; 
        10'b0001010101: data <= 18'h3ffc0; 
        10'b0001010110: data <= 18'h3ff4b; 
        10'b0001010111: data <= 18'h3fff4; 
        10'b0001011000: data <= 18'h3ff39; 
        10'b0001011001: data <= 18'h3ff7c; 
        10'b0001011010: data <= 18'h3ff13; 
        10'b0001011011: data <= 18'h3ff65; 
        10'b0001011100: data <= 18'h3ff24; 
        10'b0001011101: data <= 18'h3ff63; 
        10'b0001011110: data <= 18'h3fe81; 
        10'b0001011111: data <= 18'h3fe17; 
        10'b0001100000: data <= 18'h3fee9; 
        10'b0001100001: data <= 18'h3fefa; 
        10'b0001100010: data <= 18'h3febe; 
        10'b0001100011: data <= 18'h3ff95; 
        10'b0001100100: data <= 18'h3ffd2; 
        10'b0001100101: data <= 18'h3ff03; 
        10'b0001100110: data <= 18'h3ff68; 
        10'b0001100111: data <= 18'h3ffd0; 
        10'b0001101000: data <= 18'h3ffde; 
        10'b0001101001: data <= 18'h3ff97; 
        10'b0001101010: data <= 18'h3ff00; 
        10'b0001101011: data <= 18'h3ff54; 
        10'b0001101100: data <= 18'h3fecb; 
        10'b0001101101: data <= 18'h00024; 
        10'b0001101110: data <= 18'h00016; 
        10'b0001101111: data <= 18'h3ff36; 
        10'b0001110000: data <= 18'h3ff28; 
        10'b0001110001: data <= 18'h3ff7a; 
        10'b0001110010: data <= 18'h00016; 
        10'b0001110011: data <= 18'h0000c; 
        10'b0001110100: data <= 18'h0001e; 
        10'b0001110101: data <= 18'h3ff65; 
        10'b0001110110: data <= 18'h3ff5a; 
        10'b0001110111: data <= 18'h3fea6; 
        10'b0001111000: data <= 18'h3fdb9; 
        10'b0001111001: data <= 18'h3fcfa; 
        10'b0001111010: data <= 18'h3fb95; 
        10'b0001111011: data <= 18'h3fd2e; 
        10'b0001111100: data <= 18'h3fd28; 
        10'b0001111101: data <= 18'h3fc2f; 
        10'b0001111110: data <= 18'h3fde6; 
        10'b0001111111: data <= 18'h3fffd; 
        10'b0010000000: data <= 18'h3ffc0; 
        10'b0010000001: data <= 18'h000b6; 
        10'b0010000010: data <= 18'h3ffc9; 
        10'b0010000011: data <= 18'h3feeb; 
        10'b0010000100: data <= 18'h3fe95; 
        10'b0010000101: data <= 18'h3ff40; 
        10'b0010000110: data <= 18'h3ff63; 
        10'b0010000111: data <= 18'h3ff92; 
        10'b0010001000: data <= 18'h3ff78; 
        10'b0010001001: data <= 18'h00033; 
        10'b0010001010: data <= 18'h0001d; 
        10'b0010001011: data <= 18'h3ff9c; 
        10'b0010001100: data <= 18'h3ffae; 
        10'b0010001101: data <= 18'h00033; 
        10'b0010001110: data <= 18'h3ff51; 
        10'b0010001111: data <= 18'h3ff37; 
        10'b0010010000: data <= 18'h3ff6b; 
        10'b0010010001: data <= 18'h3fe9f; 
        10'b0010010010: data <= 18'h3fdea; 
        10'b0010010011: data <= 18'h3fdfc; 
        10'b0010010100: data <= 18'h3feae; 
        10'b0010010101: data <= 18'h3ffc1; 
        10'b0010010110: data <= 18'h00072; 
        10'b0010010111: data <= 18'h0007b; 
        10'b0010011000: data <= 18'h3ff49; 
        10'b0010011001: data <= 18'h3fefa; 
        10'b0010011010: data <= 18'h3ff62; 
        10'b0010011011: data <= 18'h3ffb6; 
        10'b0010011100: data <= 18'h00105; 
        10'b0010011101: data <= 18'h0010b; 
        10'b0010011110: data <= 18'h001fb; 
        10'b0010011111: data <= 18'h0013c; 
        10'b0010100000: data <= 18'h00132; 
        10'b0010100001: data <= 18'h00189; 
        10'b0010100010: data <= 18'h002d5; 
        10'b0010100011: data <= 18'h00269; 
        10'b0010100100: data <= 18'h001b1; 
        10'b0010100101: data <= 18'h000ef; 
        10'b0010100110: data <= 18'h00095; 
        10'b0010100111: data <= 18'h00038; 
        10'b0010101000: data <= 18'h3ff3f; 
        10'b0010101001: data <= 18'h3ff2e; 
        10'b0010101010: data <= 18'h0001b; 
        10'b0010101011: data <= 18'h3ff36; 
        10'b0010101100: data <= 18'h3fefb; 
        10'b0010101101: data <= 18'h3fd91; 
        10'b0010101110: data <= 18'h3fee8; 
        10'b0010101111: data <= 18'h3ffdf; 
        10'b0010110000: data <= 18'h3ffea; 
        10'b0010110001: data <= 18'h000fd; 
        10'b0010110010: data <= 18'h0020c; 
        10'b0010110011: data <= 18'h001b4; 
        10'b0010110100: data <= 18'h0004a; 
        10'b0010110101: data <= 18'h000a1; 
        10'b0010110110: data <= 18'h3ffb8; 
        10'b0010110111: data <= 18'h3ff07; 
        10'b0010111000: data <= 18'h3ff6a; 
        10'b0010111001: data <= 18'h3ff81; 
        10'b0010111010: data <= 18'h00006; 
        10'b0010111011: data <= 18'h001f2; 
        10'b0010111100: data <= 18'h0011d; 
        10'b0010111101: data <= 18'h00144; 
        10'b0010111110: data <= 18'h003de; 
        10'b0010111111: data <= 18'h004a6; 
        10'b0011000000: data <= 18'h0053a; 
        10'b0011000001: data <= 18'h002c4; 
        10'b0011000010: data <= 18'h0015e; 
        10'b0011000011: data <= 18'h00055; 
        10'b0011000100: data <= 18'h3ff93; 
        10'b0011000101: data <= 18'h3ffc5; 
        10'b0011000110: data <= 18'h3ffab; 
        10'b0011000111: data <= 18'h3feff; 
        10'b0011001000: data <= 18'h3fd2c; 
        10'b0011001001: data <= 18'h3fcaf; 
        10'b0011001010: data <= 18'h3fdfb; 
        10'b0011001011: data <= 18'h00043; 
        10'b0011001100: data <= 18'h00153; 
        10'b0011001101: data <= 18'h00299; 
        10'b0011001110: data <= 18'h00287; 
        10'b0011001111: data <= 18'h00235; 
        10'b0011010000: data <= 18'h000a4; 
        10'b0011010001: data <= 18'h3ffca; 
        10'b0011010010: data <= 18'h3ff4b; 
        10'b0011010011: data <= 18'h0000c; 
        10'b0011010100: data <= 18'h00118; 
        10'b0011010101: data <= 18'h000fd; 
        10'b0011010110: data <= 18'h00141; 
        10'b0011010111: data <= 18'h002cd; 
        10'b0011011000: data <= 18'h0026c; 
        10'b0011011001: data <= 18'h002e5; 
        10'b0011011010: data <= 18'h0040c; 
        10'b0011011011: data <= 18'h0056e; 
        10'b0011011100: data <= 18'h006a1; 
        10'b0011011101: data <= 18'h004c9; 
        10'b0011011110: data <= 18'h000bd; 
        10'b0011011111: data <= 18'h3ffe3; 
        10'b0011100000: data <= 18'h3ffd0; 
        10'b0011100001: data <= 18'h0002d; 
        10'b0011100010: data <= 18'h3fffc; 
        10'b0011100011: data <= 18'h3fea2; 
        10'b0011100100: data <= 18'h3fbee; 
        10'b0011100101: data <= 18'h3fc85; 
        10'b0011100110: data <= 18'h3fd7b; 
        10'b0011100111: data <= 18'h00028; 
        10'b0011101000: data <= 18'h001f8; 
        10'b0011101001: data <= 18'h00094; 
        10'b0011101010: data <= 18'h0010f; 
        10'b0011101011: data <= 18'h0020e; 
        10'b0011101100: data <= 18'h00141; 
        10'b0011101101: data <= 18'h3fe97; 
        10'b0011101110: data <= 18'h3fce9; 
        10'b0011101111: data <= 18'h3fe21; 
        10'b0011110000: data <= 18'h3feda; 
        10'b0011110001: data <= 18'h0001c; 
        10'b0011110010: data <= 18'h00051; 
        10'b0011110011: data <= 18'h00255; 
        10'b0011110100: data <= 18'h00276; 
        10'b0011110101: data <= 18'h00382; 
        10'b0011110110: data <= 18'h0058c; 
        10'b0011110111: data <= 18'h00742; 
        10'b0011111000: data <= 18'h009ae; 
        10'b0011111001: data <= 18'h00641; 
        10'b0011111010: data <= 18'h00124; 
        10'b0011111011: data <= 18'h3ffe2; 
        10'b0011111100: data <= 18'h3ff33; 
        10'b0011111101: data <= 18'h3ff88; 
        10'b0011111110: data <= 18'h3ff20; 
        10'b0011111111: data <= 18'h3fe19; 
        10'b0100000000: data <= 18'h3fdd1; 
        10'b0100000001: data <= 18'h3fdfb; 
        10'b0100000010: data <= 18'h0003f; 
        10'b0100000011: data <= 18'h3ffdc; 
        10'b0100000100: data <= 18'h001ae; 
        10'b0100000101: data <= 18'h00176; 
        10'b0100000110: data <= 18'h00197; 
        10'b0100000111: data <= 18'h0043d; 
        10'b0100001000: data <= 18'h002bc; 
        10'b0100001001: data <= 18'h3fede; 
        10'b0100001010: data <= 18'h3fc47; 
        10'b0100001011: data <= 18'h3faa9; 
        10'b0100001100: data <= 18'h3fb03; 
        10'b0100001101: data <= 18'h3fd19; 
        10'b0100001110: data <= 18'h3ff56; 
        10'b0100001111: data <= 18'h3fffb; 
        10'b0100010000: data <= 18'h00244; 
        10'b0100010001: data <= 18'h004d9; 
        10'b0100010010: data <= 18'h00704; 
        10'b0100010011: data <= 18'h00999; 
        10'b0100010100: data <= 18'h00c0f; 
        10'b0100010101: data <= 18'h007ed; 
        10'b0100010110: data <= 18'h0016b; 
        10'b0100010111: data <= 18'h3ff71; 
        10'b0100011000: data <= 18'h3ffd4; 
        10'b0100011001: data <= 18'h3ff72; 
        10'b0100011010: data <= 18'h3ff41; 
        10'b0100011011: data <= 18'h3ff66; 
        10'b0100011100: data <= 18'h3ff5d; 
        10'b0100011101: data <= 18'h3ff97; 
        10'b0100011110: data <= 18'h0015a; 
        10'b0100011111: data <= 18'h00285; 
        10'b0100100000: data <= 18'h003ef; 
        10'b0100100001: data <= 18'h0045b; 
        10'b0100100010: data <= 18'h0042a; 
        10'b0100100011: data <= 18'h0050a; 
        10'b0100100100: data <= 18'h00430; 
        10'b0100100101: data <= 18'h00338; 
        10'b0100100110: data <= 18'h3ff4f; 
        10'b0100100111: data <= 18'h3fd5e; 
        10'b0100101000: data <= 18'h3fb9c; 
        10'b0100101001: data <= 18'h3fbbf; 
        10'b0100101010: data <= 18'h3fb99; 
        10'b0100101011: data <= 18'h3fafb; 
        10'b0100101100: data <= 18'h3fc90; 
        10'b0100101101: data <= 18'h3feef; 
        10'b0100101110: data <= 18'h00095; 
        10'b0100101111: data <= 18'h00338; 
        10'b0100110000: data <= 18'h0066d; 
        10'b0100110001: data <= 18'h004d5; 
        10'b0100110010: data <= 18'h001a5; 
        10'b0100110011: data <= 18'h3ff71; 
        10'b0100110100: data <= 18'h3ff3f; 
        10'b0100110101: data <= 18'h00001; 
        10'b0100110110: data <= 18'h3ff63; 
        10'b0100110111: data <= 18'h3ff99; 
        10'b0100111000: data <= 18'h3ff61; 
        10'b0100111001: data <= 18'h3ffe9; 
        10'b0100111010: data <= 18'h00226; 
        10'b0100111011: data <= 18'h002a0; 
        10'b0100111100: data <= 18'h003cb; 
        10'b0100111101: data <= 18'h00381; 
        10'b0100111110: data <= 18'h00291; 
        10'b0100111111: data <= 18'h002d4; 
        10'b0101000000: data <= 18'h004ad; 
        10'b0101000001: data <= 18'h0045e; 
        10'b0101000010: data <= 18'h00012; 
        10'b0101000011: data <= 18'h3fd47; 
        10'b0101000100: data <= 18'h3fca0; 
        10'b0101000101: data <= 18'h3fc5e; 
        10'b0101000110: data <= 18'h3fb26; 
        10'b0101000111: data <= 18'h3f93c; 
        10'b0101001000: data <= 18'h3f62d; 
        10'b0101001001: data <= 18'h3f6fb; 
        10'b0101001010: data <= 18'h3f89c; 
        10'b0101001011: data <= 18'h3fa9c; 
        10'b0101001100: data <= 18'h3fe15; 
        10'b0101001101: data <= 18'h00036; 
        10'b0101001110: data <= 18'h0008a; 
        10'b0101001111: data <= 18'h3ffac; 
        10'b0101010000: data <= 18'h3ffaa; 
        10'b0101010001: data <= 18'h3ffb9; 
        10'b0101010010: data <= 18'h3ff98; 
        10'b0101010011: data <= 18'h3ff6f; 
        10'b0101010100: data <= 18'h3ff92; 
        10'b0101010101: data <= 18'h00117; 
        10'b0101010110: data <= 18'h00278; 
        10'b0101010111: data <= 18'h00234; 
        10'b0101011000: data <= 18'h0019e; 
        10'b0101011001: data <= 18'h000ed; 
        10'b0101011010: data <= 18'h002bc; 
        10'b0101011011: data <= 18'h005a9; 
        10'b0101011100: data <= 18'h00549; 
        10'b0101011101: data <= 18'h0056b; 
        10'b0101011110: data <= 18'h0008f; 
        10'b0101011111: data <= 18'h3fd40; 
        10'b0101100000: data <= 18'h3fae4; 
        10'b0101100001: data <= 18'h3fbdd; 
        10'b0101100010: data <= 18'h3fd31; 
        10'b0101100011: data <= 18'h3fbf8; 
        10'b0101100100: data <= 18'h3fb68; 
        10'b0101100101: data <= 18'h3f861; 
        10'b0101100110: data <= 18'h3f74e; 
        10'b0101100111: data <= 18'h3f872; 
        10'b0101101000: data <= 18'h3faf3; 
        10'b0101101001: data <= 18'h3fe91; 
        10'b0101101010: data <= 18'h00013; 
        10'b0101101011: data <= 18'h3ffff; 
        10'b0101101100: data <= 18'h3ffb3; 
        10'b0101101101: data <= 18'h3ff49; 
        10'b0101101110: data <= 18'h3ff3d; 
        10'b0101101111: data <= 18'h3ff78; 
        10'b0101110000: data <= 18'h3ffd7; 
        10'b0101110001: data <= 18'h00092; 
        10'b0101110010: data <= 18'h001a7; 
        10'b0101110011: data <= 18'h00136; 
        10'b0101110100: data <= 18'h00167; 
        10'b0101110101: data <= 18'h00128; 
        10'b0101110110: data <= 18'h003ce; 
        10'b0101110111: data <= 18'h00441; 
        10'b0101111000: data <= 18'h0032a; 
        10'b0101111001: data <= 18'h002f5; 
        10'b0101111010: data <= 18'h3ff68; 
        10'b0101111011: data <= 18'h3fcba; 
        10'b0101111100: data <= 18'h3faad; 
        10'b0101111101: data <= 18'h3fd30; 
        10'b0101111110: data <= 18'h3ff00; 
        10'b0101111111: data <= 18'h3fed8; 
        10'b0110000000: data <= 18'h3ff73; 
        10'b0110000001: data <= 18'h3fdd7; 
        10'b0110000010: data <= 18'h3fc19; 
        10'b0110000011: data <= 18'h3fa4c; 
        10'b0110000100: data <= 18'h3fbb4; 
        10'b0110000101: data <= 18'h3ff41; 
        10'b0110000110: data <= 18'h3ff30; 
        10'b0110000111: data <= 18'h3ffe2; 
        10'b0110001000: data <= 18'h3ffb6; 
        10'b0110001001: data <= 18'h3ff3a; 
        10'b0110001010: data <= 18'h3ff9e; 
        10'b0110001011: data <= 18'h3ff0b; 
        10'b0110001100: data <= 18'h3ffae; 
        10'b0110001101: data <= 18'h3ffa7; 
        10'b0110001110: data <= 18'h3fffb; 
        10'b0110001111: data <= 18'h3ffd1; 
        10'b0110010000: data <= 18'h001c0; 
        10'b0110010001: data <= 18'h002c5; 
        10'b0110010010: data <= 18'h00352; 
        10'b0110010011: data <= 18'h000a3; 
        10'b0110010100: data <= 18'h00120; 
        10'b0110010101: data <= 18'h3ffcb; 
        10'b0110010110: data <= 18'h3fda0; 
        10'b0110010111: data <= 18'h3fd44; 
        10'b0110011000: data <= 18'h3fc34; 
        10'b0110011001: data <= 18'h3fca5; 
        10'b0110011010: data <= 18'h3fcdb; 
        10'b0110011011: data <= 18'h3fe7c; 
        10'b0110011100: data <= 18'h3feb0; 
        10'b0110011101: data <= 18'h3fecf; 
        10'b0110011110: data <= 18'h3ff47; 
        10'b0110011111: data <= 18'h3fcde; 
        10'b0110100000: data <= 18'h3fde4; 
        10'b0110100001: data <= 18'h3fef1; 
        10'b0110100010: data <= 18'h3ffa0; 
        10'b0110100011: data <= 18'h3ff10; 
        10'b0110100100: data <= 18'h3ff29; 
        10'b0110100101: data <= 18'h00021; 
        10'b0110100110: data <= 18'h3ff19; 
        10'b0110100111: data <= 18'h3ffa1; 
        10'b0110101000: data <= 18'h3fea9; 
        10'b0110101001: data <= 18'h3fdfd; 
        10'b0110101010: data <= 18'h3fd2f; 
        10'b0110101011: data <= 18'h3fe22; 
        10'b0110101100: data <= 18'h000ae; 
        10'b0110101101: data <= 18'h0031e; 
        10'b0110101110: data <= 18'h0017b; 
        10'b0110101111: data <= 18'h0015d; 
        10'b0110110000: data <= 18'h0012d; 
        10'b0110110001: data <= 18'h3fef0; 
        10'b0110110010: data <= 18'h3fc79; 
        10'b0110110011: data <= 18'h3fbf2; 
        10'b0110110100: data <= 18'h3fc57; 
        10'b0110110101: data <= 18'h3fc40; 
        10'b0110110110: data <= 18'h3fd5c; 
        10'b0110110111: data <= 18'h3ffde; 
        10'b0110111000: data <= 18'h3ff1a; 
        10'b0110111001: data <= 18'h3ff3e; 
        10'b0110111010: data <= 18'h3ff18; 
        10'b0110111011: data <= 18'h3fef5; 
        10'b0110111100: data <= 18'h3ff45; 
        10'b0110111101: data <= 18'h3fffa; 
        10'b0110111110: data <= 18'h00025; 
        10'b0110111111: data <= 18'h3ff70; 
        10'b0111000000: data <= 18'h3ff7f; 
        10'b0111000001: data <= 18'h3ffac; 
        10'b0111000010: data <= 18'h3ffc8; 
        10'b0111000011: data <= 18'h3ff19; 
        10'b0111000100: data <= 18'h3ff7a; 
        10'b0111000101: data <= 18'h3fdb6; 
        10'b0111000110: data <= 18'h3fb6a; 
        10'b0111000111: data <= 18'h3fa93; 
        10'b0111001000: data <= 18'h3fc55; 
        10'b0111001001: data <= 18'h3fdf8; 
        10'b0111001010: data <= 18'h3ff32; 
        10'b0111001011: data <= 18'h3fed7; 
        10'b0111001100: data <= 18'h3ff3e; 
        10'b0111001101: data <= 18'h3fd80; 
        10'b0111001110: data <= 18'h3fb2f; 
        10'b0111001111: data <= 18'h3fc17; 
        10'b0111010000: data <= 18'h3fd29; 
        10'b0111010001: data <= 18'h3fefa; 
        10'b0111010010: data <= 18'h3ff09; 
        10'b0111010011: data <= 18'h00028; 
        10'b0111010100: data <= 18'h000cb; 
        10'b0111010101: data <= 18'h00020; 
        10'b0111010110: data <= 18'h000dc; 
        10'b0111010111: data <= 18'h00032; 
        10'b0111011000: data <= 18'h00022; 
        10'b0111011001: data <= 18'h0001f; 
        10'b0111011010: data <= 18'h3ff76; 
        10'b0111011011: data <= 18'h3ff81; 
        10'b0111011100: data <= 18'h3ff67; 
        10'b0111011101: data <= 18'h3fff6; 
        10'b0111011110: data <= 18'h3ffff; 
        10'b0111011111: data <= 18'h00011; 
        10'b0111100000: data <= 18'h3ff6b; 
        10'b0111100001: data <= 18'h0002b; 
        10'b0111100010: data <= 18'h00056; 
        10'b0111100011: data <= 18'h3fc6b; 
        10'b0111100100: data <= 18'h3f985; 
        10'b0111100101: data <= 18'h3f9ef; 
        10'b0111100110: data <= 18'h3fba8; 
        10'b0111100111: data <= 18'h3fd63; 
        10'b0111101000: data <= 18'h3fbea; 
        10'b0111101001: data <= 18'h3faba; 
        10'b0111101010: data <= 18'h3fadf; 
        10'b0111101011: data <= 18'h3fdaa; 
        10'b0111101100: data <= 18'h3fef9; 
        10'b0111101101: data <= 18'h0018d; 
        10'b0111101110: data <= 18'h0025f; 
        10'b0111101111: data <= 18'h0018c; 
        10'b0111110000: data <= 18'h00190; 
        10'b0111110001: data <= 18'h00074; 
        10'b0111110010: data <= 18'h0000d; 
        10'b0111110011: data <= 18'h000dd; 
        10'b0111110100: data <= 18'h000e0; 
        10'b0111110101: data <= 18'h3ff43; 
        10'b0111110110: data <= 18'h3fff8; 
        10'b0111110111: data <= 18'h00005; 
        10'b0111111000: data <= 18'h00016; 
        10'b0111111001: data <= 18'h3ff5f; 
        10'b0111111010: data <= 18'h3ff9a; 
        10'b0111111011: data <= 18'h3ff7d; 
        10'b0111111100: data <= 18'h00148; 
        10'b0111111101: data <= 18'h001b2; 
        10'b0111111110: data <= 18'h00407; 
        10'b0111111111: data <= 18'h000b5; 
        10'b1000000000: data <= 18'h3fc20; 
        10'b1000000001: data <= 18'h3fa5c; 
        10'b1000000010: data <= 18'h3f893; 
        10'b1000000011: data <= 18'h3f95f; 
        10'b1000000100: data <= 18'h3fb3f; 
        10'b1000000101: data <= 18'h3fd49; 
        10'b1000000110: data <= 18'h3fea5; 
        10'b1000000111: data <= 18'h3ff6f; 
        10'b1000001000: data <= 18'h3ffe6; 
        10'b1000001001: data <= 18'h001d2; 
        10'b1000001010: data <= 18'h000ea; 
        10'b1000001011: data <= 18'h001a0; 
        10'b1000001100: data <= 18'h00117; 
        10'b1000001101: data <= 18'h00195; 
        10'b1000001110: data <= 18'h0014e; 
        10'b1000001111: data <= 18'h001ce; 
        10'b1000010000: data <= 18'h000f0; 
        10'b1000010001: data <= 18'h00012; 
        10'b1000010010: data <= 18'h3ff50; 
        10'b1000010011: data <= 18'h3ffc8; 
        10'b1000010100: data <= 18'h00001; 
        10'b1000010101: data <= 18'h3ff5e; 
        10'b1000010110: data <= 18'h3ffa9; 
        10'b1000010111: data <= 18'h00023; 
        10'b1000011000: data <= 18'h001f2; 
        10'b1000011001: data <= 18'h00353; 
        10'b1000011010: data <= 18'h0047a; 
        10'b1000011011: data <= 18'h00304; 
        10'b1000011100: data <= 18'h001e9; 
        10'b1000011101: data <= 18'h0009f; 
        10'b1000011110: data <= 18'h3fe93; 
        10'b1000011111: data <= 18'h3fe7a; 
        10'b1000100000: data <= 18'h00021; 
        10'b1000100001: data <= 18'h001d3; 
        10'b1000100010: data <= 18'h000af; 
        10'b1000100011: data <= 18'h000f8; 
        10'b1000100100: data <= 18'h000fc; 
        10'b1000100101: data <= 18'h3ffb1; 
        10'b1000100110: data <= 18'h000b5; 
        10'b1000100111: data <= 18'h000b1; 
        10'b1000101000: data <= 18'h00026; 
        10'b1000101001: data <= 18'h0012f; 
        10'b1000101010: data <= 18'h00208; 
        10'b1000101011: data <= 18'h0017c; 
        10'b1000101100: data <= 18'h00020; 
        10'b1000101101: data <= 18'h3fffa; 
        10'b1000101110: data <= 18'h3fffe; 
        10'b1000101111: data <= 18'h3ff34; 
        10'b1000110000: data <= 18'h3fff6; 
        10'b1000110001: data <= 18'h3ff12; 
        10'b1000110010: data <= 18'h3ff8e; 
        10'b1000110011: data <= 18'h3ff4e; 
        10'b1000110100: data <= 18'h00043; 
        10'b1000110101: data <= 18'h00230; 
        10'b1000110110: data <= 18'h0028a; 
        10'b1000110111: data <= 18'h00318; 
        10'b1000111000: data <= 18'h00456; 
        10'b1000111001: data <= 18'h003a9; 
        10'b1000111010: data <= 18'h00338; 
        10'b1000111011: data <= 18'h004b0; 
        10'b1000111100: data <= 18'h002eb; 
        10'b1000111101: data <= 18'h00230; 
        10'b1000111110: data <= 18'h3ff62; 
        10'b1000111111: data <= 18'h3ff6f; 
        10'b1001000000: data <= 18'h0019d; 
        10'b1001000001: data <= 18'h000d3; 
        10'b1001000010: data <= 18'h00159; 
        10'b1001000011: data <= 18'h001c9; 
        10'b1001000100: data <= 18'h00190; 
        10'b1001000101: data <= 18'h0013a; 
        10'b1001000110: data <= 18'h002ef; 
        10'b1001000111: data <= 18'h00231; 
        10'b1001001000: data <= 18'h3ffb7; 
        10'b1001001001: data <= 18'h3ff16; 
        10'b1001001010: data <= 18'h3ffae; 
        10'b1001001011: data <= 18'h3ff6c; 
        10'b1001001100: data <= 18'h3ff56; 
        10'b1001001101: data <= 18'h00005; 
        10'b1001001110: data <= 18'h3ff08; 
        10'b1001001111: data <= 18'h3ffa3; 
        10'b1001010000: data <= 18'h000dd; 
        10'b1001010001: data <= 18'h3ffb9; 
        10'b1001010010: data <= 18'h0010c; 
        10'b1001010011: data <= 18'h002d5; 
        10'b1001010100: data <= 18'h00416; 
        10'b1001010101: data <= 18'h002ac; 
        10'b1001010110: data <= 18'h00244; 
        10'b1001010111: data <= 18'h00139; 
        10'b1001011000: data <= 18'h00195; 
        10'b1001011001: data <= 18'h000fc; 
        10'b1001011010: data <= 18'h00106; 
        10'b1001011011: data <= 18'h0013f; 
        10'b1001011100: data <= 18'h00053; 
        10'b1001011101: data <= 18'h00101; 
        10'b1001011110: data <= 18'h00084; 
        10'b1001011111: data <= 18'h0019f; 
        10'b1001100000: data <= 18'h00197; 
        10'b1001100001: data <= 18'h002ab; 
        10'b1001100010: data <= 18'h00348; 
        10'b1001100011: data <= 18'h000b6; 
        10'b1001100100: data <= 18'h00007; 
        10'b1001100101: data <= 18'h3ff38; 
        10'b1001100110: data <= 18'h3ff6e; 
        10'b1001100111: data <= 18'h3ff6f; 
        10'b1001101000: data <= 18'h3ffcf; 
        10'b1001101001: data <= 18'h3ff1d; 
        10'b1001101010: data <= 18'h3ff8a; 
        10'b1001101011: data <= 18'h3ff6e; 
        10'b1001101100: data <= 18'h00050; 
        10'b1001101101: data <= 18'h3ff90; 
        10'b1001101110: data <= 18'h3ff0b; 
        10'b1001101111: data <= 18'h3ffd4; 
        10'b1001110000: data <= 18'h00197; 
        10'b1001110001: data <= 18'h00252; 
        10'b1001110010: data <= 18'h00067; 
        10'b1001110011: data <= 18'h0020e; 
        10'b1001110100: data <= 18'h00353; 
        10'b1001110101: data <= 18'h0041b; 
        10'b1001110110: data <= 18'h00217; 
        10'b1001110111: data <= 18'h00051; 
        10'b1001111000: data <= 18'h0003b; 
        10'b1001111001: data <= 18'h00083; 
        10'b1001111010: data <= 18'h00113; 
        10'b1001111011: data <= 18'h00112; 
        10'b1001111100: data <= 18'h001d5; 
        10'b1001111101: data <= 18'h001a8; 
        10'b1001111110: data <= 18'h001bb; 
        10'b1001111111: data <= 18'h0009c; 
        10'b1010000000: data <= 18'h3ffe9; 
        10'b1010000001: data <= 18'h00019; 
        10'b1010000010: data <= 18'h3ffaa; 
        10'b1010000011: data <= 18'h3ffc7; 
        10'b1010000100: data <= 18'h3ff45; 
        10'b1010000101: data <= 18'h3ffa5; 
        10'b1010000110: data <= 18'h3ffcb; 
        10'b1010000111: data <= 18'h3ffb7; 
        10'b1010001000: data <= 18'h3ff4e; 
        10'b1010001001: data <= 18'h3ff8b; 
        10'b1010001010: data <= 18'h3fe9c; 
        10'b1010001011: data <= 18'h3ff5e; 
        10'b1010001100: data <= 18'h00142; 
        10'b1010001101: data <= 18'h0013b; 
        10'b1010001110: data <= 18'h0013b; 
        10'b1010001111: data <= 18'h00231; 
        10'b1010010000: data <= 18'h0021a; 
        10'b1010010001: data <= 18'h00171; 
        10'b1010010010: data <= 18'h001a8; 
        10'b1010010011: data <= 18'h00184; 
        10'b1010010100: data <= 18'h0017b; 
        10'b1010010101: data <= 18'h000af; 
        10'b1010010110: data <= 18'h3ff38; 
        10'b1010010111: data <= 18'h3ffe4; 
        10'b1010011000: data <= 18'h000ba; 
        10'b1010011001: data <= 18'h0004b; 
        10'b1010011010: data <= 18'h000f9; 
        10'b1010011011: data <= 18'h3ff64; 
        10'b1010011100: data <= 18'h0002a; 
        10'b1010011101: data <= 18'h3ff80; 
        10'b1010011110: data <= 18'h3ff7e; 
        10'b1010011111: data <= 18'h00027; 
        10'b1010100000: data <= 18'h3ffee; 
        10'b1010100001: data <= 18'h3ff85; 
        10'b1010100010: data <= 18'h3ff73; 
        10'b1010100011: data <= 18'h0002c; 
        10'b1010100100: data <= 18'h3ff0c; 
        10'b1010100101: data <= 18'h3fefd; 
        10'b1010100110: data <= 18'h3ffa3; 
        10'b1010100111: data <= 18'h3ffd1; 
        10'b1010101000: data <= 18'h3fff1; 
        10'b1010101001: data <= 18'h001a1; 
        10'b1010101010: data <= 18'h0021d; 
        10'b1010101011: data <= 18'h001a0; 
        10'b1010101100: data <= 18'h0010e; 
        10'b1010101101: data <= 18'h00178; 
        10'b1010101110: data <= 18'h002b6; 
        10'b1010101111: data <= 18'h0023e; 
        10'b1010110000: data <= 18'h00157; 
        10'b1010110001: data <= 18'h000a7; 
        10'b1010110010: data <= 18'h0013e; 
        10'b1010110011: data <= 18'h000ce; 
        10'b1010110100: data <= 18'h3fff4; 
        10'b1010110101: data <= 18'h3ffe2; 
        10'b1010110110: data <= 18'h3ffb5; 
        10'b1010110111: data <= 18'h0000d; 
        10'b1010111000: data <= 18'h3ff58; 
        10'b1010111001: data <= 18'h3ffc4; 
        10'b1010111010: data <= 18'h00019; 
        10'b1010111011: data <= 18'h3ff33; 
        10'b1010111100: data <= 18'h3ffa4; 
        10'b1010111101: data <= 18'h00009; 
        10'b1010111110: data <= 18'h00018; 
        10'b1010111111: data <= 18'h3ff29; 
        10'b1011000000: data <= 18'h3fffe; 
        10'b1011000001: data <= 18'h3ffbd; 
        10'b1011000010: data <= 18'h3ff00; 
        10'b1011000011: data <= 18'h3ffa2; 
        10'b1011000100: data <= 18'h3ff1b; 
        10'b1011000101: data <= 18'h00087; 
        10'b1011000110: data <= 18'h00065; 
        10'b1011000111: data <= 18'h0011a; 
        10'b1011001000: data <= 18'h00118; 
        10'b1011001001: data <= 18'h001eb; 
        10'b1011001010: data <= 18'h0001b; 
        10'b1011001011: data <= 18'h00092; 
        10'b1011001100: data <= 18'h0007c; 
        10'b1011001101: data <= 18'h000f1; 
        10'b1011001110: data <= 18'h3ff5f; 
        10'b1011001111: data <= 18'h3fff9; 
        10'b1011010000: data <= 18'h3fef4; 
        10'b1011010001: data <= 18'h00017; 
        10'b1011010010: data <= 18'h3ff9c; 
        10'b1011010011: data <= 18'h3ff4c; 
        10'b1011010100: data <= 18'h3ffeb; 
        10'b1011010101: data <= 18'h0000c; 
        10'b1011010110: data <= 18'h3ff1b; 
        10'b1011010111: data <= 18'h3ff87; 
        10'b1011011000: data <= 18'h3ffb8; 
        10'b1011011001: data <= 18'h3ffb1; 
        10'b1011011010: data <= 18'h3ff58; 
        10'b1011011011: data <= 18'h3ff81; 
        10'b1011011100: data <= 18'h3ff72; 
        10'b1011011101: data <= 18'h3ff8c; 
        10'b1011011110: data <= 18'h3ffd6; 
        10'b1011011111: data <= 18'h3ff59; 
        10'b1011100000: data <= 18'h3ff24; 
        10'b1011100001: data <= 18'h3ff8e; 
        10'b1011100010: data <= 18'h3ff6a; 
        10'b1011100011: data <= 18'h3ffe4; 
        10'b1011100100: data <= 18'h00004; 
        10'b1011100101: data <= 18'h3ffc6; 
        10'b1011100110: data <= 18'h3ff60; 
        10'b1011100111: data <= 18'h3ffae; 
        10'b1011101000: data <= 18'h3ffdb; 
        10'b1011101001: data <= 18'h3ff58; 
        10'b1011101010: data <= 18'h3febd; 
        10'b1011101011: data <= 18'h3fefa; 
        10'b1011101100: data <= 18'h3ffc9; 
        10'b1011101101: data <= 18'h3ffc7; 
        10'b1011101110: data <= 18'h3ff6c; 
        10'b1011101111: data <= 18'h3ffd5; 
        10'b1011110000: data <= 18'h3ff92; 
        10'b1011110001: data <= 18'h3ffb5; 
        10'b1011110010: data <= 18'h3ff78; 
        10'b1011110011: data <= 18'h3ff1b; 
        10'b1011110100: data <= 18'h3ffce; 
        10'b1011110101: data <= 18'h3ffe1; 
        10'b1011110110: data <= 18'h3ffea; 
        10'b1011110111: data <= 18'h3ffc0; 
        10'b1011111000: data <= 18'h3ff3d; 
        10'b1011111001: data <= 18'h3fff4; 
        10'b1011111010: data <= 18'h3ff7c; 
        10'b1011111011: data <= 18'h3ff70; 
        10'b1011111100: data <= 18'h0002f; 
        10'b1011111101: data <= 18'h3ff76; 
        10'b1011111110: data <= 18'h3ff63; 
        10'b1011111111: data <= 18'h3ffed; 
        10'b1100000000: data <= 18'h3ffac; 
        10'b1100000001: data <= 18'h3ff10; 
        10'b1100000010: data <= 18'h00005; 
        10'b1100000011: data <= 18'h3ffb6; 
        10'b1100000100: data <= 18'h3ff26; 
        10'b1100000101: data <= 18'h3ff0f; 
        10'b1100000110: data <= 18'h3ff4c; 
        10'b1100000111: data <= 18'h3ff0b; 
        10'b1100001000: data <= 18'h3fffc; 
        10'b1100001001: data <= 18'h3ff79; 
        10'b1100001010: data <= 18'h0002d; 
        10'b1100001011: data <= 18'h3ff30; 
        10'b1100001100: data <= 18'h3ffc1; 
        10'b1100001101: data <= 18'h3ff97; 
        10'b1100001110: data <= 18'h3ff3f; 
        10'b1100001111: data <= 18'h3ffe2; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 13) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 19'h7fee4; 
        10'b0000000001: data <= 19'h7ffd8; 
        10'b0000000010: data <= 19'h7ffd7; 
        10'b0000000011: data <= 19'h7fe82; 
        10'b0000000100: data <= 19'h7ff4c; 
        10'b0000000101: data <= 19'h7ff1c; 
        10'b0000000110: data <= 19'h7ffff; 
        10'b0000000111: data <= 19'h7ff0b; 
        10'b0000001000: data <= 19'h7ff9b; 
        10'b0000001001: data <= 19'h00052; 
        10'b0000001010: data <= 19'h7ff9b; 
        10'b0000001011: data <= 19'h7ff91; 
        10'b0000001100: data <= 19'h7fedd; 
        10'b0000001101: data <= 19'h7ffee; 
        10'b0000001110: data <= 19'h7fe7c; 
        10'b0000001111: data <= 19'h7fec0; 
        10'b0000010000: data <= 19'h7fe48; 
        10'b0000010001: data <= 19'h7fe9b; 
        10'b0000010010: data <= 19'h7ffcc; 
        10'b0000010011: data <= 19'h7ff9e; 
        10'b0000010100: data <= 19'h7fe43; 
        10'b0000010101: data <= 19'h7ff57; 
        10'b0000010110: data <= 19'h7ff85; 
        10'b0000010111: data <= 19'h7ff25; 
        10'b0000011000: data <= 19'h7fe5d; 
        10'b0000011001: data <= 19'h7ff62; 
        10'b0000011010: data <= 19'h7ff85; 
        10'b0000011011: data <= 19'h7fef0; 
        10'b0000011100: data <= 19'h7ffe6; 
        10'b0000011101: data <= 19'h7fe2d; 
        10'b0000011110: data <= 19'h7fffd; 
        10'b0000011111: data <= 19'h7fe70; 
        10'b0000100000: data <= 19'h7ffef; 
        10'b0000100001: data <= 19'h7feff; 
        10'b0000100010: data <= 19'h7ff7c; 
        10'b0000100011: data <= 19'h7fef5; 
        10'b0000100100: data <= 19'h7feb1; 
        10'b0000100101: data <= 19'h7ff86; 
        10'b0000100110: data <= 19'h00029; 
        10'b0000100111: data <= 19'h7fe7a; 
        10'b0000101000: data <= 19'h7fef1; 
        10'b0000101001: data <= 19'h7fea5; 
        10'b0000101010: data <= 19'h7fe40; 
        10'b0000101011: data <= 19'h7ffb5; 
        10'b0000101100: data <= 19'h7fed1; 
        10'b0000101101: data <= 19'h7fe9e; 
        10'b0000101110: data <= 19'h7feda; 
        10'b0000101111: data <= 19'h7fec6; 
        10'b0000110000: data <= 19'h7ff9d; 
        10'b0000110001: data <= 19'h7fe69; 
        10'b0000110010: data <= 19'h7fffa; 
        10'b0000110011: data <= 19'h7fe85; 
        10'b0000110100: data <= 19'h00005; 
        10'b0000110101: data <= 19'h7ffe1; 
        10'b0000110110: data <= 19'h7fe95; 
        10'b0000110111: data <= 19'h7ff37; 
        10'b0000111000: data <= 19'h7ff3c; 
        10'b0000111001: data <= 19'h7ffaa; 
        10'b0000111010: data <= 19'h7fef3; 
        10'b0000111011: data <= 19'h7fe43; 
        10'b0000111100: data <= 19'h7fe92; 
        10'b0000111101: data <= 19'h7ff65; 
        10'b0000111110: data <= 19'h7fff1; 
        10'b0000111111: data <= 19'h7ff87; 
        10'b0001000000: data <= 19'h7febe; 
        10'b0001000001: data <= 19'h7ff09; 
        10'b0001000010: data <= 19'h0003d; 
        10'b0001000011: data <= 19'h7fe27; 
        10'b0001000100: data <= 19'h7ffea; 
        10'b0001000101: data <= 19'h7feb3; 
        10'b0001000110: data <= 19'h7fe4e; 
        10'b0001000111: data <= 19'h7fe9f; 
        10'b0001001000: data <= 19'h7fee5; 
        10'b0001001001: data <= 19'h7ff5c; 
        10'b0001001010: data <= 19'h7ff0a; 
        10'b0001001011: data <= 19'h7ff0d; 
        10'b0001001100: data <= 19'h0006d; 
        10'b0001001101: data <= 19'h0000c; 
        10'b0001001110: data <= 19'h0002e; 
        10'b0001001111: data <= 19'h7fea9; 
        10'b0001010000: data <= 19'h7fe42; 
        10'b0001010001: data <= 19'h7ff22; 
        10'b0001010010: data <= 19'h7ffe5; 
        10'b0001010011: data <= 19'h7ff86; 
        10'b0001010100: data <= 19'h7ffac; 
        10'b0001010101: data <= 19'h7ff7f; 
        10'b0001010110: data <= 19'h7fe96; 
        10'b0001010111: data <= 19'h7ffe9; 
        10'b0001011000: data <= 19'h7fe71; 
        10'b0001011001: data <= 19'h7fef8; 
        10'b0001011010: data <= 19'h7fe26; 
        10'b0001011011: data <= 19'h7fecb; 
        10'b0001011100: data <= 19'h7fe48; 
        10'b0001011101: data <= 19'h7fec5; 
        10'b0001011110: data <= 19'h7fd02; 
        10'b0001011111: data <= 19'h7fc2e; 
        10'b0001100000: data <= 19'h7fdd2; 
        10'b0001100001: data <= 19'h7fdf4; 
        10'b0001100010: data <= 19'h7fd7d; 
        10'b0001100011: data <= 19'h7ff2b; 
        10'b0001100100: data <= 19'h7ffa4; 
        10'b0001100101: data <= 19'h7fe07; 
        10'b0001100110: data <= 19'h7fed1; 
        10'b0001100111: data <= 19'h7ffa1; 
        10'b0001101000: data <= 19'h7ffbb; 
        10'b0001101001: data <= 19'h7ff2e; 
        10'b0001101010: data <= 19'h7fdff; 
        10'b0001101011: data <= 19'h7fea8; 
        10'b0001101100: data <= 19'h7fd96; 
        10'b0001101101: data <= 19'h00047; 
        10'b0001101110: data <= 19'h0002c; 
        10'b0001101111: data <= 19'h7fe6c; 
        10'b0001110000: data <= 19'h7fe51; 
        10'b0001110001: data <= 19'h7fef5; 
        10'b0001110010: data <= 19'h0002c; 
        10'b0001110011: data <= 19'h00018; 
        10'b0001110100: data <= 19'h0003c; 
        10'b0001110101: data <= 19'h7fecb; 
        10'b0001110110: data <= 19'h7feb3; 
        10'b0001110111: data <= 19'h7fd4d; 
        10'b0001111000: data <= 19'h7fb72; 
        10'b0001111001: data <= 19'h7f9f3; 
        10'b0001111010: data <= 19'h7f72b; 
        10'b0001111011: data <= 19'h7fa5b; 
        10'b0001111100: data <= 19'h7fa50; 
        10'b0001111101: data <= 19'h7f85f; 
        10'b0001111110: data <= 19'h7fbcc; 
        10'b0001111111: data <= 19'h7fffb; 
        10'b0010000000: data <= 19'h7ff80; 
        10'b0010000001: data <= 19'h0016c; 
        10'b0010000010: data <= 19'h7ff91; 
        10'b0010000011: data <= 19'h7fdd5; 
        10'b0010000100: data <= 19'h7fd2b; 
        10'b0010000101: data <= 19'h7fe80; 
        10'b0010000110: data <= 19'h7fec6; 
        10'b0010000111: data <= 19'h7ff24; 
        10'b0010001000: data <= 19'h7feef; 
        10'b0010001001: data <= 19'h00066; 
        10'b0010001010: data <= 19'h0003a; 
        10'b0010001011: data <= 19'h7ff38; 
        10'b0010001100: data <= 19'h7ff5c; 
        10'b0010001101: data <= 19'h00065; 
        10'b0010001110: data <= 19'h7fea2; 
        10'b0010001111: data <= 19'h7fe6e; 
        10'b0010010000: data <= 19'h7fed7; 
        10'b0010010001: data <= 19'h7fd3e; 
        10'b0010010010: data <= 19'h7fbd5; 
        10'b0010010011: data <= 19'h7fbf9; 
        10'b0010010100: data <= 19'h7fd5c; 
        10'b0010010101: data <= 19'h7ff82; 
        10'b0010010110: data <= 19'h000e4; 
        10'b0010010111: data <= 19'h000f6; 
        10'b0010011000: data <= 19'h7fe92; 
        10'b0010011001: data <= 19'h7fdf5; 
        10'b0010011010: data <= 19'h7fec4; 
        10'b0010011011: data <= 19'h7ff6c; 
        10'b0010011100: data <= 19'h0020b; 
        10'b0010011101: data <= 19'h00216; 
        10'b0010011110: data <= 19'h003f5; 
        10'b0010011111: data <= 19'h00277; 
        10'b0010100000: data <= 19'h00264; 
        10'b0010100001: data <= 19'h00312; 
        10'b0010100010: data <= 19'h005aa; 
        10'b0010100011: data <= 19'h004d1; 
        10'b0010100100: data <= 19'h00361; 
        10'b0010100101: data <= 19'h001de; 
        10'b0010100110: data <= 19'h0012a; 
        10'b0010100111: data <= 19'h0006f; 
        10'b0010101000: data <= 19'h7fe7f; 
        10'b0010101001: data <= 19'h7fe5c; 
        10'b0010101010: data <= 19'h00035; 
        10'b0010101011: data <= 19'h7fe6b; 
        10'b0010101100: data <= 19'h7fdf7; 
        10'b0010101101: data <= 19'h7fb23; 
        10'b0010101110: data <= 19'h7fdd0; 
        10'b0010101111: data <= 19'h7ffbe; 
        10'b0010110000: data <= 19'h7ffd4; 
        10'b0010110001: data <= 19'h001f9; 
        10'b0010110010: data <= 19'h00419; 
        10'b0010110011: data <= 19'h00369; 
        10'b0010110100: data <= 19'h00094; 
        10'b0010110101: data <= 19'h00141; 
        10'b0010110110: data <= 19'h7ff70; 
        10'b0010110111: data <= 19'h7fe0f; 
        10'b0010111000: data <= 19'h7fed3; 
        10'b0010111001: data <= 19'h7ff02; 
        10'b0010111010: data <= 19'h0000b; 
        10'b0010111011: data <= 19'h003e4; 
        10'b0010111100: data <= 19'h0023a; 
        10'b0010111101: data <= 19'h00288; 
        10'b0010111110: data <= 19'h007bb; 
        10'b0010111111: data <= 19'h0094c; 
        10'b0011000000: data <= 19'h00a75; 
        10'b0011000001: data <= 19'h00588; 
        10'b0011000010: data <= 19'h002bb; 
        10'b0011000011: data <= 19'h000ab; 
        10'b0011000100: data <= 19'h7ff25; 
        10'b0011000101: data <= 19'h7ff8a; 
        10'b0011000110: data <= 19'h7ff55; 
        10'b0011000111: data <= 19'h7fdff; 
        10'b0011001000: data <= 19'h7fa59; 
        10'b0011001001: data <= 19'h7f95d; 
        10'b0011001010: data <= 19'h7fbf6; 
        10'b0011001011: data <= 19'h00086; 
        10'b0011001100: data <= 19'h002a5; 
        10'b0011001101: data <= 19'h00532; 
        10'b0011001110: data <= 19'h0050e; 
        10'b0011001111: data <= 19'h0046a; 
        10'b0011010000: data <= 19'h00147; 
        10'b0011010001: data <= 19'h7ff95; 
        10'b0011010010: data <= 19'h7fe97; 
        10'b0011010011: data <= 19'h00019; 
        10'b0011010100: data <= 19'h00230; 
        10'b0011010101: data <= 19'h001fb; 
        10'b0011010110: data <= 19'h00281; 
        10'b0011010111: data <= 19'h0059a; 
        10'b0011011000: data <= 19'h004d7; 
        10'b0011011001: data <= 19'h005ca; 
        10'b0011011010: data <= 19'h00818; 
        10'b0011011011: data <= 19'h00adc; 
        10'b0011011100: data <= 19'h00d42; 
        10'b0011011101: data <= 19'h00992; 
        10'b0011011110: data <= 19'h00179; 
        10'b0011011111: data <= 19'h7ffc6; 
        10'b0011100000: data <= 19'h7ff9f; 
        10'b0011100001: data <= 19'h00059; 
        10'b0011100010: data <= 19'h7fff8; 
        10'b0011100011: data <= 19'h7fd45; 
        10'b0011100100: data <= 19'h7f7dc; 
        10'b0011100101: data <= 19'h7f90a; 
        10'b0011100110: data <= 19'h7faf6; 
        10'b0011100111: data <= 19'h00050; 
        10'b0011101000: data <= 19'h003f0; 
        10'b0011101001: data <= 19'h00128; 
        10'b0011101010: data <= 19'h0021e; 
        10'b0011101011: data <= 19'h0041c; 
        10'b0011101100: data <= 19'h00281; 
        10'b0011101101: data <= 19'h7fd2f; 
        10'b0011101110: data <= 19'h7f9d2; 
        10'b0011101111: data <= 19'h7fc42; 
        10'b0011110000: data <= 19'h7fdb4; 
        10'b0011110001: data <= 19'h00038; 
        10'b0011110010: data <= 19'h000a1; 
        10'b0011110011: data <= 19'h004ab; 
        10'b0011110100: data <= 19'h004ed; 
        10'b0011110101: data <= 19'h00705; 
        10'b0011110110: data <= 19'h00b17; 
        10'b0011110111: data <= 19'h00e83; 
        10'b0011111000: data <= 19'h0135d; 
        10'b0011111001: data <= 19'h00c82; 
        10'b0011111010: data <= 19'h00247; 
        10'b0011111011: data <= 19'h7ffc4; 
        10'b0011111100: data <= 19'h7fe66; 
        10'b0011111101: data <= 19'h7ff10; 
        10'b0011111110: data <= 19'h7fe40; 
        10'b0011111111: data <= 19'h7fc33; 
        10'b0100000000: data <= 19'h7fba2; 
        10'b0100000001: data <= 19'h7fbf7; 
        10'b0100000010: data <= 19'h0007e; 
        10'b0100000011: data <= 19'h7ffb8; 
        10'b0100000100: data <= 19'h0035c; 
        10'b0100000101: data <= 19'h002eb; 
        10'b0100000110: data <= 19'h0032d; 
        10'b0100000111: data <= 19'h0087a; 
        10'b0100001000: data <= 19'h00577; 
        10'b0100001001: data <= 19'h7fdbc; 
        10'b0100001010: data <= 19'h7f88d; 
        10'b0100001011: data <= 19'h7f552; 
        10'b0100001100: data <= 19'h7f606; 
        10'b0100001101: data <= 19'h7fa32; 
        10'b0100001110: data <= 19'h7feab; 
        10'b0100001111: data <= 19'h7fff7; 
        10'b0100010000: data <= 19'h00489; 
        10'b0100010001: data <= 19'h009b2; 
        10'b0100010010: data <= 19'h00e08; 
        10'b0100010011: data <= 19'h01331; 
        10'b0100010100: data <= 19'h0181f; 
        10'b0100010101: data <= 19'h00fd9; 
        10'b0100010110: data <= 19'h002d6; 
        10'b0100010111: data <= 19'h7fee2; 
        10'b0100011000: data <= 19'h7ffa8; 
        10'b0100011001: data <= 19'h7fee4; 
        10'b0100011010: data <= 19'h7fe81; 
        10'b0100011011: data <= 19'h7fecc; 
        10'b0100011100: data <= 19'h7feba; 
        10'b0100011101: data <= 19'h7ff2e; 
        10'b0100011110: data <= 19'h002b5; 
        10'b0100011111: data <= 19'h0050b; 
        10'b0100100000: data <= 19'h007df; 
        10'b0100100001: data <= 19'h008b6; 
        10'b0100100010: data <= 19'h00853; 
        10'b0100100011: data <= 19'h00a13; 
        10'b0100100100: data <= 19'h00861; 
        10'b0100100101: data <= 19'h00670; 
        10'b0100100110: data <= 19'h7fe9f; 
        10'b0100100111: data <= 19'h7fabd; 
        10'b0100101000: data <= 19'h7f737; 
        10'b0100101001: data <= 19'h7f77f; 
        10'b0100101010: data <= 19'h7f732; 
        10'b0100101011: data <= 19'h7f5f6; 
        10'b0100101100: data <= 19'h7f921; 
        10'b0100101101: data <= 19'h7fdde; 
        10'b0100101110: data <= 19'h0012b; 
        10'b0100101111: data <= 19'h00671; 
        10'b0100110000: data <= 19'h00cda; 
        10'b0100110001: data <= 19'h009a9; 
        10'b0100110010: data <= 19'h00349; 
        10'b0100110011: data <= 19'h7fee3; 
        10'b0100110100: data <= 19'h7fe7f; 
        10'b0100110101: data <= 19'h00003; 
        10'b0100110110: data <= 19'h7fec6; 
        10'b0100110111: data <= 19'h7ff32; 
        10'b0100111000: data <= 19'h7fec2; 
        10'b0100111001: data <= 19'h7ffd3; 
        10'b0100111010: data <= 19'h0044d; 
        10'b0100111011: data <= 19'h00540; 
        10'b0100111100: data <= 19'h00797; 
        10'b0100111101: data <= 19'h00703; 
        10'b0100111110: data <= 19'h00522; 
        10'b0100111111: data <= 19'h005a7; 
        10'b0101000000: data <= 19'h0095b; 
        10'b0101000001: data <= 19'h008bd; 
        10'b0101000010: data <= 19'h00024; 
        10'b0101000011: data <= 19'h7fa8f; 
        10'b0101000100: data <= 19'h7f941; 
        10'b0101000101: data <= 19'h7f8bc; 
        10'b0101000110: data <= 19'h7f64d; 
        10'b0101000111: data <= 19'h7f277; 
        10'b0101001000: data <= 19'h7ec5a; 
        10'b0101001001: data <= 19'h7edf6; 
        10'b0101001010: data <= 19'h7f138; 
        10'b0101001011: data <= 19'h7f538; 
        10'b0101001100: data <= 19'h7fc2a; 
        10'b0101001101: data <= 19'h0006c; 
        10'b0101001110: data <= 19'h00115; 
        10'b0101001111: data <= 19'h7ff59; 
        10'b0101010000: data <= 19'h7ff53; 
        10'b0101010001: data <= 19'h7ff72; 
        10'b0101010010: data <= 19'h7ff30; 
        10'b0101010011: data <= 19'h7fede; 
        10'b0101010100: data <= 19'h7ff24; 
        10'b0101010101: data <= 19'h0022d; 
        10'b0101010110: data <= 19'h004ef; 
        10'b0101010111: data <= 19'h00467; 
        10'b0101011000: data <= 19'h0033d; 
        10'b0101011001: data <= 19'h001da; 
        10'b0101011010: data <= 19'h00578; 
        10'b0101011011: data <= 19'h00b51; 
        10'b0101011100: data <= 19'h00a92; 
        10'b0101011101: data <= 19'h00ad6; 
        10'b0101011110: data <= 19'h0011e; 
        10'b0101011111: data <= 19'h7fa81; 
        10'b0101100000: data <= 19'h7f5c7; 
        10'b0101100001: data <= 19'h7f7ba; 
        10'b0101100010: data <= 19'h7fa62; 
        10'b0101100011: data <= 19'h7f7f0; 
        10'b0101100100: data <= 19'h7f6d1; 
        10'b0101100101: data <= 19'h7f0c1; 
        10'b0101100110: data <= 19'h7ee9b; 
        10'b0101100111: data <= 19'h7f0e4; 
        10'b0101101000: data <= 19'h7f5e5; 
        10'b0101101001: data <= 19'h7fd22; 
        10'b0101101010: data <= 19'h00026; 
        10'b0101101011: data <= 19'h7fffe; 
        10'b0101101100: data <= 19'h7ff66; 
        10'b0101101101: data <= 19'h7fe92; 
        10'b0101101110: data <= 19'h7fe7a; 
        10'b0101101111: data <= 19'h7fef0; 
        10'b0101110000: data <= 19'h7ffad; 
        10'b0101110001: data <= 19'h00124; 
        10'b0101110010: data <= 19'h0034e; 
        10'b0101110011: data <= 19'h0026d; 
        10'b0101110100: data <= 19'h002cd; 
        10'b0101110101: data <= 19'h00251; 
        10'b0101110110: data <= 19'h0079d; 
        10'b0101110111: data <= 19'h00882; 
        10'b0101111000: data <= 19'h00654; 
        10'b0101111001: data <= 19'h005e9; 
        10'b0101111010: data <= 19'h7fed0; 
        10'b0101111011: data <= 19'h7f975; 
        10'b0101111100: data <= 19'h7f55a; 
        10'b0101111101: data <= 19'h7fa60; 
        10'b0101111110: data <= 19'h7fe01; 
        10'b0101111111: data <= 19'h7fdb0; 
        10'b0110000000: data <= 19'h7fee6; 
        10'b0110000001: data <= 19'h7fbaf; 
        10'b0110000010: data <= 19'h7f831; 
        10'b0110000011: data <= 19'h7f497; 
        10'b0110000100: data <= 19'h7f768; 
        10'b0110000101: data <= 19'h7fe82; 
        10'b0110000110: data <= 19'h7fe60; 
        10'b0110000111: data <= 19'h7ffc3; 
        10'b0110001000: data <= 19'h7ff6c; 
        10'b0110001001: data <= 19'h7fe74; 
        10'b0110001010: data <= 19'h7ff3c; 
        10'b0110001011: data <= 19'h7fe15; 
        10'b0110001100: data <= 19'h7ff5b; 
        10'b0110001101: data <= 19'h7ff4e; 
        10'b0110001110: data <= 19'h7fff7; 
        10'b0110001111: data <= 19'h7ffa2; 
        10'b0110010000: data <= 19'h00380; 
        10'b0110010001: data <= 19'h00589; 
        10'b0110010010: data <= 19'h006a4; 
        10'b0110010011: data <= 19'h00145; 
        10'b0110010100: data <= 19'h0023f; 
        10'b0110010101: data <= 19'h7ff95; 
        10'b0110010110: data <= 19'h7fb40; 
        10'b0110010111: data <= 19'h7fa87; 
        10'b0110011000: data <= 19'h7f868; 
        10'b0110011001: data <= 19'h7f949; 
        10'b0110011010: data <= 19'h7f9b5; 
        10'b0110011011: data <= 19'h7fcf7; 
        10'b0110011100: data <= 19'h7fd60; 
        10'b0110011101: data <= 19'h7fd9e; 
        10'b0110011110: data <= 19'h7fe8e; 
        10'b0110011111: data <= 19'h7f9bb; 
        10'b0110100000: data <= 19'h7fbc8; 
        10'b0110100001: data <= 19'h7fde3; 
        10'b0110100010: data <= 19'h7ff40; 
        10'b0110100011: data <= 19'h7fe21; 
        10'b0110100100: data <= 19'h7fe53; 
        10'b0110100101: data <= 19'h00042; 
        10'b0110100110: data <= 19'h7fe32; 
        10'b0110100111: data <= 19'h7ff43; 
        10'b0110101000: data <= 19'h7fd52; 
        10'b0110101001: data <= 19'h7fbf9; 
        10'b0110101010: data <= 19'h7fa5d; 
        10'b0110101011: data <= 19'h7fc44; 
        10'b0110101100: data <= 19'h0015c; 
        10'b0110101101: data <= 19'h0063c; 
        10'b0110101110: data <= 19'h002f6; 
        10'b0110101111: data <= 19'h002bb; 
        10'b0110110000: data <= 19'h0025b; 
        10'b0110110001: data <= 19'h7fddf; 
        10'b0110110010: data <= 19'h7f8f2; 
        10'b0110110011: data <= 19'h7f7e3; 
        10'b0110110100: data <= 19'h7f8ae; 
        10'b0110110101: data <= 19'h7f87f; 
        10'b0110110110: data <= 19'h7fab7; 
        10'b0110110111: data <= 19'h7ffbc; 
        10'b0110111000: data <= 19'h7fe34; 
        10'b0110111001: data <= 19'h7fe7c; 
        10'b0110111010: data <= 19'h7fe30; 
        10'b0110111011: data <= 19'h7fdea; 
        10'b0110111100: data <= 19'h7fe89; 
        10'b0110111101: data <= 19'h7fff4; 
        10'b0110111110: data <= 19'h0004a; 
        10'b0110111111: data <= 19'h7fee1; 
        10'b0111000000: data <= 19'h7fefe; 
        10'b0111000001: data <= 19'h7ff58; 
        10'b0111000010: data <= 19'h7ff90; 
        10'b0111000011: data <= 19'h7fe33; 
        10'b0111000100: data <= 19'h7fef4; 
        10'b0111000101: data <= 19'h7fb6b; 
        10'b0111000110: data <= 19'h7f6d3; 
        10'b0111000111: data <= 19'h7f526; 
        10'b0111001000: data <= 19'h7f8a9; 
        10'b0111001001: data <= 19'h7fbf1; 
        10'b0111001010: data <= 19'h7fe64; 
        10'b0111001011: data <= 19'h7fdaf; 
        10'b0111001100: data <= 19'h7fe7d; 
        10'b0111001101: data <= 19'h7fb00; 
        10'b0111001110: data <= 19'h7f65e; 
        10'b0111001111: data <= 19'h7f82e; 
        10'b0111010000: data <= 19'h7fa51; 
        10'b0111010001: data <= 19'h7fdf4; 
        10'b0111010010: data <= 19'h7fe13; 
        10'b0111010011: data <= 19'h00050; 
        10'b0111010100: data <= 19'h00195; 
        10'b0111010101: data <= 19'h00040; 
        10'b0111010110: data <= 19'h001b8; 
        10'b0111010111: data <= 19'h00064; 
        10'b0111011000: data <= 19'h00045; 
        10'b0111011001: data <= 19'h0003e; 
        10'b0111011010: data <= 19'h7feec; 
        10'b0111011011: data <= 19'h7ff01; 
        10'b0111011100: data <= 19'h7fece; 
        10'b0111011101: data <= 19'h7ffec; 
        10'b0111011110: data <= 19'h7ffff; 
        10'b0111011111: data <= 19'h00022; 
        10'b0111100000: data <= 19'h7fed6; 
        10'b0111100001: data <= 19'h00056; 
        10'b0111100010: data <= 19'h000ac; 
        10'b0111100011: data <= 19'h7f8d6; 
        10'b0111100100: data <= 19'h7f309; 
        10'b0111100101: data <= 19'h7f3de; 
        10'b0111100110: data <= 19'h7f74f; 
        10'b0111100111: data <= 19'h7fac6; 
        10'b0111101000: data <= 19'h7f7d4; 
        10'b0111101001: data <= 19'h7f574; 
        10'b0111101010: data <= 19'h7f5bf; 
        10'b0111101011: data <= 19'h7fb54; 
        10'b0111101100: data <= 19'h7fdf3; 
        10'b0111101101: data <= 19'h0031a; 
        10'b0111101110: data <= 19'h004bd; 
        10'b0111101111: data <= 19'h00319; 
        10'b0111110000: data <= 19'h00320; 
        10'b0111110001: data <= 19'h000e8; 
        10'b0111110010: data <= 19'h0001a; 
        10'b0111110011: data <= 19'h001ba; 
        10'b0111110100: data <= 19'h001c1; 
        10'b0111110101: data <= 19'h7fe85; 
        10'b0111110110: data <= 19'h7fff1; 
        10'b0111110111: data <= 19'h0000a; 
        10'b0111111000: data <= 19'h0002d; 
        10'b0111111001: data <= 19'h7febe; 
        10'b0111111010: data <= 19'h7ff34; 
        10'b0111111011: data <= 19'h7fefa; 
        10'b0111111100: data <= 19'h00291; 
        10'b0111111101: data <= 19'h00364; 
        10'b0111111110: data <= 19'h0080d; 
        10'b0111111111: data <= 19'h0016a; 
        10'b1000000000: data <= 19'h7f83f; 
        10'b1000000001: data <= 19'h7f4b8; 
        10'b1000000010: data <= 19'h7f127; 
        10'b1000000011: data <= 19'h7f2bd; 
        10'b1000000100: data <= 19'h7f67d; 
        10'b1000000101: data <= 19'h7fa92; 
        10'b1000000110: data <= 19'h7fd4a; 
        10'b1000000111: data <= 19'h7fedd; 
        10'b1000001000: data <= 19'h7ffcc; 
        10'b1000001001: data <= 19'h003a4; 
        10'b1000001010: data <= 19'h001d4; 
        10'b1000001011: data <= 19'h0033f; 
        10'b1000001100: data <= 19'h0022f; 
        10'b1000001101: data <= 19'h0032a; 
        10'b1000001110: data <= 19'h0029c; 
        10'b1000001111: data <= 19'h0039b; 
        10'b1000010000: data <= 19'h001e0; 
        10'b1000010001: data <= 19'h00024; 
        10'b1000010010: data <= 19'h7fea1; 
        10'b1000010011: data <= 19'h7ff8f; 
        10'b1000010100: data <= 19'h00002; 
        10'b1000010101: data <= 19'h7febb; 
        10'b1000010110: data <= 19'h7ff52; 
        10'b1000010111: data <= 19'h00046; 
        10'b1000011000: data <= 19'h003e5; 
        10'b1000011001: data <= 19'h006a6; 
        10'b1000011010: data <= 19'h008f4; 
        10'b1000011011: data <= 19'h00607; 
        10'b1000011100: data <= 19'h003d1; 
        10'b1000011101: data <= 19'h0013d; 
        10'b1000011110: data <= 19'h7fd26; 
        10'b1000011111: data <= 19'h7fcf5; 
        10'b1000100000: data <= 19'h00042; 
        10'b1000100001: data <= 19'h003a6; 
        10'b1000100010: data <= 19'h0015d; 
        10'b1000100011: data <= 19'h001f0; 
        10'b1000100100: data <= 19'h001f7; 
        10'b1000100101: data <= 19'h7ff61; 
        10'b1000100110: data <= 19'h00169; 
        10'b1000100111: data <= 19'h00161; 
        10'b1000101000: data <= 19'h0004b; 
        10'b1000101001: data <= 19'h0025d; 
        10'b1000101010: data <= 19'h00410; 
        10'b1000101011: data <= 19'h002f8; 
        10'b1000101100: data <= 19'h0003f; 
        10'b1000101101: data <= 19'h7fff3; 
        10'b1000101110: data <= 19'h7fffd; 
        10'b1000101111: data <= 19'h7fe68; 
        10'b1000110000: data <= 19'h7ffeb; 
        10'b1000110001: data <= 19'h7fe24; 
        10'b1000110010: data <= 19'h7ff1d; 
        10'b1000110011: data <= 19'h7fe9c; 
        10'b1000110100: data <= 19'h00086; 
        10'b1000110101: data <= 19'h00460; 
        10'b1000110110: data <= 19'h00514; 
        10'b1000110111: data <= 19'h00630; 
        10'b1000111000: data <= 19'h008ac; 
        10'b1000111001: data <= 19'h00753; 
        10'b1000111010: data <= 19'h0066f; 
        10'b1000111011: data <= 19'h00961; 
        10'b1000111100: data <= 19'h005d7; 
        10'b1000111101: data <= 19'h00461; 
        10'b1000111110: data <= 19'h7fec4; 
        10'b1000111111: data <= 19'h7fede; 
        10'b1001000000: data <= 19'h0033a; 
        10'b1001000001: data <= 19'h001a7; 
        10'b1001000010: data <= 19'h002b2; 
        10'b1001000011: data <= 19'h00391; 
        10'b1001000100: data <= 19'h00320; 
        10'b1001000101: data <= 19'h00274; 
        10'b1001000110: data <= 19'h005de; 
        10'b1001000111: data <= 19'h00463; 
        10'b1001001000: data <= 19'h7ff6e; 
        10'b1001001001: data <= 19'h7fe2d; 
        10'b1001001010: data <= 19'h7ff5b; 
        10'b1001001011: data <= 19'h7fed8; 
        10'b1001001100: data <= 19'h7fead; 
        10'b1001001101: data <= 19'h0000b; 
        10'b1001001110: data <= 19'h7fe10; 
        10'b1001001111: data <= 19'h7ff46; 
        10'b1001010000: data <= 19'h001ba; 
        10'b1001010001: data <= 19'h7ff73; 
        10'b1001010010: data <= 19'h00217; 
        10'b1001010011: data <= 19'h005a9; 
        10'b1001010100: data <= 19'h0082c; 
        10'b1001010101: data <= 19'h00558; 
        10'b1001010110: data <= 19'h00489; 
        10'b1001010111: data <= 19'h00272; 
        10'b1001011000: data <= 19'h0032a; 
        10'b1001011001: data <= 19'h001f7; 
        10'b1001011010: data <= 19'h0020c; 
        10'b1001011011: data <= 19'h0027f; 
        10'b1001011100: data <= 19'h000a6; 
        10'b1001011101: data <= 19'h00203; 
        10'b1001011110: data <= 19'h00107; 
        10'b1001011111: data <= 19'h0033d; 
        10'b1001100000: data <= 19'h0032e; 
        10'b1001100001: data <= 19'h00556; 
        10'b1001100010: data <= 19'h00690; 
        10'b1001100011: data <= 19'h0016b; 
        10'b1001100100: data <= 19'h0000e; 
        10'b1001100101: data <= 19'h7fe71; 
        10'b1001100110: data <= 19'h7fedd; 
        10'b1001100111: data <= 19'h7fede; 
        10'b1001101000: data <= 19'h7ff9e; 
        10'b1001101001: data <= 19'h7fe3a; 
        10'b1001101010: data <= 19'h7ff14; 
        10'b1001101011: data <= 19'h7fedd; 
        10'b1001101100: data <= 19'h0009f; 
        10'b1001101101: data <= 19'h7ff20; 
        10'b1001101110: data <= 19'h7fe16; 
        10'b1001101111: data <= 19'h7ffa9; 
        10'b1001110000: data <= 19'h0032d; 
        10'b1001110001: data <= 19'h004a5; 
        10'b1001110010: data <= 19'h000ce; 
        10'b1001110011: data <= 19'h0041d; 
        10'b1001110100: data <= 19'h006a6; 
        10'b1001110101: data <= 19'h00836; 
        10'b1001110110: data <= 19'h0042e; 
        10'b1001110111: data <= 19'h000a1; 
        10'b1001111000: data <= 19'h00076; 
        10'b1001111001: data <= 19'h00106; 
        10'b1001111010: data <= 19'h00227; 
        10'b1001111011: data <= 19'h00224; 
        10'b1001111100: data <= 19'h003ab; 
        10'b1001111101: data <= 19'h00350; 
        10'b1001111110: data <= 19'h00376; 
        10'b1001111111: data <= 19'h00138; 
        10'b1010000000: data <= 19'h7ffd2; 
        10'b1010000001: data <= 19'h00032; 
        10'b1010000010: data <= 19'h7ff55; 
        10'b1010000011: data <= 19'h7ff8d; 
        10'b1010000100: data <= 19'h7fe8a; 
        10'b1010000101: data <= 19'h7ff49; 
        10'b1010000110: data <= 19'h7ff96; 
        10'b1010000111: data <= 19'h7ff6e; 
        10'b1010001000: data <= 19'h7fe9d; 
        10'b1010001001: data <= 19'h7ff16; 
        10'b1010001010: data <= 19'h7fd38; 
        10'b1010001011: data <= 19'h7febc; 
        10'b1010001100: data <= 19'h00284; 
        10'b1010001101: data <= 19'h00277; 
        10'b1010001110: data <= 19'h00275; 
        10'b1010001111: data <= 19'h00462; 
        10'b1010010000: data <= 19'h00435; 
        10'b1010010001: data <= 19'h002e1; 
        10'b1010010010: data <= 19'h0034f; 
        10'b1010010011: data <= 19'h00308; 
        10'b1010010100: data <= 19'h002f7; 
        10'b1010010101: data <= 19'h0015d; 
        10'b1010010110: data <= 19'h7fe6f; 
        10'b1010010111: data <= 19'h7ffc8; 
        10'b1010011000: data <= 19'h00174; 
        10'b1010011001: data <= 19'h00097; 
        10'b1010011010: data <= 19'h001f2; 
        10'b1010011011: data <= 19'h7fec8; 
        10'b1010011100: data <= 19'h00054; 
        10'b1010011101: data <= 19'h7ff01; 
        10'b1010011110: data <= 19'h7fefb; 
        10'b1010011111: data <= 19'h0004e; 
        10'b1010100000: data <= 19'h7ffdc; 
        10'b1010100001: data <= 19'h7ff0b; 
        10'b1010100010: data <= 19'h7fee6; 
        10'b1010100011: data <= 19'h00057; 
        10'b1010100100: data <= 19'h7fe19; 
        10'b1010100101: data <= 19'h7fdfb; 
        10'b1010100110: data <= 19'h7ff46; 
        10'b1010100111: data <= 19'h7ffa2; 
        10'b1010101000: data <= 19'h7ffe3; 
        10'b1010101001: data <= 19'h00341; 
        10'b1010101010: data <= 19'h00439; 
        10'b1010101011: data <= 19'h00340; 
        10'b1010101100: data <= 19'h0021d; 
        10'b1010101101: data <= 19'h002f0; 
        10'b1010101110: data <= 19'h0056c; 
        10'b1010101111: data <= 19'h0047c; 
        10'b1010110000: data <= 19'h002ad; 
        10'b1010110001: data <= 19'h0014d; 
        10'b1010110010: data <= 19'h0027c; 
        10'b1010110011: data <= 19'h0019c; 
        10'b1010110100: data <= 19'h7ffe8; 
        10'b1010110101: data <= 19'h7ffc5; 
        10'b1010110110: data <= 19'h7ff69; 
        10'b1010110111: data <= 19'h0001a; 
        10'b1010111000: data <= 19'h7feb1; 
        10'b1010111001: data <= 19'h7ff88; 
        10'b1010111010: data <= 19'h00032; 
        10'b1010111011: data <= 19'h7fe66; 
        10'b1010111100: data <= 19'h7ff48; 
        10'b1010111101: data <= 19'h00011; 
        10'b1010111110: data <= 19'h00030; 
        10'b1010111111: data <= 19'h7fe52; 
        10'b1011000000: data <= 19'h7fffd; 
        10'b1011000001: data <= 19'h7ff7b; 
        10'b1011000010: data <= 19'h7fe01; 
        10'b1011000011: data <= 19'h7ff43; 
        10'b1011000100: data <= 19'h7fe35; 
        10'b1011000101: data <= 19'h0010f; 
        10'b1011000110: data <= 19'h000ca; 
        10'b1011000111: data <= 19'h00233; 
        10'b1011001000: data <= 19'h00230; 
        10'b1011001001: data <= 19'h003d6; 
        10'b1011001010: data <= 19'h00036; 
        10'b1011001011: data <= 19'h00124; 
        10'b1011001100: data <= 19'h000f7; 
        10'b1011001101: data <= 19'h001e1; 
        10'b1011001110: data <= 19'h7febe; 
        10'b1011001111: data <= 19'h7fff2; 
        10'b1011010000: data <= 19'h7fde7; 
        10'b1011010001: data <= 19'h0002e; 
        10'b1011010010: data <= 19'h7ff38; 
        10'b1011010011: data <= 19'h7fe98; 
        10'b1011010100: data <= 19'h7ffd5; 
        10'b1011010101: data <= 19'h00018; 
        10'b1011010110: data <= 19'h7fe37; 
        10'b1011010111: data <= 19'h7ff0e; 
        10'b1011011000: data <= 19'h7ff71; 
        10'b1011011001: data <= 19'h7ff62; 
        10'b1011011010: data <= 19'h7feb0; 
        10'b1011011011: data <= 19'h7ff01; 
        10'b1011011100: data <= 19'h7fee5; 
        10'b1011011101: data <= 19'h7ff18; 
        10'b1011011110: data <= 19'h7ffac; 
        10'b1011011111: data <= 19'h7feb3; 
        10'b1011100000: data <= 19'h7fe48; 
        10'b1011100001: data <= 19'h7ff1b; 
        10'b1011100010: data <= 19'h7fed3; 
        10'b1011100011: data <= 19'h7ffc7; 
        10'b1011100100: data <= 19'h00009; 
        10'b1011100101: data <= 19'h7ff8d; 
        10'b1011100110: data <= 19'h7febf; 
        10'b1011100111: data <= 19'h7ff5c; 
        10'b1011101000: data <= 19'h7ffb7; 
        10'b1011101001: data <= 19'h7feb1; 
        10'b1011101010: data <= 19'h7fd79; 
        10'b1011101011: data <= 19'h7fdf4; 
        10'b1011101100: data <= 19'h7ff91; 
        10'b1011101101: data <= 19'h7ff8f; 
        10'b1011101110: data <= 19'h7fed9; 
        10'b1011101111: data <= 19'h7ffaa; 
        10'b1011110000: data <= 19'h7ff24; 
        10'b1011110001: data <= 19'h7ff6a; 
        10'b1011110010: data <= 19'h7fef0; 
        10'b1011110011: data <= 19'h7fe36; 
        10'b1011110100: data <= 19'h7ff9b; 
        10'b1011110101: data <= 19'h7ffc2; 
        10'b1011110110: data <= 19'h7ffd5; 
        10'b1011110111: data <= 19'h7ff7f; 
        10'b1011111000: data <= 19'h7fe79; 
        10'b1011111001: data <= 19'h7ffe8; 
        10'b1011111010: data <= 19'h7fef9; 
        10'b1011111011: data <= 19'h7fee0; 
        10'b1011111100: data <= 19'h0005f; 
        10'b1011111101: data <= 19'h7feed; 
        10'b1011111110: data <= 19'h7fec7; 
        10'b1011111111: data <= 19'h7ffdb; 
        10'b1100000000: data <= 19'h7ff57; 
        10'b1100000001: data <= 19'h7fe20; 
        10'b1100000010: data <= 19'h0000a; 
        10'b1100000011: data <= 19'h7ff6c; 
        10'b1100000100: data <= 19'h7fe4d; 
        10'b1100000101: data <= 19'h7fe1d; 
        10'b1100000110: data <= 19'h7fe97; 
        10'b1100000111: data <= 19'h7fe16; 
        10'b1100001000: data <= 19'h7fff9; 
        10'b1100001001: data <= 19'h7fef2; 
        10'b1100001010: data <= 19'h0005a; 
        10'b1100001011: data <= 19'h7fe5f; 
        10'b1100001100: data <= 19'h7ff83; 
        10'b1100001101: data <= 19'h7ff2f; 
        10'b1100001110: data <= 19'h7fe7f; 
        10'b1100001111: data <= 19'h7ffc4; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 14) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 20'hffdc8; 
        10'b0000000001: data <= 20'hfffb0; 
        10'b0000000010: data <= 20'hfffae; 
        10'b0000000011: data <= 20'hffd04; 
        10'b0000000100: data <= 20'hffe99; 
        10'b0000000101: data <= 20'hffe38; 
        10'b0000000110: data <= 20'hffffd; 
        10'b0000000111: data <= 20'hffe15; 
        10'b0000001000: data <= 20'hfff35; 
        10'b0000001001: data <= 20'h000a5; 
        10'b0000001010: data <= 20'hfff35; 
        10'b0000001011: data <= 20'hfff23; 
        10'b0000001100: data <= 20'hffdba; 
        10'b0000001101: data <= 20'hfffdd; 
        10'b0000001110: data <= 20'hffcf8; 
        10'b0000001111: data <= 20'hffd80; 
        10'b0000010000: data <= 20'hffc90; 
        10'b0000010001: data <= 20'hffd35; 
        10'b0000010010: data <= 20'hfff97; 
        10'b0000010011: data <= 20'hfff3c; 
        10'b0000010100: data <= 20'hffc86; 
        10'b0000010101: data <= 20'hffeae; 
        10'b0000010110: data <= 20'hfff0b; 
        10'b0000010111: data <= 20'hffe4a; 
        10'b0000011000: data <= 20'hffcba; 
        10'b0000011001: data <= 20'hffec3; 
        10'b0000011010: data <= 20'hfff0a; 
        10'b0000011011: data <= 20'hffde1; 
        10'b0000011100: data <= 20'hfffcc; 
        10'b0000011101: data <= 20'hffc5b; 
        10'b0000011110: data <= 20'hffffa; 
        10'b0000011111: data <= 20'hffcdf; 
        10'b0000100000: data <= 20'hfffdd; 
        10'b0000100001: data <= 20'hffdff; 
        10'b0000100010: data <= 20'hffef8; 
        10'b0000100011: data <= 20'hffdea; 
        10'b0000100100: data <= 20'hffd62; 
        10'b0000100101: data <= 20'hfff0b; 
        10'b0000100110: data <= 20'h00052; 
        10'b0000100111: data <= 20'hffcf5; 
        10'b0000101000: data <= 20'hffde2; 
        10'b0000101001: data <= 20'hffd49; 
        10'b0000101010: data <= 20'hffc81; 
        10'b0000101011: data <= 20'hfff6b; 
        10'b0000101100: data <= 20'hffda1; 
        10'b0000101101: data <= 20'hffd3b; 
        10'b0000101110: data <= 20'hffdb3; 
        10'b0000101111: data <= 20'hffd8c; 
        10'b0000110000: data <= 20'hfff39; 
        10'b0000110001: data <= 20'hffcd3; 
        10'b0000110010: data <= 20'hffff3; 
        10'b0000110011: data <= 20'hffd0b; 
        10'b0000110100: data <= 20'h0000b; 
        10'b0000110101: data <= 20'hfffc2; 
        10'b0000110110: data <= 20'hffd2a; 
        10'b0000110111: data <= 20'hffe6f; 
        10'b0000111000: data <= 20'hffe79; 
        10'b0000111001: data <= 20'hfff54; 
        10'b0000111010: data <= 20'hffde6; 
        10'b0000111011: data <= 20'hffc87; 
        10'b0000111100: data <= 20'hffd23; 
        10'b0000111101: data <= 20'hffeca; 
        10'b0000111110: data <= 20'hfffe2; 
        10'b0000111111: data <= 20'hfff0f; 
        10'b0001000000: data <= 20'hffd7c; 
        10'b0001000001: data <= 20'hffe13; 
        10'b0001000010: data <= 20'h0007b; 
        10'b0001000011: data <= 20'hffc4d; 
        10'b0001000100: data <= 20'hfffd4; 
        10'b0001000101: data <= 20'hffd66; 
        10'b0001000110: data <= 20'hffc9c; 
        10'b0001000111: data <= 20'hffd3d; 
        10'b0001001000: data <= 20'hffdc9; 
        10'b0001001001: data <= 20'hffeb8; 
        10'b0001001010: data <= 20'hffe14; 
        10'b0001001011: data <= 20'hffe1b; 
        10'b0001001100: data <= 20'h000d9; 
        10'b0001001101: data <= 20'h00018; 
        10'b0001001110: data <= 20'h0005b; 
        10'b0001001111: data <= 20'hffd52; 
        10'b0001010000: data <= 20'hffc83; 
        10'b0001010001: data <= 20'hffe44; 
        10'b0001010010: data <= 20'hfffca; 
        10'b0001010011: data <= 20'hfff0d; 
        10'b0001010100: data <= 20'hfff58; 
        10'b0001010101: data <= 20'hffeff; 
        10'b0001010110: data <= 20'hffd2c; 
        10'b0001010111: data <= 20'hfffd2; 
        10'b0001011000: data <= 20'hffce3; 
        10'b0001011001: data <= 20'hffdf0; 
        10'b0001011010: data <= 20'hffc4c; 
        10'b0001011011: data <= 20'hffd95; 
        10'b0001011100: data <= 20'hffc90; 
        10'b0001011101: data <= 20'hffd8b; 
        10'b0001011110: data <= 20'hffa05; 
        10'b0001011111: data <= 20'hff85d; 
        10'b0001100000: data <= 20'hffba3; 
        10'b0001100001: data <= 20'hffbe9; 
        10'b0001100010: data <= 20'hffaf9; 
        10'b0001100011: data <= 20'hffe56; 
        10'b0001100100: data <= 20'hfff48; 
        10'b0001100101: data <= 20'hffc0e; 
        10'b0001100110: data <= 20'hffda2; 
        10'b0001100111: data <= 20'hfff41; 
        10'b0001101000: data <= 20'hfff76; 
        10'b0001101001: data <= 20'hffe5c; 
        10'b0001101010: data <= 20'hffbff; 
        10'b0001101011: data <= 20'hffd4f; 
        10'b0001101100: data <= 20'hffb2b; 
        10'b0001101101: data <= 20'h0008e; 
        10'b0001101110: data <= 20'h00059; 
        10'b0001101111: data <= 20'hffcd7; 
        10'b0001110000: data <= 20'hffca2; 
        10'b0001110001: data <= 20'hffde9; 
        10'b0001110010: data <= 20'h00057; 
        10'b0001110011: data <= 20'h00030; 
        10'b0001110100: data <= 20'h00077; 
        10'b0001110101: data <= 20'hffd95; 
        10'b0001110110: data <= 20'hffd66; 
        10'b0001110111: data <= 20'hffa99; 
        10'b0001111000: data <= 20'hff6e4; 
        10'b0001111001: data <= 20'hff3e7; 
        10'b0001111010: data <= 20'hfee56; 
        10'b0001111011: data <= 20'hff4b7; 
        10'b0001111100: data <= 20'hff49f; 
        10'b0001111101: data <= 20'hff0bd; 
        10'b0001111110: data <= 20'hff798; 
        10'b0001111111: data <= 20'hffff6; 
        10'b0010000000: data <= 20'hfff00; 
        10'b0010000001: data <= 20'h002d9; 
        10'b0010000010: data <= 20'hfff23; 
        10'b0010000011: data <= 20'hffbab; 
        10'b0010000100: data <= 20'hffa56; 
        10'b0010000101: data <= 20'hffd01; 
        10'b0010000110: data <= 20'hffd8b; 
        10'b0010000111: data <= 20'hffe48; 
        10'b0010001000: data <= 20'hffddf; 
        10'b0010001001: data <= 20'h000cc; 
        10'b0010001010: data <= 20'h00074; 
        10'b0010001011: data <= 20'hffe70; 
        10'b0010001100: data <= 20'hffeb7; 
        10'b0010001101: data <= 20'h000ca; 
        10'b0010001110: data <= 20'hffd45; 
        10'b0010001111: data <= 20'hffcdc; 
        10'b0010010000: data <= 20'hffdad; 
        10'b0010010001: data <= 20'hffa7b; 
        10'b0010010010: data <= 20'hff7aa; 
        10'b0010010011: data <= 20'hff7f2; 
        10'b0010010100: data <= 20'hffab9; 
        10'b0010010101: data <= 20'hfff03; 
        10'b0010010110: data <= 20'h001c7; 
        10'b0010010111: data <= 20'h001ec; 
        10'b0010011000: data <= 20'hffd24; 
        10'b0010011001: data <= 20'hffbea; 
        10'b0010011010: data <= 20'hffd89; 
        10'b0010011011: data <= 20'hffed8; 
        10'b0010011100: data <= 20'h00416; 
        10'b0010011101: data <= 20'h0042d; 
        10'b0010011110: data <= 20'h007eb; 
        10'b0010011111: data <= 20'h004ef; 
        10'b0010100000: data <= 20'h004c8; 
        10'b0010100001: data <= 20'h00623; 
        10'b0010100010: data <= 20'h00b53; 
        10'b0010100011: data <= 20'h009a2; 
        10'b0010100100: data <= 20'h006c2; 
        10'b0010100101: data <= 20'h003bd; 
        10'b0010100110: data <= 20'h00253; 
        10'b0010100111: data <= 20'h000de; 
        10'b0010101000: data <= 20'hffcfd; 
        10'b0010101001: data <= 20'hffcb7; 
        10'b0010101010: data <= 20'h0006b; 
        10'b0010101011: data <= 20'hffcd6; 
        10'b0010101100: data <= 20'hffbed; 
        10'b0010101101: data <= 20'hff645; 
        10'b0010101110: data <= 20'hffba1; 
        10'b0010101111: data <= 20'hfff7d; 
        10'b0010110000: data <= 20'hfffa8; 
        10'b0010110001: data <= 20'h003f3; 
        10'b0010110010: data <= 20'h00832; 
        10'b0010110011: data <= 20'h006d1; 
        10'b0010110100: data <= 20'h00128; 
        10'b0010110101: data <= 20'h00283; 
        10'b0010110110: data <= 20'hffedf; 
        10'b0010110111: data <= 20'hffc1e; 
        10'b0010111000: data <= 20'hffda6; 
        10'b0010111001: data <= 20'hffe04; 
        10'b0010111010: data <= 20'h00017; 
        10'b0010111011: data <= 20'h007c8; 
        10'b0010111100: data <= 20'h00474; 
        10'b0010111101: data <= 20'h0050f; 
        10'b0010111110: data <= 20'h00f76; 
        10'b0010111111: data <= 20'h01297; 
        10'b0011000000: data <= 20'h014ea; 
        10'b0011000001: data <= 20'h00b10; 
        10'b0011000010: data <= 20'h00577; 
        10'b0011000011: data <= 20'h00156; 
        10'b0011000100: data <= 20'hffe4b; 
        10'b0011000101: data <= 20'hfff14; 
        10'b0011000110: data <= 20'hffeaa; 
        10'b0011000111: data <= 20'hffbfe; 
        10'b0011001000: data <= 20'hff4b2; 
        10'b0011001001: data <= 20'hff2bb; 
        10'b0011001010: data <= 20'hff7ec; 
        10'b0011001011: data <= 20'h0010b; 
        10'b0011001100: data <= 20'h0054a; 
        10'b0011001101: data <= 20'h00a63; 
        10'b0011001110: data <= 20'h00a1d; 
        10'b0011001111: data <= 20'h008d5; 
        10'b0011010000: data <= 20'h0028e; 
        10'b0011010001: data <= 20'hfff2a; 
        10'b0011010010: data <= 20'hffd2d; 
        10'b0011010011: data <= 20'h00031; 
        10'b0011010100: data <= 20'h00460; 
        10'b0011010101: data <= 20'h003f5; 
        10'b0011010110: data <= 20'h00503; 
        10'b0011010111: data <= 20'h00b33; 
        10'b0011011000: data <= 20'h009af; 
        10'b0011011001: data <= 20'h00b94; 
        10'b0011011010: data <= 20'h01031; 
        10'b0011011011: data <= 20'h015b8; 
        10'b0011011100: data <= 20'h01a84; 
        10'b0011011101: data <= 20'h01325; 
        10'b0011011110: data <= 20'h002f3; 
        10'b0011011111: data <= 20'hfff8b; 
        10'b0011100000: data <= 20'hfff3e; 
        10'b0011100001: data <= 20'h000b3; 
        10'b0011100010: data <= 20'hffff0; 
        10'b0011100011: data <= 20'hffa8a; 
        10'b0011100100: data <= 20'hfefb7; 
        10'b0011100101: data <= 20'hff213; 
        10'b0011100110: data <= 20'hff5ed; 
        10'b0011100111: data <= 20'h000a0; 
        10'b0011101000: data <= 20'h007e0; 
        10'b0011101001: data <= 20'h00250; 
        10'b0011101010: data <= 20'h0043c; 
        10'b0011101011: data <= 20'h00837; 
        10'b0011101100: data <= 20'h00502; 
        10'b0011101101: data <= 20'hffa5d; 
        10'b0011101110: data <= 20'hff3a4; 
        10'b0011101111: data <= 20'hff883; 
        10'b0011110000: data <= 20'hffb68; 
        10'b0011110001: data <= 20'h00070; 
        10'b0011110010: data <= 20'h00143; 
        10'b0011110011: data <= 20'h00956; 
        10'b0011110100: data <= 20'h009da; 
        10'b0011110101: data <= 20'h00e09; 
        10'b0011110110: data <= 20'h0162f; 
        10'b0011110111: data <= 20'h01d07; 
        10'b0011111000: data <= 20'h026b9; 
        10'b0011111001: data <= 20'h01904; 
        10'b0011111010: data <= 20'h0048f; 
        10'b0011111011: data <= 20'hfff89; 
        10'b0011111100: data <= 20'hffccb; 
        10'b0011111101: data <= 20'hffe1f; 
        10'b0011111110: data <= 20'hffc80; 
        10'b0011111111: data <= 20'hff865; 
        10'b0100000000: data <= 20'hff744; 
        10'b0100000001: data <= 20'hff7ee; 
        10'b0100000010: data <= 20'h000fb; 
        10'b0100000011: data <= 20'hfff6f; 
        10'b0100000100: data <= 20'h006b8; 
        10'b0100000101: data <= 20'h005d6; 
        10'b0100000110: data <= 20'h0065a; 
        10'b0100000111: data <= 20'h010f4; 
        10'b0100001000: data <= 20'h00aef; 
        10'b0100001001: data <= 20'hffb77; 
        10'b0100001010: data <= 20'hff11a; 
        10'b0100001011: data <= 20'hfeaa4; 
        10'b0100001100: data <= 20'hfec0d; 
        10'b0100001101: data <= 20'hff464; 
        10'b0100001110: data <= 20'hffd57; 
        10'b0100001111: data <= 20'hfffed; 
        10'b0100010000: data <= 20'h00912; 
        10'b0100010001: data <= 20'h01364; 
        10'b0100010010: data <= 20'h01c10; 
        10'b0100010011: data <= 20'h02663; 
        10'b0100010100: data <= 20'h0303d; 
        10'b0100010101: data <= 20'h01fb2; 
        10'b0100010110: data <= 20'h005ad; 
        10'b0100010111: data <= 20'hffdc4; 
        10'b0100011000: data <= 20'hfff50; 
        10'b0100011001: data <= 20'hffdc9; 
        10'b0100011010: data <= 20'hffd03; 
        10'b0100011011: data <= 20'hffd97; 
        10'b0100011100: data <= 20'hffd74; 
        10'b0100011101: data <= 20'hffe5d; 
        10'b0100011110: data <= 20'h00569; 
        10'b0100011111: data <= 20'h00a16; 
        10'b0100100000: data <= 20'h00fbe; 
        10'b0100100001: data <= 20'h0116c; 
        10'b0100100010: data <= 20'h010a7; 
        10'b0100100011: data <= 20'h01427; 
        10'b0100100100: data <= 20'h010c2; 
        10'b0100100101: data <= 20'h00ce1; 
        10'b0100100110: data <= 20'hffd3e; 
        10'b0100100111: data <= 20'hff57a; 
        10'b0100101000: data <= 20'hfee6f; 
        10'b0100101001: data <= 20'hfeefe; 
        10'b0100101010: data <= 20'hfee64; 
        10'b0100101011: data <= 20'hfebed; 
        10'b0100101100: data <= 20'hff242; 
        10'b0100101101: data <= 20'hffbbb; 
        10'b0100101110: data <= 20'h00256; 
        10'b0100101111: data <= 20'h00ce2; 
        10'b0100110000: data <= 20'h019b5; 
        10'b0100110001: data <= 20'h01352; 
        10'b0100110010: data <= 20'h00693; 
        10'b0100110011: data <= 20'hffdc6; 
        10'b0100110100: data <= 20'hffcfe; 
        10'b0100110101: data <= 20'h00006; 
        10'b0100110110: data <= 20'hffd8d; 
        10'b0100110111: data <= 20'hffe65; 
        10'b0100111000: data <= 20'hffd83; 
        10'b0100111001: data <= 20'hfffa6; 
        10'b0100111010: data <= 20'h0089a; 
        10'b0100111011: data <= 20'h00a7f; 
        10'b0100111100: data <= 20'h00f2e; 
        10'b0100111101: data <= 20'h00e05; 
        10'b0100111110: data <= 20'h00a43; 
        10'b0100111111: data <= 20'h00b4e; 
        10'b0101000000: data <= 20'h012b5; 
        10'b0101000001: data <= 20'h01179; 
        10'b0101000010: data <= 20'h00047; 
        10'b0101000011: data <= 20'hff51e; 
        10'b0101000100: data <= 20'hff281; 
        10'b0101000101: data <= 20'hff177; 
        10'b0101000110: data <= 20'hfec9a; 
        10'b0101000111: data <= 20'hfe4ef; 
        10'b0101001000: data <= 20'hfd8b5; 
        10'b0101001001: data <= 20'hfdbec; 
        10'b0101001010: data <= 20'hfe270; 
        10'b0101001011: data <= 20'hfea71; 
        10'b0101001100: data <= 20'hff854; 
        10'b0101001101: data <= 20'h000d8; 
        10'b0101001110: data <= 20'h0022a; 
        10'b0101001111: data <= 20'hffeb1; 
        10'b0101010000: data <= 20'hffea7; 
        10'b0101010001: data <= 20'hffee3; 
        10'b0101010010: data <= 20'hffe61; 
        10'b0101010011: data <= 20'hffdbc; 
        10'b0101010100: data <= 20'hffe48; 
        10'b0101010101: data <= 20'h0045b; 
        10'b0101010110: data <= 20'h009de; 
        10'b0101010111: data <= 20'h008ce; 
        10'b0101011000: data <= 20'h00679; 
        10'b0101011001: data <= 20'h003b5; 
        10'b0101011010: data <= 20'h00aef; 
        10'b0101011011: data <= 20'h016a3; 
        10'b0101011100: data <= 20'h01525; 
        10'b0101011101: data <= 20'h015ac; 
        10'b0101011110: data <= 20'h0023c; 
        10'b0101011111: data <= 20'hff502; 
        10'b0101100000: data <= 20'hfeb8e; 
        10'b0101100001: data <= 20'hfef73; 
        10'b0101100010: data <= 20'hff4c5; 
        10'b0101100011: data <= 20'hfefe1; 
        10'b0101100100: data <= 20'hfeda2; 
        10'b0101100101: data <= 20'hfe183; 
        10'b0101100110: data <= 20'hfdd37; 
        10'b0101100111: data <= 20'hfe1c7; 
        10'b0101101000: data <= 20'hfebcb; 
        10'b0101101001: data <= 20'hffa43; 
        10'b0101101010: data <= 20'h0004c; 
        10'b0101101011: data <= 20'hffffb; 
        10'b0101101100: data <= 20'hffecd; 
        10'b0101101101: data <= 20'hffd24; 
        10'b0101101110: data <= 20'hffcf4; 
        10'b0101101111: data <= 20'hffde1; 
        10'b0101110000: data <= 20'hfff5a; 
        10'b0101110001: data <= 20'h00248; 
        10'b0101110010: data <= 20'h0069c; 
        10'b0101110011: data <= 20'h004d9; 
        10'b0101110100: data <= 20'h0059a; 
        10'b0101110101: data <= 20'h004a1; 
        10'b0101110110: data <= 20'h00f3a; 
        10'b0101110111: data <= 20'h01104; 
        10'b0101111000: data <= 20'h00ca8; 
        10'b0101111001: data <= 20'h00bd3; 
        10'b0101111010: data <= 20'hffda0; 
        10'b0101111011: data <= 20'hff2ea; 
        10'b0101111100: data <= 20'hfeab4; 
        10'b0101111101: data <= 20'hff4bf; 
        10'b0101111110: data <= 20'hffc01; 
        10'b0101111111: data <= 20'hffb60; 
        10'b0110000000: data <= 20'hffdcc; 
        10'b0110000001: data <= 20'hff75d; 
        10'b0110000010: data <= 20'hff062; 
        10'b0110000011: data <= 20'hfe92e; 
        10'b0110000100: data <= 20'hfeed0; 
        10'b0110000101: data <= 20'hffd05; 
        10'b0110000110: data <= 20'hffcc1; 
        10'b0110000111: data <= 20'hfff87; 
        10'b0110001000: data <= 20'hffed9; 
        10'b0110001001: data <= 20'hffce7; 
        10'b0110001010: data <= 20'hffe79; 
        10'b0110001011: data <= 20'hffc2b; 
        10'b0110001100: data <= 20'hffeb6; 
        10'b0110001101: data <= 20'hffe9c; 
        10'b0110001110: data <= 20'hfffee; 
        10'b0110001111: data <= 20'hfff45; 
        10'b0110010000: data <= 20'h00700; 
        10'b0110010001: data <= 20'h00b12; 
        10'b0110010010: data <= 20'h00d49; 
        10'b0110010011: data <= 20'h0028b; 
        10'b0110010100: data <= 20'h0047f; 
        10'b0110010101: data <= 20'hfff2b; 
        10'b0110010110: data <= 20'hff67f; 
        10'b0110010111: data <= 20'hff50e; 
        10'b0110011000: data <= 20'hff0cf; 
        10'b0110011001: data <= 20'hff292; 
        10'b0110011010: data <= 20'hff36b; 
        10'b0110011011: data <= 20'hff9ef; 
        10'b0110011100: data <= 20'hffac0; 
        10'b0110011101: data <= 20'hffb3b; 
        10'b0110011110: data <= 20'hffd1b; 
        10'b0110011111: data <= 20'hff377; 
        10'b0110100000: data <= 20'hff790; 
        10'b0110100001: data <= 20'hffbc5; 
        10'b0110100010: data <= 20'hffe7f; 
        10'b0110100011: data <= 20'hffc42; 
        10'b0110100100: data <= 20'hffca5; 
        10'b0110100101: data <= 20'h00084; 
        10'b0110100110: data <= 20'hffc63; 
        10'b0110100111: data <= 20'hffe86; 
        10'b0110101000: data <= 20'hffaa3; 
        10'b0110101001: data <= 20'hff7f2; 
        10'b0110101010: data <= 20'hff4ba; 
        10'b0110101011: data <= 20'hff888; 
        10'b0110101100: data <= 20'h002b7; 
        10'b0110101101: data <= 20'h00c78; 
        10'b0110101110: data <= 20'h005ec; 
        10'b0110101111: data <= 20'h00576; 
        10'b0110110000: data <= 20'h004b5; 
        10'b0110110001: data <= 20'hffbbf; 
        10'b0110110010: data <= 20'hff1e5; 
        10'b0110110011: data <= 20'hfefc6; 
        10'b0110110100: data <= 20'hff15c; 
        10'b0110110101: data <= 20'hff0ff; 
        10'b0110110110: data <= 20'hff56f; 
        10'b0110110111: data <= 20'hfff77; 
        10'b0110111000: data <= 20'hffc69; 
        10'b0110111001: data <= 20'hffcf8; 
        10'b0110111010: data <= 20'hffc5f; 
        10'b0110111011: data <= 20'hffbd4; 
        10'b0110111100: data <= 20'hffd13; 
        10'b0110111101: data <= 20'hfffe9; 
        10'b0110111110: data <= 20'h00095; 
        10'b0110111111: data <= 20'hffdc1; 
        10'b0111000000: data <= 20'hffdfb; 
        10'b0111000001: data <= 20'hffeb0; 
        10'b0111000010: data <= 20'hfff20; 
        10'b0111000011: data <= 20'hffc66; 
        10'b0111000100: data <= 20'hffde7; 
        10'b0111000101: data <= 20'hff6d7; 
        10'b0111000110: data <= 20'hfeda6; 
        10'b0111000111: data <= 20'hfea4c; 
        10'b0111001000: data <= 20'hff153; 
        10'b0111001001: data <= 20'hff7e1; 
        10'b0111001010: data <= 20'hffcc7; 
        10'b0111001011: data <= 20'hffb5d; 
        10'b0111001100: data <= 20'hffcfa; 
        10'b0111001101: data <= 20'hff5ff; 
        10'b0111001110: data <= 20'hfecbc; 
        10'b0111001111: data <= 20'hff05c; 
        10'b0111010000: data <= 20'hff4a3; 
        10'b0111010001: data <= 20'hffbe8; 
        10'b0111010010: data <= 20'hffc26; 
        10'b0111010011: data <= 20'h0009f; 
        10'b0111010100: data <= 20'h0032b; 
        10'b0111010101: data <= 20'h00080; 
        10'b0111010110: data <= 20'h00370; 
        10'b0111010111: data <= 20'h000c8; 
        10'b0111011000: data <= 20'h00089; 
        10'b0111011001: data <= 20'h0007c; 
        10'b0111011010: data <= 20'hffdd8; 
        10'b0111011011: data <= 20'hffe02; 
        10'b0111011100: data <= 20'hffd9c; 
        10'b0111011101: data <= 20'hfffd7; 
        10'b0111011110: data <= 20'hffffd; 
        10'b0111011111: data <= 20'h00043; 
        10'b0111100000: data <= 20'hffdad; 
        10'b0111100001: data <= 20'h000ab; 
        10'b0111100010: data <= 20'h00157; 
        10'b0111100011: data <= 20'hff1ab; 
        10'b0111100100: data <= 20'hfe613; 
        10'b0111100101: data <= 20'hfe7bd; 
        10'b0111100110: data <= 20'hfee9e; 
        10'b0111100111: data <= 20'hff58b; 
        10'b0111101000: data <= 20'hfefa7; 
        10'b0111101001: data <= 20'hfeae7; 
        10'b0111101010: data <= 20'hfeb7e; 
        10'b0111101011: data <= 20'hff6a9; 
        10'b0111101100: data <= 20'hffbe5; 
        10'b0111101101: data <= 20'h00633; 
        10'b0111101110: data <= 20'h0097b; 
        10'b0111101111: data <= 20'h00631; 
        10'b0111110000: data <= 20'h00640; 
        10'b0111110001: data <= 20'h001d1; 
        10'b0111110010: data <= 20'h00034; 
        10'b0111110011: data <= 20'h00373; 
        10'b0111110100: data <= 20'h00382; 
        10'b0111110101: data <= 20'hffd0b; 
        10'b0111110110: data <= 20'hfffe1; 
        10'b0111110111: data <= 20'h00015; 
        10'b0111111000: data <= 20'h00059; 
        10'b0111111001: data <= 20'hffd7c; 
        10'b0111111010: data <= 20'hffe69; 
        10'b0111111011: data <= 20'hffdf4; 
        10'b0111111100: data <= 20'h00521; 
        10'b0111111101: data <= 20'h006c7; 
        10'b0111111110: data <= 20'h0101a; 
        10'b0111111111: data <= 20'h002d5; 
        10'b1000000000: data <= 20'hff07f; 
        10'b1000000001: data <= 20'hfe96f; 
        10'b1000000010: data <= 20'hfe24e; 
        10'b1000000011: data <= 20'hfe57a; 
        10'b1000000100: data <= 20'hfecfb; 
        10'b1000000101: data <= 20'hff523; 
        10'b1000000110: data <= 20'hffa94; 
        10'b1000000111: data <= 20'hffdbb; 
        10'b1000001000: data <= 20'hfff98; 
        10'b1000001001: data <= 20'h00747; 
        10'b1000001010: data <= 20'h003a9; 
        10'b1000001011: data <= 20'h0067e; 
        10'b1000001100: data <= 20'h0045d; 
        10'b1000001101: data <= 20'h00655; 
        10'b1000001110: data <= 20'h00538; 
        10'b1000001111: data <= 20'h00737; 
        10'b1000010000: data <= 20'h003bf; 
        10'b1000010001: data <= 20'h00047; 
        10'b1000010010: data <= 20'hffd42; 
        10'b1000010011: data <= 20'hfff1e; 
        10'b1000010100: data <= 20'h00004; 
        10'b1000010101: data <= 20'hffd76; 
        10'b1000010110: data <= 20'hffea4; 
        10'b1000010111: data <= 20'h0008b; 
        10'b1000011000: data <= 20'h007c9; 
        10'b1000011001: data <= 20'h00d4d; 
        10'b1000011010: data <= 20'h011e8; 
        10'b1000011011: data <= 20'h00c0e; 
        10'b1000011100: data <= 20'h007a3; 
        10'b1000011101: data <= 20'h0027a; 
        10'b1000011110: data <= 20'hffa4d; 
        10'b1000011111: data <= 20'hff9ea; 
        10'b1000100000: data <= 20'h00084; 
        10'b1000100001: data <= 20'h0074c; 
        10'b1000100010: data <= 20'h002ba; 
        10'b1000100011: data <= 20'h003e0; 
        10'b1000100100: data <= 20'h003ef; 
        10'b1000100101: data <= 20'hffec3; 
        10'b1000100110: data <= 20'h002d3; 
        10'b1000100111: data <= 20'h002c2; 
        10'b1000101000: data <= 20'h00096; 
        10'b1000101001: data <= 20'h004bb; 
        10'b1000101010: data <= 20'h0081f; 
        10'b1000101011: data <= 20'h005f0; 
        10'b1000101100: data <= 20'h0007f; 
        10'b1000101101: data <= 20'hfffe7; 
        10'b1000101110: data <= 20'hffff9; 
        10'b1000101111: data <= 20'hffccf; 
        10'b1000110000: data <= 20'hfffd7; 
        10'b1000110001: data <= 20'hffc47; 
        10'b1000110010: data <= 20'hffe3a; 
        10'b1000110011: data <= 20'hffd39; 
        10'b1000110100: data <= 20'h0010b; 
        10'b1000110101: data <= 20'h008c0; 
        10'b1000110110: data <= 20'h00a29; 
        10'b1000110111: data <= 20'h00c60; 
        10'b1000111000: data <= 20'h01158; 
        10'b1000111001: data <= 20'h00ea6; 
        10'b1000111010: data <= 20'h00cde; 
        10'b1000111011: data <= 20'h012c2; 
        10'b1000111100: data <= 20'h00bad; 
        10'b1000111101: data <= 20'h008c2; 
        10'b1000111110: data <= 20'hffd89; 
        10'b1000111111: data <= 20'hffdbc; 
        10'b1001000000: data <= 20'h00674; 
        10'b1001000001: data <= 20'h0034d; 
        10'b1001000010: data <= 20'h00564; 
        10'b1001000011: data <= 20'h00722; 
        10'b1001000100: data <= 20'h0063f; 
        10'b1001000101: data <= 20'h004e8; 
        10'b1001000110: data <= 20'h00bbc; 
        10'b1001000111: data <= 20'h008c5; 
        10'b1001001000: data <= 20'hffedb; 
        10'b1001001001: data <= 20'hffc5a; 
        10'b1001001010: data <= 20'hffeb6; 
        10'b1001001011: data <= 20'hffdb0; 
        10'b1001001100: data <= 20'hffd59; 
        10'b1001001101: data <= 20'h00015; 
        10'b1001001110: data <= 20'hffc21; 
        10'b1001001111: data <= 20'hffe8c; 
        10'b1001010000: data <= 20'h00373; 
        10'b1001010001: data <= 20'hffee5; 
        10'b1001010010: data <= 20'h0042f; 
        10'b1001010011: data <= 20'h00b52; 
        10'b1001010100: data <= 20'h01059; 
        10'b1001010101: data <= 20'h00ab1; 
        10'b1001010110: data <= 20'h00912; 
        10'b1001010111: data <= 20'h004e3; 
        10'b1001011000: data <= 20'h00654; 
        10'b1001011001: data <= 20'h003ee; 
        10'b1001011010: data <= 20'h00418; 
        10'b1001011011: data <= 20'h004fd; 
        10'b1001011100: data <= 20'h0014c; 
        10'b1001011101: data <= 20'h00405; 
        10'b1001011110: data <= 20'h0020f; 
        10'b1001011111: data <= 20'h0067b; 
        10'b1001100000: data <= 20'h0065c; 
        10'b1001100001: data <= 20'h00aab; 
        10'b1001100010: data <= 20'h00d1f; 
        10'b1001100011: data <= 20'h002d6; 
        10'b1001100100: data <= 20'h0001d; 
        10'b1001100101: data <= 20'hffce2; 
        10'b1001100110: data <= 20'hffdba; 
        10'b1001100111: data <= 20'hffdbd; 
        10'b1001101000: data <= 20'hfff3b; 
        10'b1001101001: data <= 20'hffc74; 
        10'b1001101010: data <= 20'hffe29; 
        10'b1001101011: data <= 20'hffdb9; 
        10'b1001101100: data <= 20'h0013f; 
        10'b1001101101: data <= 20'hffe40; 
        10'b1001101110: data <= 20'hffc2c; 
        10'b1001101111: data <= 20'hfff51; 
        10'b1001110000: data <= 20'h0065a; 
        10'b1001110001: data <= 20'h0094a; 
        10'b1001110010: data <= 20'h0019c; 
        10'b1001110011: data <= 20'h00839; 
        10'b1001110100: data <= 20'h00d4d; 
        10'b1001110101: data <= 20'h0106c; 
        10'b1001110110: data <= 20'h0085c; 
        10'b1001110111: data <= 20'h00143; 
        10'b1001111000: data <= 20'h000ec; 
        10'b1001111001: data <= 20'h0020d; 
        10'b1001111010: data <= 20'h0044e; 
        10'b1001111011: data <= 20'h00448; 
        10'b1001111100: data <= 20'h00756; 
        10'b1001111101: data <= 20'h006a0; 
        10'b1001111110: data <= 20'h006ec; 
        10'b1001111111: data <= 20'h0026f; 
        10'b1010000000: data <= 20'hfffa5; 
        10'b1010000001: data <= 20'h00063; 
        10'b1010000010: data <= 20'hffea9; 
        10'b1010000011: data <= 20'hfff1a; 
        10'b1010000100: data <= 20'hffd14; 
        10'b1010000101: data <= 20'hffe93; 
        10'b1010000110: data <= 20'hfff2c; 
        10'b1010000111: data <= 20'hffedc; 
        10'b1010001000: data <= 20'hffd3a; 
        10'b1010001001: data <= 20'hffe2b; 
        10'b1010001010: data <= 20'hffa70; 
        10'b1010001011: data <= 20'hffd78; 
        10'b1010001100: data <= 20'h00508; 
        10'b1010001101: data <= 20'h004ed; 
        10'b1010001110: data <= 20'h004ea; 
        10'b1010001111: data <= 20'h008c4; 
        10'b1010010000: data <= 20'h0086a; 
        10'b1010010001: data <= 20'h005c3; 
        10'b1010010010: data <= 20'h0069e; 
        10'b1010010011: data <= 20'h00610; 
        10'b1010010100: data <= 20'h005ee; 
        10'b1010010101: data <= 20'h002ba; 
        10'b1010010110: data <= 20'hffcde; 
        10'b1010010111: data <= 20'hfff90; 
        10'b1010011000: data <= 20'h002e8; 
        10'b1010011001: data <= 20'h0012e; 
        10'b1010011010: data <= 20'h003e5; 
        10'b1010011011: data <= 20'hffd90; 
        10'b1010011100: data <= 20'h000a7; 
        10'b1010011101: data <= 20'hffe02; 
        10'b1010011110: data <= 20'hffdf6; 
        10'b1010011111: data <= 20'h0009c; 
        10'b1010100000: data <= 20'hfffb8; 
        10'b1010100001: data <= 20'hffe16; 
        10'b1010100010: data <= 20'hffdcb; 
        10'b1010100011: data <= 20'h000ae; 
        10'b1010100100: data <= 20'hffc31; 
        10'b1010100101: data <= 20'hffbf5; 
        10'b1010100110: data <= 20'hffe8c; 
        10'b1010100111: data <= 20'hfff43; 
        10'b1010101000: data <= 20'hfffc6; 
        10'b1010101001: data <= 20'h00683; 
        10'b1010101010: data <= 20'h00873; 
        10'b1010101011: data <= 20'h00681; 
        10'b1010101100: data <= 20'h00439; 
        10'b1010101101: data <= 20'h005e1; 
        10'b1010101110: data <= 20'h00ad8; 
        10'b1010101111: data <= 20'h008f9; 
        10'b1010110000: data <= 20'h0055a; 
        10'b1010110001: data <= 20'h0029a; 
        10'b1010110010: data <= 20'h004f8; 
        10'b1010110011: data <= 20'h00339; 
        10'b1010110100: data <= 20'hfffd0; 
        10'b1010110101: data <= 20'hfff89; 
        10'b1010110110: data <= 20'hffed2; 
        10'b1010110111: data <= 20'h00034; 
        10'b1010111000: data <= 20'hffd61; 
        10'b1010111001: data <= 20'hfff0f; 
        10'b1010111010: data <= 20'h00064; 
        10'b1010111011: data <= 20'hffccb; 
        10'b1010111100: data <= 20'hffe91; 
        10'b1010111101: data <= 20'h00022; 
        10'b1010111110: data <= 20'h00061; 
        10'b1010111111: data <= 20'hffca3; 
        10'b1011000000: data <= 20'hffffa; 
        10'b1011000001: data <= 20'hffef6; 
        10'b1011000010: data <= 20'hffc02; 
        10'b1011000011: data <= 20'hffe86; 
        10'b1011000100: data <= 20'hffc6a; 
        10'b1011000101: data <= 20'h0021e; 
        10'b1011000110: data <= 20'h00193; 
        10'b1011000111: data <= 20'h00467; 
        10'b1011001000: data <= 20'h00461; 
        10'b1011001001: data <= 20'h007ad; 
        10'b1011001010: data <= 20'h0006c; 
        10'b1011001011: data <= 20'h00249; 
        10'b1011001100: data <= 20'h001ee; 
        10'b1011001101: data <= 20'h003c2; 
        10'b1011001110: data <= 20'hffd7b; 
        10'b1011001111: data <= 20'hfffe4; 
        10'b1011010000: data <= 20'hffbcf; 
        10'b1011010001: data <= 20'h0005c; 
        10'b1011010010: data <= 20'hffe70; 
        10'b1011010011: data <= 20'hffd2f; 
        10'b1011010100: data <= 20'hfffab; 
        10'b1011010101: data <= 20'h00031; 
        10'b1011010110: data <= 20'hffc6e; 
        10'b1011010111: data <= 20'hffe1d; 
        10'b1011011000: data <= 20'hffee2; 
        10'b1011011001: data <= 20'hffec5; 
        10'b1011011010: data <= 20'hffd60; 
        10'b1011011011: data <= 20'hffe02; 
        10'b1011011100: data <= 20'hffdca; 
        10'b1011011101: data <= 20'hffe2f; 
        10'b1011011110: data <= 20'hfff59; 
        10'b1011011111: data <= 20'hffd65; 
        10'b1011100000: data <= 20'hffc90; 
        10'b1011100001: data <= 20'hffe36; 
        10'b1011100010: data <= 20'hffda7; 
        10'b1011100011: data <= 20'hfff8e; 
        10'b1011100100: data <= 20'h00012; 
        10'b1011100101: data <= 20'hfff19; 
        10'b1011100110: data <= 20'hffd7e; 
        10'b1011100111: data <= 20'hffeb8; 
        10'b1011101000: data <= 20'hfff6d; 
        10'b1011101001: data <= 20'hffd62; 
        10'b1011101010: data <= 20'hffaf2; 
        10'b1011101011: data <= 20'hffbe9; 
        10'b1011101100: data <= 20'hfff23; 
        10'b1011101101: data <= 20'hfff1e; 
        10'b1011101110: data <= 20'hffdb1; 
        10'b1011101111: data <= 20'hfff53; 
        10'b1011110000: data <= 20'hffe48; 
        10'b1011110001: data <= 20'hffed3; 
        10'b1011110010: data <= 20'hffddf; 
        10'b1011110011: data <= 20'hffc6d; 
        10'b1011110100: data <= 20'hfff36; 
        10'b1011110101: data <= 20'hfff84; 
        10'b1011110110: data <= 20'hfffa9; 
        10'b1011110111: data <= 20'hffefe; 
        10'b1011111000: data <= 20'hffcf2; 
        10'b1011111001: data <= 20'hfffcf; 
        10'b1011111010: data <= 20'hffdf1; 
        10'b1011111011: data <= 20'hffdc0; 
        10'b1011111100: data <= 20'h000be; 
        10'b1011111101: data <= 20'hffdda; 
        10'b1011111110: data <= 20'hffd8d; 
        10'b1011111111: data <= 20'hfffb5; 
        10'b1100000000: data <= 20'hffeaf; 
        10'b1100000001: data <= 20'hffc41; 
        10'b1100000010: data <= 20'h00015; 
        10'b1100000011: data <= 20'hffed9; 
        10'b1100000100: data <= 20'hffc9a; 
        10'b1100000101: data <= 20'hffc3b; 
        10'b1100000110: data <= 20'hffd2e; 
        10'b1100000111: data <= 20'hffc2c; 
        10'b1100001000: data <= 20'hffff2; 
        10'b1100001001: data <= 20'hffde4; 
        10'b1100001010: data <= 20'h000b4; 
        10'b1100001011: data <= 20'hffcbf; 
        10'b1100001100: data <= 20'hfff06; 
        10'b1100001101: data <= 20'hffe5e; 
        10'b1100001110: data <= 20'hffcfd; 
        10'b1100001111: data <= 20'hfff88; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 15) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 21'h1ffb91; 
        10'b0000000001: data <= 21'h1fff60; 
        10'b0000000010: data <= 21'h1fff5d; 
        10'b0000000011: data <= 21'h1ffa09; 
        10'b0000000100: data <= 21'h1ffd31; 
        10'b0000000101: data <= 21'h1ffc70; 
        10'b0000000110: data <= 21'h1ffffb; 
        10'b0000000111: data <= 21'h1ffc2a; 
        10'b0000001000: data <= 21'h1ffe6a; 
        10'b0000001001: data <= 21'h000149; 
        10'b0000001010: data <= 21'h1ffe6a; 
        10'b0000001011: data <= 21'h1ffe46; 
        10'b0000001100: data <= 21'h1ffb73; 
        10'b0000001101: data <= 21'h1fffba; 
        10'b0000001110: data <= 21'h1ff9ef; 
        10'b0000001111: data <= 21'h1ffb00; 
        10'b0000010000: data <= 21'h1ff921; 
        10'b0000010001: data <= 21'h1ffa6b; 
        10'b0000010010: data <= 21'h1fff2e; 
        10'b0000010011: data <= 21'h1ffe77; 
        10'b0000010100: data <= 21'h1ff90c; 
        10'b0000010101: data <= 21'h1ffd5c; 
        10'b0000010110: data <= 21'h1ffe16; 
        10'b0000010111: data <= 21'h1ffc93; 
        10'b0000011000: data <= 21'h1ff973; 
        10'b0000011001: data <= 21'h1ffd87; 
        10'b0000011010: data <= 21'h1ffe13; 
        10'b0000011011: data <= 21'h1ffbc1; 
        10'b0000011100: data <= 21'h1fff98; 
        10'b0000011101: data <= 21'h1ff8b6; 
        10'b0000011110: data <= 21'h1ffff3; 
        10'b0000011111: data <= 21'h1ff9bf; 
        10'b0000100000: data <= 21'h1fffbb; 
        10'b0000100001: data <= 21'h1ffbfe; 
        10'b0000100010: data <= 21'h1ffdf1; 
        10'b0000100011: data <= 21'h1ffbd3; 
        10'b0000100100: data <= 21'h1ffac5; 
        10'b0000100101: data <= 21'h1ffe16; 
        10'b0000100110: data <= 21'h0000a5; 
        10'b0000100111: data <= 21'h1ff9ea; 
        10'b0000101000: data <= 21'h1ffbc5; 
        10'b0000101001: data <= 21'h1ffa92; 
        10'b0000101010: data <= 21'h1ff902; 
        10'b0000101011: data <= 21'h1ffed5; 
        10'b0000101100: data <= 21'h1ffb43; 
        10'b0000101101: data <= 21'h1ffa76; 
        10'b0000101110: data <= 21'h1ffb67; 
        10'b0000101111: data <= 21'h1ffb18; 
        10'b0000110000: data <= 21'h1ffe72; 
        10'b0000110001: data <= 21'h1ff9a6; 
        10'b0000110010: data <= 21'h1fffe6; 
        10'b0000110011: data <= 21'h1ffa16; 
        10'b0000110100: data <= 21'h000016; 
        10'b0000110101: data <= 21'h1fff84; 
        10'b0000110110: data <= 21'h1ffa55; 
        10'b0000110111: data <= 21'h1ffcde; 
        10'b0000111000: data <= 21'h1ffcf1; 
        10'b0000111001: data <= 21'h1ffea8; 
        10'b0000111010: data <= 21'h1ffbcc; 
        10'b0000111011: data <= 21'h1ff90d; 
        10'b0000111100: data <= 21'h1ffa46; 
        10'b0000111101: data <= 21'h1ffd94; 
        10'b0000111110: data <= 21'h1fffc4; 
        10'b0000111111: data <= 21'h1ffe1d; 
        10'b0001000000: data <= 21'h1ffaf8; 
        10'b0001000001: data <= 21'h1ffc25; 
        10'b0001000010: data <= 21'h0000f6; 
        10'b0001000011: data <= 21'h1ff89b; 
        10'b0001000100: data <= 21'h1fffa7; 
        10'b0001000101: data <= 21'h1ffacb; 
        10'b0001000110: data <= 21'h1ff938; 
        10'b0001000111: data <= 21'h1ffa7b; 
        10'b0001001000: data <= 21'h1ffb93; 
        10'b0001001001: data <= 21'h1ffd70; 
        10'b0001001010: data <= 21'h1ffc28; 
        10'b0001001011: data <= 21'h1ffc36; 
        10'b0001001100: data <= 21'h0001b2; 
        10'b0001001101: data <= 21'h000030; 
        10'b0001001110: data <= 21'h0000b6; 
        10'b0001001111: data <= 21'h1ffaa4; 
        10'b0001010000: data <= 21'h1ff907; 
        10'b0001010001: data <= 21'h1ffc87; 
        10'b0001010010: data <= 21'h1fff93; 
        10'b0001010011: data <= 21'h1ffe19; 
        10'b0001010100: data <= 21'h1ffeb1; 
        10'b0001010101: data <= 21'h1ffdfe; 
        10'b0001010110: data <= 21'h1ffa58; 
        10'b0001010111: data <= 21'h1fffa3; 
        10'b0001011000: data <= 21'h1ff9c6; 
        10'b0001011001: data <= 21'h1ffbe1; 
        10'b0001011010: data <= 21'h1ff898; 
        10'b0001011011: data <= 21'h1ffb2a; 
        10'b0001011100: data <= 21'h1ff91f; 
        10'b0001011101: data <= 21'h1ffb16; 
        10'b0001011110: data <= 21'h1ff40a; 
        10'b0001011111: data <= 21'h1ff0ba; 
        10'b0001100000: data <= 21'h1ff747; 
        10'b0001100001: data <= 21'h1ff7d2; 
        10'b0001100010: data <= 21'h1ff5f3; 
        10'b0001100011: data <= 21'h1ffcac; 
        10'b0001100100: data <= 21'h1ffe8f; 
        10'b0001100101: data <= 21'h1ff81b; 
        10'b0001100110: data <= 21'h1ffb43; 
        10'b0001100111: data <= 21'h1ffe83; 
        10'b0001101000: data <= 21'h1ffeed; 
        10'b0001101001: data <= 21'h1ffcb7; 
        10'b0001101010: data <= 21'h1ff7fd; 
        10'b0001101011: data <= 21'h1ffa9f; 
        10'b0001101100: data <= 21'h1ff656; 
        10'b0001101101: data <= 21'h00011d; 
        10'b0001101110: data <= 21'h0000b2; 
        10'b0001101111: data <= 21'h1ff9af; 
        10'b0001110000: data <= 21'h1ff943; 
        10'b0001110001: data <= 21'h1ffbd3; 
        10'b0001110010: data <= 21'h0000af; 
        10'b0001110011: data <= 21'h000060; 
        10'b0001110100: data <= 21'h0000ee; 
        10'b0001110101: data <= 21'h1ffb2b; 
        10'b0001110110: data <= 21'h1ffacd; 
        10'b0001110111: data <= 21'h1ff532; 
        10'b0001111000: data <= 21'h1fedc7; 
        10'b0001111001: data <= 21'h1fe7ce; 
        10'b0001111010: data <= 21'h1fdcac; 
        10'b0001111011: data <= 21'h1fe96e; 
        10'b0001111100: data <= 21'h1fe93f; 
        10'b0001111101: data <= 21'h1fe17a; 
        10'b0001111110: data <= 21'h1fef30; 
        10'b0001111111: data <= 21'h1fffec; 
        10'b0010000000: data <= 21'h1ffe01; 
        10'b0010000001: data <= 21'h0005b1; 
        10'b0010000010: data <= 21'h1ffe46; 
        10'b0010000011: data <= 21'h1ff756; 
        10'b0010000100: data <= 21'h1ff4ab; 
        10'b0010000101: data <= 21'h1ffa02; 
        10'b0010000110: data <= 21'h1ffb17; 
        10'b0010000111: data <= 21'h1ffc90; 
        10'b0010001000: data <= 21'h1ffbbe; 
        10'b0010001001: data <= 21'h000198; 
        10'b0010001010: data <= 21'h0000e8; 
        10'b0010001011: data <= 21'h1ffce0; 
        10'b0010001100: data <= 21'h1ffd6e; 
        10'b0010001101: data <= 21'h000195; 
        10'b0010001110: data <= 21'h1ffa89; 
        10'b0010001111: data <= 21'h1ff9b9; 
        10'b0010010000: data <= 21'h1ffb5b; 
        10'b0010010001: data <= 21'h1ff4f7; 
        10'b0010010010: data <= 21'h1fef54; 
        10'b0010010011: data <= 21'h1fefe3; 
        10'b0010010100: data <= 21'h1ff572; 
        10'b0010010101: data <= 21'h1ffe07; 
        10'b0010010110: data <= 21'h00038e; 
        10'b0010010111: data <= 21'h0003d8; 
        10'b0010011000: data <= 21'h1ffa49; 
        10'b0010011001: data <= 21'h1ff7d3; 
        10'b0010011010: data <= 21'h1ffb12; 
        10'b0010011011: data <= 21'h1ffdb1; 
        10'b0010011100: data <= 21'h00082b; 
        10'b0010011101: data <= 21'h00085a; 
        10'b0010011110: data <= 21'h000fd5; 
        10'b0010011111: data <= 21'h0009dd; 
        10'b0010100000: data <= 21'h000990; 
        10'b0010100001: data <= 21'h000c46; 
        10'b0010100010: data <= 21'h0016a7; 
        10'b0010100011: data <= 21'h001345; 
        10'b0010100100: data <= 21'h000d85; 
        10'b0010100101: data <= 21'h000779; 
        10'b0010100110: data <= 21'h0004a6; 
        10'b0010100111: data <= 21'h0001bd; 
        10'b0010101000: data <= 21'h1ff9fa; 
        10'b0010101001: data <= 21'h1ff96e; 
        10'b0010101010: data <= 21'h0000d6; 
        10'b0010101011: data <= 21'h1ff9ac; 
        10'b0010101100: data <= 21'h1ff7da; 
        10'b0010101101: data <= 21'h1fec8a; 
        10'b0010101110: data <= 21'h1ff742; 
        10'b0010101111: data <= 21'h1ffefa; 
        10'b0010110000: data <= 21'h1fff50; 
        10'b0010110001: data <= 21'h0007e5; 
        10'b0010110010: data <= 21'h001064; 
        10'b0010110011: data <= 21'h000da3; 
        10'b0010110100: data <= 21'h000251; 
        10'b0010110101: data <= 21'h000506; 
        10'b0010110110: data <= 21'h1ffdbf; 
        10'b0010110111: data <= 21'h1ff83b; 
        10'b0010111000: data <= 21'h1ffb4d; 
        10'b0010111001: data <= 21'h1ffc09; 
        10'b0010111010: data <= 21'h00002d; 
        10'b0010111011: data <= 21'h000f8f; 
        10'b0010111100: data <= 21'h0008e7; 
        10'b0010111101: data <= 21'h000a1e; 
        10'b0010111110: data <= 21'h001eed; 
        10'b0010111111: data <= 21'h00252f; 
        10'b0011000000: data <= 21'h0029d4; 
        10'b0011000001: data <= 21'h001620; 
        10'b0011000010: data <= 21'h000aee; 
        10'b0011000011: data <= 21'h0002ab; 
        10'b0011000100: data <= 21'h1ffc95; 
        10'b0011000101: data <= 21'h1ffe28; 
        10'b0011000110: data <= 21'h1ffd54; 
        10'b0011000111: data <= 21'h1ff7fb; 
        10'b0011001000: data <= 21'h1fe963; 
        10'b0011001001: data <= 21'h1fe576; 
        10'b0011001010: data <= 21'h1fefd8; 
        10'b0011001011: data <= 21'h000216; 
        10'b0011001100: data <= 21'h000a95; 
        10'b0011001101: data <= 21'h0014c6; 
        10'b0011001110: data <= 21'h00143a; 
        10'b0011001111: data <= 21'h0011a9; 
        10'b0011010000: data <= 21'h00051c; 
        10'b0011010001: data <= 21'h1ffe54; 
        10'b0011010010: data <= 21'h1ffa5a; 
        10'b0011010011: data <= 21'h000062; 
        10'b0011010100: data <= 21'h0008c0; 
        10'b0011010101: data <= 21'h0007ea; 
        10'b0011010110: data <= 21'h000a05; 
        10'b0011010111: data <= 21'h001667; 
        10'b0011011000: data <= 21'h00135e; 
        10'b0011011001: data <= 21'h001729; 
        10'b0011011010: data <= 21'h002062; 
        10'b0011011011: data <= 21'h002b70; 
        10'b0011011100: data <= 21'h003507; 
        10'b0011011101: data <= 21'h002649; 
        10'b0011011110: data <= 21'h0005e6; 
        10'b0011011111: data <= 21'h1fff17; 
        10'b0011100000: data <= 21'h1ffe7d; 
        10'b0011100001: data <= 21'h000166; 
        10'b0011100010: data <= 21'h1fffe0; 
        10'b0011100011: data <= 21'h1ff513; 
        10'b0011100100: data <= 21'h1fdf6e; 
        10'b0011100101: data <= 21'h1fe427; 
        10'b0011100110: data <= 21'h1febd9; 
        10'b0011100111: data <= 21'h00013f; 
        10'b0011101000: data <= 21'h000fc0; 
        10'b0011101001: data <= 21'h0004a0; 
        10'b0011101010: data <= 21'h000877; 
        10'b0011101011: data <= 21'h00106e; 
        10'b0011101100: data <= 21'h000a05; 
        10'b0011101101: data <= 21'h1ff4ba; 
        10'b0011101110: data <= 21'h1fe748; 
        10'b0011101111: data <= 21'h1ff107; 
        10'b0011110000: data <= 21'h1ff6d0; 
        10'b0011110001: data <= 21'h0000e1; 
        10'b0011110010: data <= 21'h000285; 
        10'b0011110011: data <= 21'h0012ab; 
        10'b0011110100: data <= 21'h0013b4; 
        10'b0011110101: data <= 21'h001c12; 
        10'b0011110110: data <= 21'h002c5e; 
        10'b0011110111: data <= 21'h003a0d; 
        10'b0011111000: data <= 21'h004d72; 
        10'b0011111001: data <= 21'h003209; 
        10'b0011111010: data <= 21'h00091e; 
        10'b0011111011: data <= 21'h1fff12; 
        10'b0011111100: data <= 21'h1ff997; 
        10'b0011111101: data <= 21'h1ffc3e; 
        10'b0011111110: data <= 21'h1ff901; 
        10'b0011111111: data <= 21'h1ff0cb; 
        10'b0100000000: data <= 21'h1fee87; 
        10'b0100000001: data <= 21'h1fefdb; 
        10'b0100000010: data <= 21'h0001f7; 
        10'b0100000011: data <= 21'h1ffedf; 
        10'b0100000100: data <= 21'h000d71; 
        10'b0100000101: data <= 21'h000bad; 
        10'b0100000110: data <= 21'h000cb5; 
        10'b0100000111: data <= 21'h0021e8; 
        10'b0100001000: data <= 21'h0015de; 
        10'b0100001001: data <= 21'h1ff6ef; 
        10'b0100001010: data <= 21'h1fe234; 
        10'b0100001011: data <= 21'h1fd549; 
        10'b0100001100: data <= 21'h1fd81a; 
        10'b0100001101: data <= 21'h1fe8c8; 
        10'b0100001110: data <= 21'h1ffaad; 
        10'b0100001111: data <= 21'h1fffdb; 
        10'b0100010000: data <= 21'h001223; 
        10'b0100010001: data <= 21'h0026c8; 
        10'b0100010010: data <= 21'h003820; 
        10'b0100010011: data <= 21'h004cc5; 
        10'b0100010100: data <= 21'h00607b; 
        10'b0100010101: data <= 21'h003f64; 
        10'b0100010110: data <= 21'h000b5a; 
        10'b0100010111: data <= 21'h1ffb87; 
        10'b0100011000: data <= 21'h1ffea0; 
        10'b0100011001: data <= 21'h1ffb92; 
        10'b0100011010: data <= 21'h1ffa06; 
        10'b0100011011: data <= 21'h1ffb2f; 
        10'b0100011100: data <= 21'h1ffae8; 
        10'b0100011101: data <= 21'h1ffcb9; 
        10'b0100011110: data <= 21'h000ad3; 
        10'b0100011111: data <= 21'h00142c; 
        10'b0100100000: data <= 21'h001f7b; 
        10'b0100100001: data <= 21'h0022d7; 
        10'b0100100010: data <= 21'h00214d; 
        10'b0100100011: data <= 21'h00284e; 
        10'b0100100100: data <= 21'h002183; 
        10'b0100100101: data <= 21'h0019c1; 
        10'b0100100110: data <= 21'h1ffa7b; 
        10'b0100100111: data <= 21'h1feaf3; 
        10'b0100101000: data <= 21'h1fdcdd; 
        10'b0100101001: data <= 21'h1fddfb; 
        10'b0100101010: data <= 21'h1fdcc9; 
        10'b0100101011: data <= 21'h1fd7d9; 
        10'b0100101100: data <= 21'h1fe484; 
        10'b0100101101: data <= 21'h1ff777; 
        10'b0100101110: data <= 21'h0004ac; 
        10'b0100101111: data <= 21'h0019c3; 
        10'b0100110000: data <= 21'h003369; 
        10'b0100110001: data <= 21'h0026a4; 
        10'b0100110010: data <= 21'h000d25; 
        10'b0100110011: data <= 21'h1ffb8c; 
        10'b0100110100: data <= 21'h1ff9fb; 
        10'b0100110101: data <= 21'h00000b; 
        10'b0100110110: data <= 21'h1ffb19; 
        10'b0100110111: data <= 21'h1ffcca; 
        10'b0100111000: data <= 21'h1ffb06; 
        10'b0100111001: data <= 21'h1fff4c; 
        10'b0100111010: data <= 21'h001133; 
        10'b0100111011: data <= 21'h0014ff; 
        10'b0100111100: data <= 21'h001e5c; 
        10'b0100111101: data <= 21'h001c0a; 
        10'b0100111110: data <= 21'h001486; 
        10'b0100111111: data <= 21'h00169d; 
        10'b0101000000: data <= 21'h00256b; 
        10'b0101000001: data <= 21'h0022f2; 
        10'b0101000010: data <= 21'h00008f; 
        10'b0101000011: data <= 21'h1fea3b; 
        10'b0101000100: data <= 21'h1fe503; 
        10'b0101000101: data <= 21'h1fe2ee; 
        10'b0101000110: data <= 21'h1fd934; 
        10'b0101000111: data <= 21'h1fc9de; 
        10'b0101001000: data <= 21'h1fb169; 
        10'b0101001001: data <= 21'h1fb7d9; 
        10'b0101001010: data <= 21'h1fc4df; 
        10'b0101001011: data <= 21'h1fd4e2; 
        10'b0101001100: data <= 21'h1ff0a8; 
        10'b0101001101: data <= 21'h0001b0; 
        10'b0101001110: data <= 21'h000453; 
        10'b0101001111: data <= 21'h1ffd62; 
        10'b0101010000: data <= 21'h1ffd4e; 
        10'b0101010001: data <= 21'h1ffdc7; 
        10'b0101010010: data <= 21'h1ffcc2; 
        10'b0101010011: data <= 21'h1ffb79; 
        10'b0101010100: data <= 21'h1ffc90; 
        10'b0101010101: data <= 21'h0008b6; 
        10'b0101010110: data <= 21'h0013bd; 
        10'b0101010111: data <= 21'h00119c; 
        10'b0101011000: data <= 21'h000cf2; 
        10'b0101011001: data <= 21'h00076a; 
        10'b0101011010: data <= 21'h0015de; 
        10'b0101011011: data <= 21'h002d45; 
        10'b0101011100: data <= 21'h002a49; 
        10'b0101011101: data <= 21'h002b59; 
        10'b0101011110: data <= 21'h000478; 
        10'b0101011111: data <= 21'h1fea04; 
        10'b0101100000: data <= 21'h1fd71c; 
        10'b0101100001: data <= 21'h1fdee7; 
        10'b0101100010: data <= 21'h1fe98a; 
        10'b0101100011: data <= 21'h1fdfc1; 
        10'b0101100100: data <= 21'h1fdb44; 
        10'b0101100101: data <= 21'h1fc305; 
        10'b0101100110: data <= 21'h1fba6e; 
        10'b0101100111: data <= 21'h1fc38e; 
        10'b0101101000: data <= 21'h1fd795; 
        10'b0101101001: data <= 21'h1ff486; 
        10'b0101101010: data <= 21'h000099; 
        10'b0101101011: data <= 21'h1ffff6; 
        10'b0101101100: data <= 21'h1ffd99; 
        10'b0101101101: data <= 21'h1ffa48; 
        10'b0101101110: data <= 21'h1ff9e9; 
        10'b0101101111: data <= 21'h1ffbc1; 
        10'b0101110000: data <= 21'h1ffeb5; 
        10'b0101110001: data <= 21'h000490; 
        10'b0101110010: data <= 21'h000d39; 
        10'b0101110011: data <= 21'h0009b2; 
        10'b0101110100: data <= 21'h000b35; 
        10'b0101110101: data <= 21'h000942; 
        10'b0101110110: data <= 21'h001e74; 
        10'b0101110111: data <= 21'h002207; 
        10'b0101111000: data <= 21'h001950; 
        10'b0101111001: data <= 21'h0017a5; 
        10'b0101111010: data <= 21'h1ffb40; 
        10'b0101111011: data <= 21'h1fe5d3; 
        10'b0101111100: data <= 21'h1fd567; 
        10'b0101111101: data <= 21'h1fe97e; 
        10'b0101111110: data <= 21'h1ff802; 
        10'b0101111111: data <= 21'h1ff6c0; 
        10'b0110000000: data <= 21'h1ffb98; 
        10'b0110000001: data <= 21'h1feeba; 
        10'b0110000010: data <= 21'h1fe0c5; 
        10'b0110000011: data <= 21'h1fd25d; 
        10'b0110000100: data <= 21'h1fdda1; 
        10'b0110000101: data <= 21'h1ffa09; 
        10'b0110000110: data <= 21'h1ff982; 
        10'b0110000111: data <= 21'h1fff0d; 
        10'b0110001000: data <= 21'h1ffdb1; 
        10'b0110001001: data <= 21'h1ff9cf; 
        10'b0110001010: data <= 21'h1ffcf1; 
        10'b0110001011: data <= 21'h1ff855; 
        10'b0110001100: data <= 21'h1ffd6d; 
        10'b0110001101: data <= 21'h1ffd38; 
        10'b0110001110: data <= 21'h1fffdc; 
        10'b0110001111: data <= 21'h1ffe89; 
        10'b0110010000: data <= 21'h000dff; 
        10'b0110010001: data <= 21'h001624; 
        10'b0110010010: data <= 21'h001a91; 
        10'b0110010011: data <= 21'h000516; 
        10'b0110010100: data <= 21'h0008fd; 
        10'b0110010101: data <= 21'h1ffe56; 
        10'b0110010110: data <= 21'h1fecfe; 
        10'b0110010111: data <= 21'h1fea1c; 
        10'b0110011000: data <= 21'h1fe19e; 
        10'b0110011001: data <= 21'h1fe524; 
        10'b0110011010: data <= 21'h1fe6d6; 
        10'b0110011011: data <= 21'h1ff3dd; 
        10'b0110011100: data <= 21'h1ff57f; 
        10'b0110011101: data <= 21'h1ff676; 
        10'b0110011110: data <= 21'h1ffa37; 
        10'b0110011111: data <= 21'h1fe6ee; 
        10'b0110100000: data <= 21'h1fef20; 
        10'b0110100001: data <= 21'h1ff78b; 
        10'b0110100010: data <= 21'h1ffcfe; 
        10'b0110100011: data <= 21'h1ff884; 
        10'b0110100100: data <= 21'h1ff94a; 
        10'b0110100101: data <= 21'h000108; 
        10'b0110100110: data <= 21'h1ff8c7; 
        10'b0110100111: data <= 21'h1ffd0c; 
        10'b0110101000: data <= 21'h1ff547; 
        10'b0110101001: data <= 21'h1fefe4; 
        10'b0110101010: data <= 21'h1fe974; 
        10'b0110101011: data <= 21'h1ff110; 
        10'b0110101100: data <= 21'h00056f; 
        10'b0110101101: data <= 21'h0018f0; 
        10'b0110101110: data <= 21'h000bd8; 
        10'b0110101111: data <= 21'h000aeb; 
        10'b0110110000: data <= 21'h00096a; 
        10'b0110110001: data <= 21'h1ff77d; 
        10'b0110110010: data <= 21'h1fe3ca; 
        10'b0110110011: data <= 21'h1fdf8d; 
        10'b0110110100: data <= 21'h1fe2b7; 
        10'b0110110101: data <= 21'h1fe1fd; 
        10'b0110110110: data <= 21'h1feade; 
        10'b0110110111: data <= 21'h1ffeee; 
        10'b0110111000: data <= 21'h1ff8d2; 
        10'b0110111001: data <= 21'h1ff9f0; 
        10'b0110111010: data <= 21'h1ff8be; 
        10'b0110111011: data <= 21'h1ff7a8; 
        10'b0110111100: data <= 21'h1ffa26; 
        10'b0110111101: data <= 21'h1fffd2; 
        10'b0110111110: data <= 21'h000129; 
        10'b0110111111: data <= 21'h1ffb82; 
        10'b0111000000: data <= 21'h1ffbf7; 
        10'b0111000001: data <= 21'h1ffd61; 
        10'b0111000010: data <= 21'h1ffe40; 
        10'b0111000011: data <= 21'h1ff8cc; 
        10'b0111000100: data <= 21'h1ffbce; 
        10'b0111000101: data <= 21'h1fedae; 
        10'b0111000110: data <= 21'h1fdb4d; 
        10'b0111000111: data <= 21'h1fd499; 
        10'b0111001000: data <= 21'h1fe2a5; 
        10'b0111001001: data <= 21'h1fefc3; 
        10'b0111001010: data <= 21'h1ff98e; 
        10'b0111001011: data <= 21'h1ff6bb; 
        10'b0111001100: data <= 21'h1ff9f4; 
        10'b0111001101: data <= 21'h1febff; 
        10'b0111001110: data <= 21'h1fd979; 
        10'b0111001111: data <= 21'h1fe0b8; 
        10'b0111010000: data <= 21'h1fe946; 
        10'b0111010001: data <= 21'h1ff7d0; 
        10'b0111010010: data <= 21'h1ff84c; 
        10'b0111010011: data <= 21'h00013f; 
        10'b0111010100: data <= 21'h000655; 
        10'b0111010101: data <= 21'h000101; 
        10'b0111010110: data <= 21'h0006e1; 
        10'b0111010111: data <= 21'h000191; 
        10'b0111011000: data <= 21'h000113; 
        10'b0111011001: data <= 21'h0000f8; 
        10'b0111011010: data <= 21'h1ffbb0; 
        10'b0111011011: data <= 21'h1ffc05; 
        10'b0111011100: data <= 21'h1ffb38; 
        10'b0111011101: data <= 21'h1fffae; 
        10'b0111011110: data <= 21'h1ffffa; 
        10'b0111011111: data <= 21'h000087; 
        10'b0111100000: data <= 21'h1ffb5a; 
        10'b0111100001: data <= 21'h000157; 
        10'b0111100010: data <= 21'h0002ae; 
        10'b0111100011: data <= 21'h1fe356; 
        10'b0111100100: data <= 21'h1fcc26; 
        10'b0111100101: data <= 21'h1fcf7a; 
        10'b0111100110: data <= 21'h1fdd3c; 
        10'b0111100111: data <= 21'h1feb16; 
        10'b0111101000: data <= 21'h1fdf4e; 
        10'b0111101001: data <= 21'h1fd5cf; 
        10'b0111101010: data <= 21'h1fd6fb; 
        10'b0111101011: data <= 21'h1fed52; 
        10'b0111101100: data <= 21'h1ff7cb; 
        10'b0111101101: data <= 21'h000c66; 
        10'b0111101110: data <= 21'h0012f5; 
        10'b0111101111: data <= 21'h000c63; 
        10'b0111110000: data <= 21'h000c7f; 
        10'b0111110001: data <= 21'h0003a2; 
        10'b0111110010: data <= 21'h000068; 
        10'b0111110011: data <= 21'h0006e7; 
        10'b0111110100: data <= 21'h000704; 
        10'b0111110101: data <= 21'h1ffa15; 
        10'b0111110110: data <= 21'h1fffc2; 
        10'b0111110111: data <= 21'h00002a; 
        10'b0111111000: data <= 21'h0000b2; 
        10'b0111111001: data <= 21'h1ffaf7; 
        10'b0111111010: data <= 21'h1ffcd2; 
        10'b0111111011: data <= 21'h1ffbe9; 
        10'b0111111100: data <= 21'h000a42; 
        10'b0111111101: data <= 21'h000d8e; 
        10'b0111111110: data <= 21'h002035; 
        10'b0111111111: data <= 21'h0005aa; 
        10'b1000000000: data <= 21'h1fe0fd; 
        10'b1000000001: data <= 21'h1fd2de; 
        10'b1000000010: data <= 21'h1fc49c; 
        10'b1000000011: data <= 21'h1fcaf4; 
        10'b1000000100: data <= 21'h1fd9f5; 
        10'b1000000101: data <= 21'h1fea47; 
        10'b1000000110: data <= 21'h1ff528; 
        10'b1000000111: data <= 21'h1ffb76; 
        10'b1000001000: data <= 21'h1fff2f; 
        10'b1000001001: data <= 21'h000e8f; 
        10'b1000001010: data <= 21'h000752; 
        10'b1000001011: data <= 21'h000cfc; 
        10'b1000001100: data <= 21'h0008ba; 
        10'b1000001101: data <= 21'h000caa; 
        10'b1000001110: data <= 21'h000a6f; 
        10'b1000001111: data <= 21'h000e6d; 
        10'b1000010000: data <= 21'h00077f; 
        10'b1000010001: data <= 21'h00008f; 
        10'b1000010010: data <= 21'h1ffa84; 
        10'b1000010011: data <= 21'h1ffe3d; 
        10'b1000010100: data <= 21'h000009; 
        10'b1000010101: data <= 21'h1ffaed; 
        10'b1000010110: data <= 21'h1ffd47; 
        10'b1000010111: data <= 21'h000117; 
        10'b1000011000: data <= 21'h000f92; 
        10'b1000011001: data <= 21'h001a9a; 
        10'b1000011010: data <= 21'h0023d1; 
        10'b1000011011: data <= 21'h00181c; 
        10'b1000011100: data <= 21'h000f45; 
        10'b1000011101: data <= 21'h0004f5; 
        10'b1000011110: data <= 21'h1ff499; 
        10'b1000011111: data <= 21'h1ff3d4; 
        10'b1000100000: data <= 21'h000108; 
        10'b1000100001: data <= 21'h000e98; 
        10'b1000100010: data <= 21'h000574; 
        10'b1000100011: data <= 21'h0007c0; 
        10'b1000100100: data <= 21'h0007de; 
        10'b1000100101: data <= 21'h1ffd85; 
        10'b1000100110: data <= 21'h0005a6; 
        10'b1000100111: data <= 21'h000585; 
        10'b1000101000: data <= 21'h00012d; 
        10'b1000101001: data <= 21'h000975; 
        10'b1000101010: data <= 21'h00103e; 
        10'b1000101011: data <= 21'h000be0; 
        10'b1000101100: data <= 21'h0000fd; 
        10'b1000101101: data <= 21'h1fffce; 
        10'b1000101110: data <= 21'h1ffff2; 
        10'b1000101111: data <= 21'h1ff99e; 
        10'b1000110000: data <= 21'h1fffad; 
        10'b1000110001: data <= 21'h1ff88e; 
        10'b1000110010: data <= 21'h1ffc74; 
        10'b1000110011: data <= 21'h1ffa71; 
        10'b1000110100: data <= 21'h000216; 
        10'b1000110101: data <= 21'h00117f; 
        10'b1000110110: data <= 21'h001451; 
        10'b1000110111: data <= 21'h0018c1; 
        10'b1000111000: data <= 21'h0022b0; 
        10'b1000111001: data <= 21'h001d4b; 
        10'b1000111010: data <= 21'h0019bd; 
        10'b1000111011: data <= 21'h002584; 
        10'b1000111100: data <= 21'h00175b; 
        10'b1000111101: data <= 21'h001184; 
        10'b1000111110: data <= 21'h1ffb11; 
        10'b1000111111: data <= 21'h1ffb78; 
        10'b1001000000: data <= 21'h000ce8; 
        10'b1001000001: data <= 21'h00069a; 
        10'b1001000010: data <= 21'h000ac8; 
        10'b1001000011: data <= 21'h000e45; 
        10'b1001000100: data <= 21'h000c7f; 
        10'b1001000101: data <= 21'h0009d0; 
        10'b1001000110: data <= 21'h001778; 
        10'b1001000111: data <= 21'h00118a; 
        10'b1001001000: data <= 21'h1ffdb7; 
        10'b1001001001: data <= 21'h1ff8b4; 
        10'b1001001010: data <= 21'h1ffd6c; 
        10'b1001001011: data <= 21'h1ffb5f; 
        10'b1001001100: data <= 21'h1ffab2; 
        10'b1001001101: data <= 21'h00002b; 
        10'b1001001110: data <= 21'h1ff842; 
        10'b1001001111: data <= 21'h1ffd18; 
        10'b1001010000: data <= 21'h0006e7; 
        10'b1001010001: data <= 21'h1ffdcb; 
        10'b1001010010: data <= 21'h00085e; 
        10'b1001010011: data <= 21'h0016a4; 
        10'b1001010100: data <= 21'h0020b1; 
        10'b1001010101: data <= 21'h001562; 
        10'b1001010110: data <= 21'h001223; 
        10'b1001010111: data <= 21'h0009c7; 
        10'b1001011000: data <= 21'h000ca7; 
        10'b1001011001: data <= 21'h0007dc; 
        10'b1001011010: data <= 21'h00082f; 
        10'b1001011011: data <= 21'h0009fa; 
        10'b1001011100: data <= 21'h000298; 
        10'b1001011101: data <= 21'h00080a; 
        10'b1001011110: data <= 21'h00041e; 
        10'b1001011111: data <= 21'h000cf5; 
        10'b1001100000: data <= 21'h000cb9; 
        10'b1001100001: data <= 21'h001557; 
        10'b1001100010: data <= 21'h001a3f; 
        10'b1001100011: data <= 21'h0005ac; 
        10'b1001100100: data <= 21'h000039; 
        10'b1001100101: data <= 21'h1ff9c4; 
        10'b1001100110: data <= 21'h1ffb73; 
        10'b1001100111: data <= 21'h1ffb79; 
        10'b1001101000: data <= 21'h1ffe76; 
        10'b1001101001: data <= 21'h1ff8e8; 
        10'b1001101010: data <= 21'h1ffc51; 
        10'b1001101011: data <= 21'h1ffb73; 
        10'b1001101100: data <= 21'h00027e; 
        10'b1001101101: data <= 21'h1ffc81; 
        10'b1001101110: data <= 21'h1ff857; 
        10'b1001101111: data <= 21'h1ffea2; 
        10'b1001110000: data <= 21'h000cb5; 
        10'b1001110001: data <= 21'h001294; 
        10'b1001110010: data <= 21'h000339; 
        10'b1001110011: data <= 21'h001072; 
        10'b1001110100: data <= 21'h001a99; 
        10'b1001110101: data <= 21'h0020d8; 
        10'b1001110110: data <= 21'h0010b8; 
        10'b1001110111: data <= 21'h000286; 
        10'b1001111000: data <= 21'h0001d8; 
        10'b1001111001: data <= 21'h00041a; 
        10'b1001111010: data <= 21'h00089b; 
        10'b1001111011: data <= 21'h000890; 
        10'b1001111100: data <= 21'h000eac; 
        10'b1001111101: data <= 21'h000d41; 
        10'b1001111110: data <= 21'h000dd7; 
        10'b1001111111: data <= 21'h0004de; 
        10'b1010000000: data <= 21'h1fff4a; 
        10'b1010000001: data <= 21'h0000c6; 
        10'b1010000010: data <= 21'h1ffd52; 
        10'b1010000011: data <= 21'h1ffe35; 
        10'b1010000100: data <= 21'h1ffa28; 
        10'b1010000101: data <= 21'h1ffd26; 
        10'b1010000110: data <= 21'h1ffe59; 
        10'b1010000111: data <= 21'h1ffdb8; 
        10'b1010001000: data <= 21'h1ffa74; 
        10'b1010001001: data <= 21'h1ffc57; 
        10'b1010001010: data <= 21'h1ff4e1; 
        10'b1010001011: data <= 21'h1ffaf1; 
        10'b1010001100: data <= 21'h000a10; 
        10'b1010001101: data <= 21'h0009da; 
        10'b1010001110: data <= 21'h0009d5; 
        10'b1010001111: data <= 21'h001188; 
        10'b1010010000: data <= 21'h0010d3; 
        10'b1010010001: data <= 21'h000b85; 
        10'b1010010010: data <= 21'h000d3d; 
        10'b1010010011: data <= 21'h000c1f; 
        10'b1010010100: data <= 21'h000bdc; 
        10'b1010010101: data <= 21'h000574; 
        10'b1010010110: data <= 21'h1ff9bd; 
        10'b1010010111: data <= 21'h1fff20; 
        10'b1010011000: data <= 21'h0005d0; 
        10'b1010011001: data <= 21'h00025c; 
        10'b1010011010: data <= 21'h0007ca; 
        10'b1010011011: data <= 21'h1ffb20; 
        10'b1010011100: data <= 21'h00014e; 
        10'b1010011101: data <= 21'h1ffc03; 
        10'b1010011110: data <= 21'h1ffbec; 
        10'b1010011111: data <= 21'h000138; 
        10'b1010100000: data <= 21'h1fff71; 
        10'b1010100001: data <= 21'h1ffc2b; 
        10'b1010100010: data <= 21'h1ffb96; 
        10'b1010100011: data <= 21'h00015d; 
        10'b1010100100: data <= 21'h1ff863; 
        10'b1010100101: data <= 21'h1ff7ea; 
        10'b1010100110: data <= 21'h1ffd18; 
        10'b1010100111: data <= 21'h1ffe86; 
        10'b1010101000: data <= 21'h1fff8c; 
        10'b1010101001: data <= 21'h000d05; 
        10'b1010101010: data <= 21'h0010e6; 
        10'b1010101011: data <= 21'h000d02; 
        10'b1010101100: data <= 21'h000872; 
        10'b1010101101: data <= 21'h000bc2; 
        10'b1010101110: data <= 21'h0015b0; 
        10'b1010101111: data <= 21'h0011f1; 
        10'b1010110000: data <= 21'h000ab4; 
        10'b1010110001: data <= 21'h000534; 
        10'b1010110010: data <= 21'h0009f0; 
        10'b1010110011: data <= 21'h000671; 
        10'b1010110100: data <= 21'h1fffa1; 
        10'b1010110101: data <= 21'h1fff12; 
        10'b1010110110: data <= 21'h1ffda4; 
        10'b1010110111: data <= 21'h000068; 
        10'b1010111000: data <= 21'h1ffac2; 
        10'b1010111001: data <= 21'h1ffe1e; 
        10'b1010111010: data <= 21'h0000c9; 
        10'b1010111011: data <= 21'h1ff997; 
        10'b1010111100: data <= 21'h1ffd22; 
        10'b1010111101: data <= 21'h000045; 
        10'b1010111110: data <= 21'h0000c1; 
        10'b1010111111: data <= 21'h1ff946; 
        10'b1011000000: data <= 21'h1ffff4; 
        10'b1011000001: data <= 21'h1ffdeb; 
        10'b1011000010: data <= 21'h1ff803; 
        10'b1011000011: data <= 21'h1ffd0d; 
        10'b1011000100: data <= 21'h1ff8d4; 
        10'b1011000101: data <= 21'h00043b; 
        10'b1011000110: data <= 21'h000327; 
        10'b1011000111: data <= 21'h0008cd; 
        10'b1011001000: data <= 21'h0008c1; 
        10'b1011001001: data <= 21'h000f5a; 
        10'b1011001010: data <= 21'h0000d8; 
        10'b1011001011: data <= 21'h000492; 
        10'b1011001100: data <= 21'h0003dd; 
        10'b1011001101: data <= 21'h000784; 
        10'b1011001110: data <= 21'h1ffaf7; 
        10'b1011001111: data <= 21'h1fffc8; 
        10'b1011010000: data <= 21'h1ff79d; 
        10'b1011010001: data <= 21'h0000b8; 
        10'b1011010010: data <= 21'h1ffcdf; 
        10'b1011010011: data <= 21'h1ffa5f; 
        10'b1011010100: data <= 21'h1fff56; 
        10'b1011010101: data <= 21'h000062; 
        10'b1011010110: data <= 21'h1ff8db; 
        10'b1011010111: data <= 21'h1ffc3a; 
        10'b1011011000: data <= 21'h1ffdc4; 
        10'b1011011001: data <= 21'h1ffd8a; 
        10'b1011011010: data <= 21'h1ffac0; 
        10'b1011011011: data <= 21'h1ffc05; 
        10'b1011011100: data <= 21'h1ffb93; 
        10'b1011011101: data <= 21'h1ffc5e; 
        10'b1011011110: data <= 21'h1ffeb2; 
        10'b1011011111: data <= 21'h1ffacb; 
        10'b1011100000: data <= 21'h1ff920; 
        10'b1011100001: data <= 21'h1ffc6d; 
        10'b1011100010: data <= 21'h1ffb4e; 
        10'b1011100011: data <= 21'h1fff1c; 
        10'b1011100100: data <= 21'h000024; 
        10'b1011100101: data <= 21'h1ffe33; 
        10'b1011100110: data <= 21'h1ffafd; 
        10'b1011100111: data <= 21'h1ffd70; 
        10'b1011101000: data <= 21'h1ffeda; 
        10'b1011101001: data <= 21'h1ffac4; 
        10'b1011101010: data <= 21'h1ff5e4; 
        10'b1011101011: data <= 21'h1ff7d1; 
        10'b1011101100: data <= 21'h1ffe45; 
        10'b1011101101: data <= 21'h1ffe3b; 
        10'b1011101110: data <= 21'h1ffb63; 
        10'b1011101111: data <= 21'h1ffea6; 
        10'b1011110000: data <= 21'h1ffc90; 
        10'b1011110001: data <= 21'h1ffda6; 
        10'b1011110010: data <= 21'h1ffbbf; 
        10'b1011110011: data <= 21'h1ff8d9; 
        10'b1011110100: data <= 21'h1ffe6c; 
        10'b1011110101: data <= 21'h1fff08; 
        10'b1011110110: data <= 21'h1fff52; 
        10'b1011110111: data <= 21'h1ffdfd; 
        10'b1011111000: data <= 21'h1ff9e4; 
        10'b1011111001: data <= 21'h1fff9e; 
        10'b1011111010: data <= 21'h1ffbe3; 
        10'b1011111011: data <= 21'h1ffb7f; 
        10'b1011111100: data <= 21'h00017c; 
        10'b1011111101: data <= 21'h1ffbb4; 
        10'b1011111110: data <= 21'h1ffb1a; 
        10'b1011111111: data <= 21'h1fff6b; 
        10'b1100000000: data <= 21'h1ffd5e; 
        10'b1100000001: data <= 21'h1ff881; 
        10'b1100000010: data <= 21'h00002a; 
        10'b1100000011: data <= 21'h1ffdb2; 
        10'b1100000100: data <= 21'h1ff933; 
        10'b1100000101: data <= 21'h1ff876; 
        10'b1100000110: data <= 21'h1ffa5c; 
        10'b1100000111: data <= 21'h1ff859; 
        10'b1100001000: data <= 21'h1fffe4; 
        10'b1100001001: data <= 21'h1ffbc8; 
        10'b1100001010: data <= 21'h000168; 
        10'b1100001011: data <= 21'h1ff97e; 
        10'b1100001100: data <= 21'h1ffe0b; 
        10'b1100001101: data <= 21'h1ffcbc; 
        10'b1100001110: data <= 21'h1ff9fa; 
        10'b1100001111: data <= 21'h1fff0f; 
      endcase 
    end 
  end 
endgenerate 
generate 
  if (WGHT_FRC == 16) begin  
    always @(posedge clk) 
      begin 
        case(address) 
        10'b0000000000: data <= 22'h3ff722; 
        10'b0000000001: data <= 22'h3ffebf; 
        10'b0000000010: data <= 22'h3ffeb9; 
        10'b0000000011: data <= 22'h3ff412; 
        10'b0000000100: data <= 22'h3ffa62; 
        10'b0000000101: data <= 22'h3ff8e0; 
        10'b0000000110: data <= 22'h3ffff6; 
        10'b0000000111: data <= 22'h3ff854; 
        10'b0000001000: data <= 22'h3ffcd5; 
        10'b0000001001: data <= 22'h000292; 
        10'b0000001010: data <= 22'h3ffcd4; 
        10'b0000001011: data <= 22'h3ffc8b; 
        10'b0000001100: data <= 22'h3ff6e7; 
        10'b0000001101: data <= 22'h3fff73; 
        10'b0000001110: data <= 22'h3ff3de; 
        10'b0000001111: data <= 22'h3ff600; 
        10'b0000010000: data <= 22'h3ff242; 
        10'b0000010001: data <= 22'h3ff4d6; 
        10'b0000010010: data <= 22'h3ffe5c; 
        10'b0000010011: data <= 22'h3ffcee; 
        10'b0000010100: data <= 22'h3ff218; 
        10'b0000010101: data <= 22'h3ffab8; 
        10'b0000010110: data <= 22'h3ffc2b; 
        10'b0000010111: data <= 22'h3ff927; 
        10'b0000011000: data <= 22'h3ff2e7; 
        10'b0000011001: data <= 22'h3ffb0e; 
        10'b0000011010: data <= 22'h3ffc27; 
        10'b0000011011: data <= 22'h3ff782; 
        10'b0000011100: data <= 22'h3fff30; 
        10'b0000011101: data <= 22'h3ff16c; 
        10'b0000011110: data <= 22'h3fffe7; 
        10'b0000011111: data <= 22'h3ff37d; 
        10'b0000100000: data <= 22'h3fff76; 
        10'b0000100001: data <= 22'h3ff7fb; 
        10'b0000100010: data <= 22'h3ffbe1; 
        10'b0000100011: data <= 22'h3ff7a6; 
        10'b0000100100: data <= 22'h3ff58a; 
        10'b0000100101: data <= 22'h3ffc2c; 
        10'b0000100110: data <= 22'h000149; 
        10'b0000100111: data <= 22'h3ff3d3; 
        10'b0000101000: data <= 22'h3ff78a; 
        10'b0000101001: data <= 22'h3ff525; 
        10'b0000101010: data <= 22'h3ff203; 
        10'b0000101011: data <= 22'h3ffdaa; 
        10'b0000101100: data <= 22'h3ff686; 
        10'b0000101101: data <= 22'h3ff4ec; 
        10'b0000101110: data <= 22'h3ff6ce; 
        10'b0000101111: data <= 22'h3ff62f; 
        10'b0000110000: data <= 22'h3ffce5; 
        10'b0000110001: data <= 22'h3ff34c; 
        10'b0000110010: data <= 22'h3fffcc; 
        10'b0000110011: data <= 22'h3ff42c; 
        10'b0000110100: data <= 22'h00002b; 
        10'b0000110101: data <= 22'h3fff09; 
        10'b0000110110: data <= 22'h3ff4aa; 
        10'b0000110111: data <= 22'h3ff9bc; 
        10'b0000111000: data <= 22'h3ff9e2; 
        10'b0000111001: data <= 22'h3ffd50; 
        10'b0000111010: data <= 22'h3ff798; 
        10'b0000111011: data <= 22'h3ff21a; 
        10'b0000111100: data <= 22'h3ff48c; 
        10'b0000111101: data <= 22'h3ffb27; 
        10'b0000111110: data <= 22'h3fff87; 
        10'b0000111111: data <= 22'h3ffc3b; 
        10'b0001000000: data <= 22'h3ff5f0; 
        10'b0001000001: data <= 22'h3ff84a; 
        10'b0001000010: data <= 22'h0001ec; 
        10'b0001000011: data <= 22'h3ff136; 
        10'b0001000100: data <= 22'h3fff4f; 
        10'b0001000101: data <= 22'h3ff597; 
        10'b0001000110: data <= 22'h3ff26f; 
        10'b0001000111: data <= 22'h3ff4f5; 
        10'b0001001000: data <= 22'h3ff725; 
        10'b0001001001: data <= 22'h3ffae0; 
        10'b0001001010: data <= 22'h3ff850; 
        10'b0001001011: data <= 22'h3ff86c; 
        10'b0001001100: data <= 22'h000365; 
        10'b0001001101: data <= 22'h000060; 
        10'b0001001110: data <= 22'h00016d; 
        10'b0001001111: data <= 22'h3ff548; 
        10'b0001010000: data <= 22'h3ff20e; 
        10'b0001010001: data <= 22'h3ff90f; 
        10'b0001010010: data <= 22'h3fff26; 
        10'b0001010011: data <= 22'h3ffc33; 
        10'b0001010100: data <= 22'h3ffd61; 
        10'b0001010101: data <= 22'h3ffbfc; 
        10'b0001010110: data <= 22'h3ff4b1; 
        10'b0001010111: data <= 22'h3fff46; 
        10'b0001011000: data <= 22'h3ff38b; 
        10'b0001011001: data <= 22'h3ff7c2; 
        10'b0001011010: data <= 22'h3ff130; 
        10'b0001011011: data <= 22'h3ff655; 
        10'b0001011100: data <= 22'h3ff23f; 
        10'b0001011101: data <= 22'h3ff62b; 
        10'b0001011110: data <= 22'h3fe814; 
        10'b0001011111: data <= 22'h3fe173; 
        10'b0001100000: data <= 22'h3fee8e; 
        10'b0001100001: data <= 22'h3fefa3; 
        10'b0001100010: data <= 22'h3febe6; 
        10'b0001100011: data <= 22'h3ff958; 
        10'b0001100100: data <= 22'h3ffd1f; 
        10'b0001100101: data <= 22'h3ff037; 
        10'b0001100110: data <= 22'h3ff686; 
        10'b0001100111: data <= 22'h3ffd05; 
        10'b0001101000: data <= 22'h3ffdd9; 
        10'b0001101001: data <= 22'h3ff96f; 
        10'b0001101010: data <= 22'h3feffb; 
        10'b0001101011: data <= 22'h3ff53d; 
        10'b0001101100: data <= 22'h3fecac; 
        10'b0001101101: data <= 22'h000239; 
        10'b0001101110: data <= 22'h000164; 
        10'b0001101111: data <= 22'h3ff35d; 
        10'b0001110000: data <= 22'h3ff287; 
        10'b0001110001: data <= 22'h3ff7a6; 
        10'b0001110010: data <= 22'h00015e; 
        10'b0001110011: data <= 22'h0000c0; 
        10'b0001110100: data <= 22'h0001dd; 
        10'b0001110101: data <= 22'h3ff656; 
        10'b0001110110: data <= 22'h3ff599; 
        10'b0001110111: data <= 22'h3fea64; 
        10'b0001111000: data <= 22'h3fdb8e; 
        10'b0001111001: data <= 22'h3fcf9b; 
        10'b0001111010: data <= 22'h3fb958; 
        10'b0001111011: data <= 22'h3fd2dc; 
        10'b0001111100: data <= 22'h3fd27e; 
        10'b0001111101: data <= 22'h3fc2f5; 
        10'b0001111110: data <= 22'h3fde61; 
        10'b0001111111: data <= 22'h3fffd8; 
        10'b0010000000: data <= 22'h3ffc02; 
        10'b0010000001: data <= 22'h000b63; 
        10'b0010000010: data <= 22'h3ffc8b; 
        10'b0010000011: data <= 22'h3feeab; 
        10'b0010000100: data <= 22'h3fe956; 
        10'b0010000101: data <= 22'h3ff404; 
        10'b0010000110: data <= 22'h3ff62e; 
        10'b0010000111: data <= 22'h3ff91f; 
        10'b0010001000: data <= 22'h3ff77c; 
        10'b0010001001: data <= 22'h000330; 
        10'b0010001010: data <= 22'h0001d0; 
        10'b0010001011: data <= 22'h3ff9bf; 
        10'b0010001100: data <= 22'h3ffadc; 
        10'b0010001101: data <= 22'h000329; 
        10'b0010001110: data <= 22'h3ff513; 
        10'b0010001111: data <= 22'h3ff371; 
        10'b0010010000: data <= 22'h3ff6b5; 
        10'b0010010001: data <= 22'h3fe9ed; 
        10'b0010010010: data <= 22'h3fdea8; 
        10'b0010010011: data <= 22'h3fdfc7; 
        10'b0010010100: data <= 22'h3feae3; 
        10'b0010010101: data <= 22'h3ffc0d; 
        10'b0010010110: data <= 22'h00071d; 
        10'b0010010111: data <= 22'h0007b0; 
        10'b0010011000: data <= 22'h3ff491; 
        10'b0010011001: data <= 22'h3fefa7; 
        10'b0010011010: data <= 22'h3ff623; 
        10'b0010011011: data <= 22'h3ffb62; 
        10'b0010011100: data <= 22'h001057; 
        10'b0010011101: data <= 22'h0010b4; 
        10'b0010011110: data <= 22'h001faa; 
        10'b0010011111: data <= 22'h0013ba; 
        10'b0010100000: data <= 22'h001321; 
        10'b0010100001: data <= 22'h00188d; 
        10'b0010100010: data <= 22'h002d4e; 
        10'b0010100011: data <= 22'h002689; 
        10'b0010100100: data <= 22'h001b0a; 
        10'b0010100101: data <= 22'h000ef3; 
        10'b0010100110: data <= 22'h00094d; 
        10'b0010100111: data <= 22'h00037a; 
        10'b0010101000: data <= 22'h3ff3f5; 
        10'b0010101001: data <= 22'h3ff2dd; 
        10'b0010101010: data <= 22'h0001ac; 
        10'b0010101011: data <= 22'h3ff359; 
        10'b0010101100: data <= 22'h3fefb5; 
        10'b0010101101: data <= 22'h3fd915; 
        10'b0010101110: data <= 22'h3fee84; 
        10'b0010101111: data <= 22'h3ffdf4; 
        10'b0010110000: data <= 22'h3ffea0; 
        10'b0010110001: data <= 22'h000fca; 
        10'b0010110010: data <= 22'h0020c8; 
        10'b0010110011: data <= 22'h001b46; 
        10'b0010110100: data <= 22'h0004a2; 
        10'b0010110101: data <= 22'h000a0b; 
        10'b0010110110: data <= 22'h3ffb7e; 
        10'b0010110111: data <= 22'h3ff077; 
        10'b0010111000: data <= 22'h3ff69a; 
        10'b0010111001: data <= 22'h3ff812; 
        10'b0010111010: data <= 22'h00005b; 
        10'b0010111011: data <= 22'h001f1f; 
        10'b0010111100: data <= 22'h0011cf; 
        10'b0010111101: data <= 22'h00143c; 
        10'b0010111110: data <= 22'h003dda; 
        10'b0010111111: data <= 22'h004a5e; 
        10'b0011000000: data <= 22'h0053a8; 
        10'b0011000001: data <= 22'h002c40; 
        10'b0011000010: data <= 22'h0015db; 
        10'b0011000011: data <= 22'h000557; 
        10'b0011000100: data <= 22'h3ff92a; 
        10'b0011000101: data <= 22'h3ffc50; 
        10'b0011000110: data <= 22'h3ffaa8; 
        10'b0011000111: data <= 22'h3feff6; 
        10'b0011001000: data <= 22'h3fd2c6; 
        10'b0011001001: data <= 22'h3fcaec; 
        10'b0011001010: data <= 22'h3fdfb0; 
        10'b0011001011: data <= 22'h00042d; 
        10'b0011001100: data <= 22'h001529; 
        10'b0011001101: data <= 22'h00298d; 
        10'b0011001110: data <= 22'h002873; 
        10'b0011001111: data <= 22'h002353; 
        10'b0011010000: data <= 22'h000a39; 
        10'b0011010001: data <= 22'h3ffca8; 
        10'b0011010010: data <= 22'h3ff4b4; 
        10'b0011010011: data <= 22'h0000c5; 
        10'b0011010100: data <= 22'h00117f; 
        10'b0011010101: data <= 22'h000fd5; 
        10'b0011010110: data <= 22'h00140b; 
        10'b0011010111: data <= 22'h002ccd; 
        10'b0011011000: data <= 22'h0026bc; 
        10'b0011011001: data <= 22'h002e52; 
        10'b0011011010: data <= 22'h0040c3; 
        10'b0011011011: data <= 22'h0056df; 
        10'b0011011100: data <= 22'h006a0f; 
        10'b0011011101: data <= 22'h004c93; 
        10'b0011011110: data <= 22'h000bcb; 
        10'b0011011111: data <= 22'h3ffe2e; 
        10'b0011100000: data <= 22'h3ffcfa; 
        10'b0011100001: data <= 22'h0002cc; 
        10'b0011100010: data <= 22'h3fffc0; 
        10'b0011100011: data <= 22'h3fea26; 
        10'b0011100100: data <= 22'h3fbedd; 
        10'b0011100101: data <= 22'h3fc84e; 
        10'b0011100110: data <= 22'h3fd7b3; 
        10'b0011100111: data <= 22'h00027f; 
        10'b0011101000: data <= 22'h001f80; 
        10'b0011101001: data <= 22'h000941; 
        10'b0011101010: data <= 22'h0010ee; 
        10'b0011101011: data <= 22'h0020dc; 
        10'b0011101100: data <= 22'h001409; 
        10'b0011101101: data <= 22'h3fe974; 
        10'b0011101110: data <= 22'h3fce8f; 
        10'b0011101111: data <= 22'h3fe20d; 
        10'b0011110000: data <= 22'h3feda1; 
        10'b0011110001: data <= 22'h0001c2; 
        10'b0011110010: data <= 22'h00050a; 
        10'b0011110011: data <= 22'h002556; 
        10'b0011110100: data <= 22'h002767; 
        10'b0011110101: data <= 22'h003824; 
        10'b0011110110: data <= 22'h0058bb; 
        10'b0011110111: data <= 22'h00741b; 
        10'b0011111000: data <= 22'h009ae4; 
        10'b0011111001: data <= 22'h006412; 
        10'b0011111010: data <= 22'h00123b; 
        10'b0011111011: data <= 22'h3ffe23; 
        10'b0011111100: data <= 22'h3ff32d; 
        10'b0011111101: data <= 22'h3ff87d; 
        10'b0011111110: data <= 22'h3ff201; 
        10'b0011111111: data <= 22'h3fe195; 
        10'b0100000000: data <= 22'h3fdd0e; 
        10'b0100000001: data <= 22'h3fdfb6; 
        10'b0100000010: data <= 22'h0003ed; 
        10'b0100000011: data <= 22'h3ffdbe; 
        10'b0100000100: data <= 22'h001ae1; 
        10'b0100000101: data <= 22'h001759; 
        10'b0100000110: data <= 22'h00196a; 
        10'b0100000111: data <= 22'h0043cf; 
        10'b0100001000: data <= 22'h002bbc; 
        10'b0100001001: data <= 22'h3fedde; 
        10'b0100001010: data <= 22'h3fc468; 
        10'b0100001011: data <= 22'h3faa92; 
        10'b0100001100: data <= 22'h3fb033; 
        10'b0100001101: data <= 22'h3fd190; 
        10'b0100001110: data <= 22'h3ff55b; 
        10'b0100001111: data <= 22'h3fffb5; 
        10'b0100010000: data <= 22'h002447; 
        10'b0100010001: data <= 22'h004d91; 
        10'b0100010010: data <= 22'h007040; 
        10'b0100010011: data <= 22'h00998b; 
        10'b0100010100: data <= 22'h00c0f6; 
        10'b0100010101: data <= 22'h007ec8; 
        10'b0100010110: data <= 22'h0016b4; 
        10'b0100010111: data <= 22'h3ff70e; 
        10'b0100011000: data <= 22'h3ffd40; 
        10'b0100011001: data <= 22'h3ff724; 
        10'b0100011010: data <= 22'h3ff40c; 
        10'b0100011011: data <= 22'h3ff65d; 
        10'b0100011100: data <= 22'h3ff5d0; 
        10'b0100011101: data <= 22'h3ff973; 
        10'b0100011110: data <= 22'h0015a6; 
        10'b0100011111: data <= 22'h002857; 
        10'b0100100000: data <= 22'h003ef6; 
        10'b0100100001: data <= 22'h0045af; 
        10'b0100100010: data <= 22'h00429a; 
        10'b0100100011: data <= 22'h00509b; 
        10'b0100100100: data <= 22'h004306; 
        10'b0100100101: data <= 22'h003383; 
        10'b0100100110: data <= 22'h3ff4f6; 
        10'b0100100111: data <= 22'h3fd5e6; 
        10'b0100101000: data <= 22'h3fb9bb; 
        10'b0100101001: data <= 22'h3fbbf7; 
        10'b0100101010: data <= 22'h3fb991; 
        10'b0100101011: data <= 22'h3fafb3; 
        10'b0100101100: data <= 22'h3fc907; 
        10'b0100101101: data <= 22'h3feeed; 
        10'b0100101110: data <= 22'h000958; 
        10'b0100101111: data <= 22'h003386; 
        10'b0100110000: data <= 22'h0066d2; 
        10'b0100110001: data <= 22'h004d48; 
        10'b0100110010: data <= 22'h001a4a; 
        10'b0100110011: data <= 22'h3ff718; 
        10'b0100110100: data <= 22'h3ff3f7; 
        10'b0100110101: data <= 22'h000016; 
        10'b0100110110: data <= 22'h3ff633; 
        10'b0100110111: data <= 22'h3ff994; 
        10'b0100111000: data <= 22'h3ff60d; 
        10'b0100111001: data <= 22'h3ffe97; 
        10'b0100111010: data <= 22'h002267; 
        10'b0100111011: data <= 22'h0029fd; 
        10'b0100111100: data <= 22'h003cb7; 
        10'b0100111101: data <= 22'h003814; 
        10'b0100111110: data <= 22'h00290d; 
        10'b0100111111: data <= 22'h002d39; 
        10'b0101000000: data <= 22'h004ad5; 
        10'b0101000001: data <= 22'h0045e5; 
        10'b0101000010: data <= 22'h00011e; 
        10'b0101000011: data <= 22'h3fd477; 
        10'b0101000100: data <= 22'h3fca06; 
        10'b0101000101: data <= 22'h3fc5dc; 
        10'b0101000110: data <= 22'h3fb268; 
        10'b0101000111: data <= 22'h3f93bc; 
        10'b0101001000: data <= 22'h3f62d2; 
        10'b0101001001: data <= 22'h3f6fb2; 
        10'b0101001010: data <= 22'h3f89be; 
        10'b0101001011: data <= 22'h3fa9c3; 
        10'b0101001100: data <= 22'h3fe150; 
        10'b0101001101: data <= 22'h000360; 
        10'b0101001110: data <= 22'h0008a6; 
        10'b0101001111: data <= 22'h3ffac5; 
        10'b0101010000: data <= 22'h3ffa9b; 
        10'b0101010001: data <= 22'h3ffb8d; 
        10'b0101010010: data <= 22'h3ff984; 
        10'b0101010011: data <= 22'h3ff6f2; 
        10'b0101010100: data <= 22'h3ff920; 
        10'b0101010101: data <= 22'h00116b; 
        10'b0101010110: data <= 22'h002779; 
        10'b0101010111: data <= 22'h002339; 
        10'b0101011000: data <= 22'h0019e4; 
        10'b0101011001: data <= 22'h000ed3; 
        10'b0101011010: data <= 22'h002bbc; 
        10'b0101011011: data <= 22'h005a8b; 
        10'b0101011100: data <= 22'h005493; 
        10'b0101011101: data <= 22'h0056b2; 
        10'b0101011110: data <= 22'h0008f0; 
        10'b0101011111: data <= 22'h3fd407; 
        10'b0101100000: data <= 22'h3fae38; 
        10'b0101100001: data <= 22'h3fbdcd; 
        10'b0101100010: data <= 22'h3fd314; 
        10'b0101100011: data <= 22'h3fbf83; 
        10'b0101100100: data <= 22'h3fb688; 
        10'b0101100101: data <= 22'h3f860b; 
        10'b0101100110: data <= 22'h3f74dc; 
        10'b0101100111: data <= 22'h3f871d; 
        10'b0101101000: data <= 22'h3faf2a; 
        10'b0101101001: data <= 22'h3fe90d; 
        10'b0101101010: data <= 22'h000131; 
        10'b0101101011: data <= 22'h3fffed; 
        10'b0101101100: data <= 22'h3ffb32; 
        10'b0101101101: data <= 22'h3ff490; 
        10'b0101101110: data <= 22'h3ff3d2; 
        10'b0101101111: data <= 22'h3ff783; 
        10'b0101110000: data <= 22'h3ffd6a; 
        10'b0101110001: data <= 22'h00091f; 
        10'b0101110010: data <= 22'h001a71; 
        10'b0101110011: data <= 22'h001364; 
        10'b0101110100: data <= 22'h00166a; 
        10'b0101110101: data <= 22'h001284; 
        10'b0101110110: data <= 22'h003ce7; 
        10'b0101110111: data <= 22'h00440f; 
        10'b0101111000: data <= 22'h0032a0; 
        10'b0101111001: data <= 22'h002f4b; 
        10'b0101111010: data <= 22'h3ff680; 
        10'b0101111011: data <= 22'h3fcba7; 
        10'b0101111100: data <= 22'h3faacf; 
        10'b0101111101: data <= 22'h3fd2fd; 
        10'b0101111110: data <= 22'h3ff005; 
        10'b0101111111: data <= 22'h3fed80; 
        10'b0110000000: data <= 22'h3ff730; 
        10'b0110000001: data <= 22'h3fdd74; 
        10'b0110000010: data <= 22'h3fc18a; 
        10'b0110000011: data <= 22'h3fa4b9; 
        10'b0110000100: data <= 22'h3fbb42; 
        10'b0110000101: data <= 22'h3ff412; 
        10'b0110000110: data <= 22'h3ff303; 
        10'b0110000111: data <= 22'h3ffe1b; 
        10'b0110001000: data <= 22'h3ffb62; 
        10'b0110001001: data <= 22'h3ff39e; 
        10'b0110001010: data <= 22'h3ff9e3; 
        10'b0110001011: data <= 22'h3ff0aa; 
        10'b0110001100: data <= 22'h3ffada; 
        10'b0110001101: data <= 22'h3ffa6f; 
        10'b0110001110: data <= 22'h3fffb8; 
        10'b0110001111: data <= 22'h3ffd12; 
        10'b0110010000: data <= 22'h001bff; 
        10'b0110010001: data <= 22'h002c49; 
        10'b0110010010: data <= 22'h003522; 
        10'b0110010011: data <= 22'h000a2b; 
        10'b0110010100: data <= 22'h0011fa; 
        10'b0110010101: data <= 22'h3ffcac; 
        10'b0110010110: data <= 22'h3fd9fc; 
        10'b0110010111: data <= 22'h3fd439; 
        10'b0110011000: data <= 22'h3fc33d; 
        10'b0110011001: data <= 22'h3fca48; 
        10'b0110011010: data <= 22'h3fcdab; 
        10'b0110011011: data <= 22'h3fe7bb; 
        10'b0110011100: data <= 22'h3feafe; 
        10'b0110011101: data <= 22'h3fecec; 
        10'b0110011110: data <= 22'h3ff46d; 
        10'b0110011111: data <= 22'h3fcddc; 
        10'b0110100000: data <= 22'h3fde40; 
        10'b0110100001: data <= 22'h3fef15; 
        10'b0110100010: data <= 22'h3ff9fc; 
        10'b0110100011: data <= 22'h3ff108; 
        10'b0110100100: data <= 22'h3ff295; 
        10'b0110100101: data <= 22'h00020f; 
        10'b0110100110: data <= 22'h3ff18d; 
        10'b0110100111: data <= 22'h3ffa18; 
        10'b0110101000: data <= 22'h3fea8e; 
        10'b0110101001: data <= 22'h3fdfc8; 
        10'b0110101010: data <= 22'h3fd2e8; 
        10'b0110101011: data <= 22'h3fe220; 
        10'b0110101100: data <= 22'h000ade; 
        10'b0110101101: data <= 22'h0031e0; 
        10'b0110101110: data <= 22'h0017b0; 
        10'b0110101111: data <= 22'h0015d7; 
        10'b0110110000: data <= 22'h0012d4; 
        10'b0110110001: data <= 22'h3feefa; 
        10'b0110110010: data <= 22'h3fc793; 
        10'b0110110011: data <= 22'h3fbf19; 
        10'b0110110100: data <= 22'h3fc56e; 
        10'b0110110101: data <= 22'h3fc3fa; 
        10'b0110110110: data <= 22'h3fd5bb; 
        10'b0110110111: data <= 22'h3ffddd; 
        10'b0110111000: data <= 22'h3ff1a4; 
        10'b0110111001: data <= 22'h3ff3e1; 
        10'b0110111010: data <= 22'h3ff17c; 
        10'b0110111011: data <= 22'h3fef51; 
        10'b0110111100: data <= 22'h3ff44b; 
        10'b0110111101: data <= 22'h3fffa4; 
        10'b0110111110: data <= 22'h000253; 
        10'b0110111111: data <= 22'h3ff705; 
        10'b0111000000: data <= 22'h3ff7ed; 
        10'b0111000001: data <= 22'h3ffac2; 
        10'b0111000010: data <= 22'h3ffc80; 
        10'b0111000011: data <= 22'h3ff197; 
        10'b0111000100: data <= 22'h3ff79c; 
        10'b0111000101: data <= 22'h3fdb5c; 
        10'b0111000110: data <= 22'h3fb699; 
        10'b0111000111: data <= 22'h3fa932; 
        10'b0111001000: data <= 22'h3fc54b; 
        10'b0111001001: data <= 22'h3fdf85; 
        10'b0111001010: data <= 22'h3ff31c; 
        10'b0111001011: data <= 22'h3fed76; 
        10'b0111001100: data <= 22'h3ff3e7; 
        10'b0111001101: data <= 22'h3fd7fe; 
        10'b0111001110: data <= 22'h3fb2f2; 
        10'b0111001111: data <= 22'h3fc16f; 
        10'b0111010000: data <= 22'h3fd28c; 
        10'b0111010001: data <= 22'h3fefa0; 
        10'b0111010010: data <= 22'h3ff098; 
        10'b0111010011: data <= 22'h00027e; 
        10'b0111010100: data <= 22'h000cab; 
        10'b0111010101: data <= 22'h000202; 
        10'b0111010110: data <= 22'h000dc2; 
        10'b0111010111: data <= 22'h000321; 
        10'b0111011000: data <= 22'h000226; 
        10'b0111011001: data <= 22'h0001f0; 
        10'b0111011010: data <= 22'h3ff75f; 
        10'b0111011011: data <= 22'h3ff809; 
        10'b0111011100: data <= 22'h3ff66f; 
        10'b0111011101: data <= 22'h3fff5d; 
        10'b0111011110: data <= 22'h3ffff4; 
        10'b0111011111: data <= 22'h00010d; 
        10'b0111100000: data <= 22'h3ff6b3; 
        10'b0111100001: data <= 22'h0002ad; 
        10'b0111100010: data <= 22'h00055d; 
        10'b0111100011: data <= 22'h3fc6ad; 
        10'b0111100100: data <= 22'h3f984c; 
        10'b0111100101: data <= 22'h3f9ef3; 
        10'b0111100110: data <= 22'h3fba78; 
        10'b0111100111: data <= 22'h3fd62c; 
        10'b0111101000: data <= 22'h3fbe9c; 
        10'b0111101001: data <= 22'h3fab9d; 
        10'b0111101010: data <= 22'h3fadf6; 
        10'b0111101011: data <= 22'h3fdaa4; 
        10'b0111101100: data <= 22'h3fef95; 
        10'b0111101101: data <= 22'h0018cc; 
        10'b0111101110: data <= 22'h0025ea; 
        10'b0111101111: data <= 22'h0018c6; 
        10'b0111110000: data <= 22'h0018ff; 
        10'b0111110001: data <= 22'h000743; 
        10'b0111110010: data <= 22'h0000d0; 
        10'b0111110011: data <= 22'h000dce; 
        10'b0111110100: data <= 22'h000e08; 
        10'b0111110101: data <= 22'h3ff42b; 
        10'b0111110110: data <= 22'h3fff85; 
        10'b0111110111: data <= 22'h000054; 
        10'b0111111000: data <= 22'h000165; 
        10'b0111111001: data <= 22'h3ff5ef; 
        10'b0111111010: data <= 22'h3ff9a4; 
        10'b0111111011: data <= 22'h3ff7d2; 
        10'b0111111100: data <= 22'h001485; 
        10'b0111111101: data <= 22'h001b1d; 
        10'b0111111110: data <= 22'h00406a; 
        10'b0111111111: data <= 22'h000b54; 
        10'b1000000000: data <= 22'h3fc1fb; 
        10'b1000000001: data <= 22'h3fa5bc; 
        10'b1000000010: data <= 22'h3f8938; 
        10'b1000000011: data <= 22'h3f95e8; 
        10'b1000000100: data <= 22'h3fb3eb; 
        10'b1000000101: data <= 22'h3fd48d; 
        10'b1000000110: data <= 22'h3fea50; 
        10'b1000000111: data <= 22'h3ff6eb; 
        10'b1000001000: data <= 22'h3ffe5f; 
        10'b1000001001: data <= 22'h001d1e; 
        10'b1000001010: data <= 22'h000ea4; 
        10'b1000001011: data <= 22'h0019f8; 
        10'b1000001100: data <= 22'h001175; 
        10'b1000001101: data <= 22'h001954; 
        10'b1000001110: data <= 22'h0014df; 
        10'b1000001111: data <= 22'h001cdb; 
        10'b1000010000: data <= 22'h000efd; 
        10'b1000010001: data <= 22'h00011e; 
        10'b1000010010: data <= 22'h3ff508; 
        10'b1000010011: data <= 22'h3ffc7a; 
        10'b1000010100: data <= 22'h000011; 
        10'b1000010101: data <= 22'h3ff5d9; 
        10'b1000010110: data <= 22'h3ffa8f; 
        10'b1000010111: data <= 22'h00022d; 
        10'b1000011000: data <= 22'h001f24; 
        10'b1000011001: data <= 22'h003534; 
        10'b1000011010: data <= 22'h0047a2; 
        10'b1000011011: data <= 22'h003038; 
        10'b1000011100: data <= 22'h001e8b; 
        10'b1000011101: data <= 22'h0009ea; 
        10'b1000011110: data <= 22'h3fe933; 
        10'b1000011111: data <= 22'h3fe7a8; 
        10'b1000100000: data <= 22'h00020f; 
        10'b1000100001: data <= 22'h001d30; 
        10'b1000100010: data <= 22'h000ae9; 
        10'b1000100011: data <= 22'h000f80; 
        10'b1000100100: data <= 22'h000fbc; 
        10'b1000100101: data <= 22'h3ffb0a; 
        10'b1000100110: data <= 22'h000b4b; 
        10'b1000100111: data <= 22'h000b09; 
        10'b1000101000: data <= 22'h00025a; 
        10'b1000101001: data <= 22'h0012ea; 
        10'b1000101010: data <= 22'h00207c; 
        10'b1000101011: data <= 22'h0017bf; 
        10'b1000101100: data <= 22'h0001fb; 
        10'b1000101101: data <= 22'h3fff9c; 
        10'b1000101110: data <= 22'h3fffe4; 
        10'b1000101111: data <= 22'h3ff33d; 
        10'b1000110000: data <= 22'h3fff5b; 
        10'b1000110001: data <= 22'h3ff11d; 
        10'b1000110010: data <= 22'h3ff8e8; 
        10'b1000110011: data <= 22'h3ff4e3; 
        10'b1000110100: data <= 22'h00042c; 
        10'b1000110101: data <= 22'h0022fe; 
        10'b1000110110: data <= 22'h0028a2; 
        10'b1000110111: data <= 22'h003182; 
        10'b1000111000: data <= 22'h004560; 
        10'b1000111001: data <= 22'h003a97; 
        10'b1000111010: data <= 22'h00337a; 
        10'b1000111011: data <= 22'h004b07; 
        10'b1000111100: data <= 22'h002eb6; 
        10'b1000111101: data <= 22'h002308; 
        10'b1000111110: data <= 22'h3ff623; 
        10'b1000111111: data <= 22'h3ff6f1; 
        10'b1001000000: data <= 22'h0019d0; 
        10'b1001000001: data <= 22'h000d35; 
        10'b1001000010: data <= 22'h001591; 
        10'b1001000011: data <= 22'h001c8a; 
        10'b1001000100: data <= 22'h0018fe; 
        10'b1001000101: data <= 22'h0013a1; 
        10'b1001000110: data <= 22'h002ef0; 
        10'b1001000111: data <= 22'h002315; 
        10'b1001001000: data <= 22'h3ffb6e; 
        10'b1001001001: data <= 22'h3ff168; 
        10'b1001001010: data <= 22'h3ffad8; 
        10'b1001001011: data <= 22'h3ff6bf; 
        10'b1001001100: data <= 22'h3ff564; 
        10'b1001001101: data <= 22'h000055; 
        10'b1001001110: data <= 22'h3ff084; 
        10'b1001001111: data <= 22'h3ffa30; 
        10'b1001010000: data <= 22'h000dce; 
        10'b1001010001: data <= 22'h3ffb96; 
        10'b1001010010: data <= 22'h0010bb; 
        10'b1001010011: data <= 22'h002d49; 
        10'b1001010100: data <= 22'h004162; 
        10'b1001010101: data <= 22'h002ac4; 
        10'b1001010110: data <= 22'h002447; 
        10'b1001010111: data <= 22'h00138d; 
        10'b1001011000: data <= 22'h00194e; 
        10'b1001011001: data <= 22'h000fb9; 
        10'b1001011010: data <= 22'h00105e; 
        10'b1001011011: data <= 22'h0013f4; 
        10'b1001011100: data <= 22'h000530; 
        10'b1001011101: data <= 22'h001014; 
        10'b1001011110: data <= 22'h00083c; 
        10'b1001011111: data <= 22'h0019eb; 
        10'b1001100000: data <= 22'h001972; 
        10'b1001100001: data <= 22'h002aae; 
        10'b1001100010: data <= 22'h00347e; 
        10'b1001100011: data <= 22'h000b58; 
        10'b1001100100: data <= 22'h000073; 
        10'b1001100101: data <= 22'h3ff388; 
        10'b1001100110: data <= 22'h3ff6e7; 
        10'b1001100111: data <= 22'h3ff6f3; 
        10'b1001101000: data <= 22'h3ffced; 
        10'b1001101001: data <= 22'h3ff1d0; 
        10'b1001101010: data <= 22'h3ff8a2; 
        10'b1001101011: data <= 22'h3ff6e6; 
        10'b1001101100: data <= 22'h0004fc; 
        10'b1001101101: data <= 22'h3ff902; 
        10'b1001101110: data <= 22'h3ff0ae; 
        10'b1001101111: data <= 22'h3ffd45; 
        10'b1001110000: data <= 22'h00196a; 
        10'b1001110001: data <= 22'h002527; 
        10'b1001110010: data <= 22'h000672; 
        10'b1001110011: data <= 22'h0020e5; 
        10'b1001110100: data <= 22'h003533; 
        10'b1001110101: data <= 22'h0041b0; 
        10'b1001110110: data <= 22'h002171; 
        10'b1001110111: data <= 22'h00050b; 
        10'b1001111000: data <= 22'h0003b1; 
        10'b1001111001: data <= 22'h000833; 
        10'b1001111010: data <= 22'h001137; 
        10'b1001111011: data <= 22'h001120; 
        10'b1001111100: data <= 22'h001d57; 
        10'b1001111101: data <= 22'h001a82; 
        10'b1001111110: data <= 22'h001baf; 
        10'b1001111111: data <= 22'h0009bd; 
        10'b1010000000: data <= 22'h3ffe93; 
        10'b1010000001: data <= 22'h00018d; 
        10'b1010000010: data <= 22'h3ffaa5; 
        10'b1010000011: data <= 22'h3ffc6a; 
        10'b1010000100: data <= 22'h3ff450; 
        10'b1010000101: data <= 22'h3ffa4b; 
        10'b1010000110: data <= 22'h3ffcb1; 
        10'b1010000111: data <= 22'h3ffb71; 
        10'b1010001000: data <= 22'h3ff4e8; 
        10'b1010001001: data <= 22'h3ff8ae; 
        10'b1010001010: data <= 22'h3fe9c1; 
        10'b1010001011: data <= 22'h3ff5e1; 
        10'b1010001100: data <= 22'h001420; 
        10'b1010001101: data <= 22'h0013b4; 
        10'b1010001110: data <= 22'h0013a9; 
        10'b1010001111: data <= 22'h00230f; 
        10'b1010010000: data <= 22'h0021a7; 
        10'b1010010001: data <= 22'h00170a; 
        10'b1010010010: data <= 22'h001a7a; 
        10'b1010010011: data <= 22'h00183f; 
        10'b1010010100: data <= 22'h0017b8; 
        10'b1010010101: data <= 22'h000ae8; 
        10'b1010010110: data <= 22'h3ff379; 
        10'b1010010111: data <= 22'h3ffe3f; 
        10'b1010011000: data <= 22'h000ba0; 
        10'b1010011001: data <= 22'h0004b8; 
        10'b1010011010: data <= 22'h000f93; 
        10'b1010011011: data <= 22'h3ff640; 
        10'b1010011100: data <= 22'h00029c; 
        10'b1010011101: data <= 22'h3ff806; 
        10'b1010011110: data <= 22'h3ff7d9; 
        10'b1010011111: data <= 22'h00026f; 
        10'b1010100000: data <= 22'h3ffee2; 
        10'b1010100001: data <= 22'h3ff857; 
        10'b1010100010: data <= 22'h3ff72d; 
        10'b1010100011: data <= 22'h0002ba; 
        10'b1010100100: data <= 22'h3ff0c6; 
        10'b1010100101: data <= 22'h3fefd5; 
        10'b1010100110: data <= 22'h3ffa30; 
        10'b1010100111: data <= 22'h3ffd0d; 
        10'b1010101000: data <= 22'h3fff18; 
        10'b1010101001: data <= 22'h001a0a; 
        10'b1010101010: data <= 22'h0021cc; 
        10'b1010101011: data <= 22'h001a03; 
        10'b1010101100: data <= 22'h0010e4; 
        10'b1010101101: data <= 22'h001784; 
        10'b1010101110: data <= 22'h002b61; 
        10'b1010101111: data <= 22'h0023e3; 
        10'b1010110000: data <= 22'h001568; 
        10'b1010110001: data <= 22'h000a69; 
        10'b1010110010: data <= 22'h0013e0; 
        10'b1010110011: data <= 22'h000ce2; 
        10'b1010110100: data <= 22'h3fff42; 
        10'b1010110101: data <= 22'h3ffe24; 
        10'b1010110110: data <= 22'h3ffb48; 
        10'b1010110111: data <= 22'h0000d1; 
        10'b1010111000: data <= 22'h3ff585; 
        10'b1010111001: data <= 22'h3ffc3c; 
        10'b1010111010: data <= 22'h000192; 
        10'b1010111011: data <= 22'h3ff32e; 
        10'b1010111100: data <= 22'h3ffa43; 
        10'b1010111101: data <= 22'h00008a; 
        10'b1010111110: data <= 22'h000183; 
        10'b1010111111: data <= 22'h3ff28d; 
        10'b1011000000: data <= 22'h3fffe8; 
        10'b1011000001: data <= 22'h3ffbd7; 
        10'b1011000010: data <= 22'h3ff006; 
        10'b1011000011: data <= 22'h3ffa1a; 
        10'b1011000100: data <= 22'h3ff1a9; 
        10'b1011000101: data <= 22'h000876; 
        10'b1011000110: data <= 22'h00064e; 
        10'b1011000111: data <= 22'h00119a; 
        10'b1011001000: data <= 22'h001183; 
        10'b1011001001: data <= 22'h001eb4; 
        10'b1011001010: data <= 22'h0001af; 
        10'b1011001011: data <= 22'h000924; 
        10'b1011001100: data <= 22'h0007b9; 
        10'b1011001101: data <= 22'h000f09; 
        10'b1011001110: data <= 22'h3ff5ee; 
        10'b1011001111: data <= 22'h3fff8f; 
        10'b1011010000: data <= 22'h3fef3b; 
        10'b1011010001: data <= 22'h000171; 
        10'b1011010010: data <= 22'h3ff9bf; 
        10'b1011010011: data <= 22'h3ff4be; 
        10'b1011010100: data <= 22'h3ffeab; 
        10'b1011010101: data <= 22'h0000c4; 
        10'b1011010110: data <= 22'h3ff1b6; 
        10'b1011010111: data <= 22'h3ff874; 
        10'b1011011000: data <= 22'h3ffb88; 
        10'b1011011001: data <= 22'h3ffb13; 
        10'b1011011010: data <= 22'h3ff57f; 
        10'b1011011011: data <= 22'h3ff80a; 
        10'b1011011100: data <= 22'h3ff726; 
        10'b1011011101: data <= 22'h3ff8bd; 
        10'b1011011110: data <= 22'h3ffd64; 
        10'b1011011111: data <= 22'h3ff595; 
        10'b1011100000: data <= 22'h3ff23f; 
        10'b1011100001: data <= 22'h3ff8da; 
        10'b1011100010: data <= 22'h3ff69b; 
        10'b1011100011: data <= 22'h3ffe39; 
        10'b1011100100: data <= 22'h000047; 
        10'b1011100101: data <= 22'h3ffc66; 
        10'b1011100110: data <= 22'h3ff5fa; 
        10'b1011100111: data <= 22'h3ffae1; 
        10'b1011101000: data <= 22'h3ffdb5; 
        10'b1011101001: data <= 22'h3ff587; 
        10'b1011101010: data <= 22'h3febc8; 
        10'b1011101011: data <= 22'h3fefa2; 
        10'b1011101100: data <= 22'h3ffc8a; 
        10'b1011101101: data <= 22'h3ffc77; 
        10'b1011101110: data <= 22'h3ff6c5; 
        10'b1011101111: data <= 22'h3ffd4d; 
        10'b1011110000: data <= 22'h3ff91f; 
        10'b1011110001: data <= 22'h3ffb4d; 
        10'b1011110010: data <= 22'h3ff77e; 
        10'b1011110011: data <= 22'h3ff1b2; 
        10'b1011110100: data <= 22'h3ffcd9; 
        10'b1011110101: data <= 22'h3ffe10; 
        10'b1011110110: data <= 22'h3ffea4; 
        10'b1011110111: data <= 22'h3ffbfa; 
        10'b1011111000: data <= 22'h3ff3c9; 
        10'b1011111001: data <= 22'h3fff3d; 
        10'b1011111010: data <= 22'h3ff7c5; 
        10'b1011111011: data <= 22'h3ff6ff; 
        10'b1011111100: data <= 22'h0002f8; 
        10'b1011111101: data <= 22'h3ff767; 
        10'b1011111110: data <= 22'h3ff634; 
        10'b1011111111: data <= 22'h3ffed6; 
        10'b1100000000: data <= 22'h3ffabc; 
        10'b1100000001: data <= 22'h3ff103; 
        10'b1100000010: data <= 22'h000054; 
        10'b1100000011: data <= 22'h3ffb63; 
        10'b1100000100: data <= 22'h3ff266; 
        10'b1100000101: data <= 22'h3ff0eb; 
        10'b1100000110: data <= 22'h3ff4b8; 
        10'b1100000111: data <= 22'h3ff0b1; 
        10'b1100001000: data <= 22'h3fffc7; 
        10'b1100001001: data <= 22'h3ff790; 
        10'b1100001010: data <= 22'h0002cf; 
        10'b1100001011: data <= 22'h3ff2fc; 
        10'b1100001100: data <= 22'h3ffc16; 
        10'b1100001101: data <= 22'h3ff977; 
        10'b1100001110: data <= 22'h3ff3f5; 
        10'b1100001111: data <= 22'h3ffe1e; 
      endcase 
    end 
  end 
endgenerate 
assign dout = data; 
endmodule
