`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// WEIGHT MEMORY
// This code create bram for 1 of 10 weights strings
// and send element with input address from the string to out.
//////////////////////////////////////////////////////////////////////////////////

module ROM_weights #( 
    parameter int BITS = 24 // bit depth
)(
    input logic clk, // clock
    input logic [9:0] address, // address of current element from string
    output [BITS-1:0] dout // current element from string
);

(* rom_style = "block" *) reg [BITS-1:0] data;

always @(posedge clk)
begin
case(address)
    10'b000000000: data <= 24'hFFFF7B; 
    10'b000000001: data <= 24'h00004B; 
    10'b000000010: data <= 24'hFFFFD6; 
    10'b000000011: data <= 24'hFFFFEC; 
    10'b000000100: data <= 24'h000059; 
    10'b000000101: data <= 24'hFFFFF6; 
    10'b000000110: data <= 24'hFFFFAB; 
    10'b000000111: data <= 24'hFFFFA6; 
    10'b000001000: data <= 24'hFFFFEB; 
    10'b000001001: data <= 24'hFFFFD3; 
    10'b000001010: data <= 24'h000063; 
    10'b000001011: data <= 24'hFFFFF8; 
    10'b000001100: data <= 24'h00002D; 
    10'b000001101: data <= 24'hFFFF7E; 
    10'b000001110: data <= 24'hFFFFF8; 
    10'b000001111: data <= 24'hFFFF4E; 
    10'b000010000: data <= 24'hFFFF6C; 
    10'b000010001: data <= 24'hFFFFD8; 
    10'b000010010: data <= 24'hFFFF68; 
    10'b000010011: data <= 24'h000062; 
    10'b000010100: data <= 24'hFFFF6B; 
    10'b000010101: data <= 24'hFFFFD0; 
    10'b000010110: data <= 24'hFFFF60; 
    10'b000010111: data <= 24'hFFFFEF; 
    10'b000011000: data <= 24'h000031; 
    10'b000011001: data <= 24'hFFFFDC; 
    10'b000011010: data <= 24'hFFFFF8; 
    10'b000011011: data <= 24'hFFFFFA; 
    10'b000011100: data <= 24'h000038; 
    10'b000011101: data <= 24'h000045; 
    10'b000011110: data <= 24'h000016; 
    10'b000011111: data <= 24'hFFFF64; 
    10'b000100000: data <= 24'hFFFF5C; 
    10'b000100001: data <= 24'h000008; 
    10'b000100010: data <= 24'hFFFF7E; 
    10'b000100011: data <= 24'hFFFFDB; 
    10'b000100100: data <= 24'hFFFF9B; 
    10'b000100101: data <= 24'hFFFF49; 
    10'b000100110: data <= 24'hFFFF8B; 
    10'b000100111: data <= 24'h000009; 
    10'b000101000: data <= 24'h00006F; 
    10'b000101001: data <= 24'hFFFF67; 
    10'b000101010: data <= 24'hFFFFAD; 
    10'b000101011: data <= 24'h000030; 
    10'b000101100: data <= 24'hFFFF81; 
    10'b000101101: data <= 24'hFFFF53; 
    10'b000101110: data <= 24'h000020; 
    10'b000101111: data <= 24'h00004D; 
    10'b000110000: data <= 24'hFFFF7B; 
    10'b000110001: data <= 24'h000024; 
    10'b000110010: data <= 24'hFFFF8F; 
    10'b000110011: data <= 24'hFFFF71; 
    10'b000110100: data <= 24'hFFFFE3; 
    10'b000110101: data <= 24'h000009; 
    10'b000110110: data <= 24'hFFFFD2; 
    10'b000110111: data <= 24'h00005F; 
    10'b000111000: data <= 24'hFFFF5A; 
    10'b000111001: data <= 24'hFFFF9A; 
    10'b000111010: data <= 24'hFFFF90; 
    10'b000111011: data <= 24'h00002F; 
    10'b000111100: data <= 24'h00000C; 
    10'b000111101: data <= 24'hFFFF54; 
    10'b000111110: data <= 24'hFFFFD7; 
    10'b000111111: data <= 24'h00005B; 
    10'b001000000: data <= 24'hFFFFC8; 
    10'b001000001: data <= 24'hFFFF85; 
    10'b001000010: data <= 24'hFFFF89; 
    10'b001000011: data <= 24'hFFFF35; 
    10'b001000100: data <= 24'hFFFF28; 
    10'b001000101: data <= 24'hFFFFB5; 
    10'b001000110: data <= 24'hFFFF20; 
    10'b001000111: data <= 24'hFFFEE1; 
    10'b001001000: data <= 24'hFFFF2F; 
    10'b001001001: data <= 24'hFFFFC9; 
    10'b001001010: data <= 24'hFFFF4E; 
    10'b001001011: data <= 24'hFFFF1B; 
    10'b001001100: data <= 24'hFFFFD8; 
    10'b001001101: data <= 24'h000044; 
    10'b001001110: data <= 24'h00000C; 
    10'b001001111: data <= 24'hFFFF81; 
    10'b001010000: data <= 24'h000056; 
    10'b001010001: data <= 24'hFFFF49; 
    10'b001010010: data <= 24'hFFFFD3; 
    10'b001010011: data <= 24'h000029; 
    10'b001010100: data <= 24'hFFFF55; 
    10'b001010101: data <= 24'hFFFFD7; 
    10'b001010110: data <= 24'h000060; 
    10'b001010111: data <= 24'hFFFF5A; 
    10'b001011000: data <= 24'hFFFF89; 
    10'b001011001: data <= 24'h00004D; 
    10'b001011010: data <= 24'h00001F; 
    10'b001011011: data <= 24'h000003; 
    10'b001011100: data <= 24'h00000C; 
    10'b001011101: data <= 24'hFFFFD4; 
    10'b001011110: data <= 24'hFFFFC6; 
    10'b001011111: data <= 24'hFFFF1E; 
    10'b001100000: data <= 24'hFFFECB; 
    10'b001100001: data <= 24'hFFFF51; 
    10'b001100010: data <= 24'hFFFF0E; 
    10'b001100011: data <= 24'hFFFEEE; 
    10'b001100100: data <= 24'h00002D; 
    10'b001100101: data <= 24'h000015; 
    10'b001100110: data <= 24'hFFFECF; 
    10'b001100111: data <= 24'hFFFEFB; 
    10'b001101000: data <= 24'hFFFE8A; 
    10'b001101001: data <= 24'hFFFEF6; 
    10'b001101010: data <= 24'hFFFEBF; 
    10'b001101011: data <= 24'hFFFF21; 
    10'b001101100: data <= 24'hFFFF65; 
    10'b001101101: data <= 24'h00003A; 
    10'b001101110: data <= 24'h000038; 
    10'b001101111: data <= 24'hFFFFA7; 
    10'b001110000: data <= 24'h000016; 
    10'b001110001: data <= 24'hFFFF53; 
    10'b001110010: data <= 24'hFFFF86; 
    10'b001110011: data <= 24'hFFFF57; 
    10'b001110100: data <= 24'hFFFF41; 
    10'b001110101: data <= 24'hFFFFE7; 
    10'b001110110: data <= 24'hFFFFCC; 
    10'b001110111: data <= 24'hFFFF54; 
    10'b001111000: data <= 24'hFFFFC6; 
    10'b001111001: data <= 24'hFFFFDA; 
    10'b001111010: data <= 24'hFFFEEA; 
    10'b001111011: data <= 24'hFFFEEE; 
    10'b001111100: data <= 24'hFFFEF2; 
    10'b001111101: data <= 24'hFFFEFE; 
    10'b001111110: data <= 24'hFFFFB9; 
    10'b001111111: data <= 24'hFFFFE4; 
    10'b010000000: data <= 24'hFFFF2B; 
    10'b010000001: data <= 24'hFFFF38; 
    10'b010000010: data <= 24'hFFFF32; 
    10'b010000011: data <= 24'hFFFEE1; 
    10'b010000100: data <= 24'hFFFF8B; 
    10'b010000101: data <= 24'hFFFE8F; 
    10'b010000110: data <= 24'hFFFF70; 
    10'b010000111: data <= 24'hFFFFEB; 
    10'b010001000: data <= 24'hFFFF5F; 
    10'b010001001: data <= 24'hFFFFB7; 
    10'b010001010: data <= 24'hFFFFA1; 
    10'b010001011: data <= 24'hFFFFF0; 
    10'b010001100: data <= 24'h00002D; 
    10'b010001101: data <= 24'hFFFFAE; 
    10'b010001110: data <= 24'hFFFFFC; 
    10'b010001111: data <= 24'hFFFF68; 
    10'b010010000: data <= 24'hFFFFD6; 
    10'b010010001: data <= 24'hFFFFB6; 
    10'b010010010: data <= 24'hFFFFC9; 
    10'b010010011: data <= 24'hFFFF8D; 
    10'b010010100: data <= 24'hFFFFCC; 
    10'b010010101: data <= 24'hFFFF31; 
    10'b010010110: data <= 24'hFFFFA2; 
    10'b010010111: data <= 24'h00003C; 
    10'b010011000: data <= 24'h0000F1; 
    10'b010011001: data <= 24'h00020A; 
    10'b010011010: data <= 24'h000277; 
    10'b010011011: data <= 24'h000270; 
    10'b010011100: data <= 24'h0002BE; 
    10'b010011101: data <= 24'h0002F3; 
    10'b010011110: data <= 24'h00031F; 
    10'b010011111: data <= 24'h000119; 
    10'b010100000: data <= 24'h000032; 
    10'b010100001: data <= 24'h000082; 
    10'b010100010: data <= 24'hFFFFBF; 
    10'b010100011: data <= 24'hFFFFF6; 
    10'b010100100: data <= 24'hFFFEAA; 
    10'b010100101: data <= 24'hFFFF08; 
    10'b010100110: data <= 24'hFFFFEE; 
    10'b010100111: data <= 24'hFFFF7C; 
    10'b010101000: data <= 24'hFFFFBB; 
    10'b010101001: data <= 24'hFFFFDF; 
    10'b010101010: data <= 24'h000012; 
    10'b010101011: data <= 24'hFFFFC7; 
    10'b010101100: data <= 24'h000002; 
    10'b010101101: data <= 24'h000008; 
    10'b010101110: data <= 24'h000013; 
    10'b010101111: data <= 24'hFFFFF8; 
    10'b010110000: data <= 24'hFFFF54; 
    10'b010110001: data <= 24'hFFFEDC; 
    10'b010110010: data <= 24'h00009F; 
    10'b010110011: data <= 24'hFFFFE6; 
    10'b010110100: data <= 24'h0001B1; 
    10'b010110101: data <= 24'h00017F; 
    10'b010110110: data <= 24'h00016D; 
    10'b010110111: data <= 24'h00021F; 
    10'b010111000: data <= 24'h000296; 
    10'b010111001: data <= 24'h0003AA; 
    10'b010111010: data <= 24'h000368; 
    10'b010111011: data <= 24'h0002E8; 
    10'b010111100: data <= 24'h0002CD; 
    10'b010111101: data <= 24'h000333; 
    10'b010111110: data <= 24'h0001D0; 
    10'b010111111: data <= 24'h0000A6; 
    10'b011000000: data <= 24'hFFFE9C; 
    10'b011000001: data <= 24'hFFFE8D; 
    10'b011000010: data <= 24'hFFFF05; 
    10'b011000011: data <= 24'h000025; 
    10'b011000100: data <= 24'h000055; 
    10'b011000101: data <= 24'h00000D; 
    10'b011000110: data <= 24'hFFFFEE; 
    10'b011000111: data <= 24'hFFFF25; 
    10'b011001000: data <= 24'hFFFEAD; 
    10'b011001001: data <= 24'hFFFFE2; 
    10'b011001010: data <= 24'hFFFF77; 
    10'b011001011: data <= 24'h000002; 
    10'b011001100: data <= 24'hFFFF61; 
    10'b011001101: data <= 24'hFFFFD1; 
    10'b011001110: data <= 24'h00001E; 
    10'b011001111: data <= 24'h000135; 
    10'b011010000: data <= 24'h000283; 
    10'b011010001: data <= 24'h000250; 
    10'b011010010: data <= 24'h0000F2; 
    10'b011010011: data <= 24'h00017A; 
    10'b011010100: data <= 24'h00021B; 
    10'b011010101: data <= 24'h0003EF; 
    10'b011010110: data <= 24'h0002E5; 
    10'b011010111: data <= 24'h000288; 
    10'b011011000: data <= 24'h000109; 
    10'b011011001: data <= 24'h0001FD; 
    10'b011011010: data <= 24'h00022F; 
    10'b011011011: data <= 24'h00011E; 
    10'b011011100: data <= 24'hFFFF26; 
    10'b011011101: data <= 24'hFFFE9B; 
    10'b011011110: data <= 24'hFFFEC0; 
    10'b011011111: data <= 24'hFFFFEC; 
    10'b011100000: data <= 24'h000060; 
    10'b011100001: data <= 24'h000023; 
    10'b011100010: data <= 24'hFFFFD6; 
    10'b011100011: data <= 24'hFFFFFE; 
    10'b011100100: data <= 24'hFFFF07; 
    10'b011100101: data <= 24'hFFFF3F; 
    10'b011100110: data <= 24'hFFFF61; 
    10'b011100111: data <= 24'hFFFF3D; 
    10'b011101000: data <= 24'hFFFF99; 
    10'b011101001: data <= 24'hFFFF93; 
    10'b011101010: data <= 24'h000131; 
    10'b011101011: data <= 24'h000141; 
    10'b011101100: data <= 24'h0000A4; 
    10'b011101101: data <= 24'h000045; 
    10'b011101110: data <= 24'h000072; 
    10'b011101111: data <= 24'h0001C5; 
    10'b011110000: data <= 24'h000529; 
    10'b011110001: data <= 24'h00041B; 
    10'b011110010: data <= 24'h0003D0; 
    10'b011110011: data <= 24'h000133; 
    10'b011110100: data <= 24'h000102; 
    10'b011110101: data <= 24'h0000EC; 
    10'b011110110: data <= 24'h000243; 
    10'b011110111: data <= 24'h0003F1; 
    10'b011111000: data <= 24'hFFFF90; 
    10'b011111001: data <= 24'hFFFEB0; 
    10'b011111010: data <= 24'hFFFFDE; 
    10'b011111011: data <= 24'hFFFF4F; 
    10'b011111100: data <= 24'hFFFFE4; 
    10'b011111101: data <= 24'hFFFFEF; 
    10'b011111110: data <= 24'h00001D; 
    10'b011111111: data <= 24'h000016; 
    10'b100000000: data <= 24'hFFFEC8; 
    10'b100000001: data <= 24'hFFFF21; 
    10'b100000010: data <= 24'hFFFEC1; 
    10'b100000011: data <= 24'hFFFF49; 
    10'b100000100: data <= 24'hFFFF4B; 
    10'b100000101: data <= 24'hFFFFA3; 
    10'b100000110: data <= 24'h0000DB; 
    10'b100000111: data <= 24'hFFFF44; 
    10'b100001000: data <= 24'h00006D; 
    10'b100001001: data <= 24'h00014A; 
    10'b100001010: data <= 24'h000126; 
    10'b100001011: data <= 24'h0000FA; 
    10'b100001100: data <= 24'h0002D3; 
    10'b100001101: data <= 24'h0003C4; 
    10'b100001110: data <= 24'h000454; 
    10'b100001111: data <= 24'h000281; 
    10'b100010000: data <= 24'h0000C3; 
    10'b100010001: data <= 24'hFFFFDB; 
    10'b100010010: data <= 24'h0001DB; 
    10'b100010011: data <= 24'h000402; 
    10'b100010100: data <= 24'h00012B; 
    10'b100010101: data <= 24'hFFFF03; 
    10'b100010110: data <= 24'h000003; 
    10'b100010111: data <= 24'hFFFFE0; 
    10'b100011000: data <= 24'hFFFF5D; 
    10'b100011001: data <= 24'h00004F; 
    10'b100011010: data <= 24'hFFFF77; 
    10'b100011011: data <= 24'hFFFF07; 
    10'b100011100: data <= 24'hFFFF1C; 
    10'b100011101: data <= 24'hFFFF4B; 
    10'b100011110: data <= 24'hFFFF67; 
    10'b100011111: data <= 24'h000014; 
    10'b100100000: data <= 24'h000068; 
    10'b100100001: data <= 24'hFFFFE7; 
    10'b100100010: data <= 24'hFFFF51; 
    10'b100100011: data <= 24'h000038; 
    10'b100100100: data <= 24'h000047; 
    10'b100100101: data <= 24'hFFFFD6; 
    10'b100100110: data <= 24'hFFFEA3; 
    10'b100100111: data <= 24'hFFFDA9; 
    10'b100101000: data <= 24'hFFFE98; 
    10'b100101001: data <= 24'h00015B; 
    10'b100101010: data <= 24'h000372; 
    10'b100101011: data <= 24'h000392; 
    10'b100101100: data <= 24'h000328; 
    10'b100101101: data <= 24'h00024A; 
    10'b100101110: data <= 24'h000364; 
    10'b100101111: data <= 24'h0004A4; 
    10'b100110000: data <= 24'h000235; 
    10'b100110001: data <= 24'hFFFF16; 
    10'b100110010: data <= 24'hFFFF15; 
    10'b100110011: data <= 24'hFFFF4D; 
    10'b100110100: data <= 24'hFFFF86; 
    10'b100110101: data <= 24'hFFFF5D; 
    10'b100110110: data <= 24'h000044; 
    10'b100110111: data <= 24'hFFFFCD; 
    10'b100111000: data <= 24'hFFFE42; 
    10'b100111001: data <= 24'hFFFFA0; 
    10'b100111010: data <= 24'h000045; 
    10'b100111011: data <= 24'h000150; 
    10'b100111100: data <= 24'h0000FC; 
    10'b100111101: data <= 24'hFFFF9F; 
    10'b100111110: data <= 24'h000058; 
    10'b100111111: data <= 24'h000008; 
    10'b101000000: data <= 24'h0000AD; 
    10'b101000001: data <= 24'hFFFF89; 
    10'b101000010: data <= 24'hFFFC4E; 
    10'b101000011: data <= 24'hFFF929; 
    10'b101000100: data <= 24'hFFF990; 
    10'b101000101: data <= 24'hFFFD7C; 
    10'b101000110: data <= 24'hFFFFAA; 
    10'b101000111: data <= 24'h0001D0; 
    10'b101001000: data <= 24'h0002E7; 
    10'b101001001: data <= 24'h0002B0; 
    10'b101001010: data <= 24'h0003AB; 
    10'b101001011: data <= 24'h000429; 
    10'b101001100: data <= 24'h0002FE; 
    10'b101001101: data <= 24'hFFFF6C; 
    10'b101001110: data <= 24'hFFFFF6; 
    10'b101001111: data <= 24'hFFFF42; 
    10'b101010000: data <= 24'hFFFF80; 
    10'b101010001: data <= 24'hFFFFD7; 
    10'b101010010: data <= 24'hFFFFC5; 
    10'b101010011: data <= 24'hFFFFCF; 
    10'b101010100: data <= 24'hFFFF04; 
    10'b101010101: data <= 24'h000028; 
    10'b101010110: data <= 24'h00016E; 
    10'b101010111: data <= 24'h00017F; 
    10'b101011000: data <= 24'h0000B9; 
    10'b101011001: data <= 24'hFFFFCC; 
    10'b101011010: data <= 24'h000106; 
    10'b101011011: data <= 24'h0000BA; 
    10'b101011100: data <= 24'h000157; 
    10'b101011101: data <= 24'hFFFEE5; 
    10'b101011110: data <= 24'hFFF8C1; 
    10'b101011111: data <= 24'hFFF706; 
    10'b101100000: data <= 24'hFFF710; 
    10'b101100001: data <= 24'hFFFB1D; 
    10'b101100010: data <= 24'hFFFF22; 
    10'b101100011: data <= 24'hFFFFA4; 
    10'b101100100: data <= 24'h000070; 
    10'b101100101: data <= 24'h000140; 
    10'b101100110: data <= 24'h0004C2; 
    10'b101100111: data <= 24'h00045A; 
    10'b101101000: data <= 24'h000306; 
    10'b101101001: data <= 24'h00001B; 
    10'b101101010: data <= 24'hFFFF86; 
    10'b101101011: data <= 24'hFFFF84; 
    10'b101101100: data <= 24'hFFFF4A; 
    10'b101101101: data <= 24'hFFFFFB; 
    10'b101101110: data <= 24'h00003F; 
    10'b101101111: data <= 24'hFFFF52; 
    10'b101110000: data <= 24'hFFFFBD; 
    10'b101110001: data <= 24'h0000E3; 
    10'b101110010: data <= 24'h0001BC; 
    10'b101110011: data <= 24'h00023D; 
    10'b101110100: data <= 24'h0001B1; 
    10'b101110101: data <= 24'h00012F; 
    10'b101110110: data <= 24'h00019E; 
    10'b101110111: data <= 24'h000142; 
    10'b101111000: data <= 24'h0000E8; 
    10'b101111001: data <= 24'hFFFB96; 
    10'b101111010: data <= 24'hFFF8BE; 
    10'b101111011: data <= 24'hFFF6C7; 
    10'b101111100: data <= 24'hFFF86D; 
    10'b101111101: data <= 24'hFFFC3D; 
    10'b101111110: data <= 24'hFFFE29; 
    10'b101111111: data <= 24'hFFFD88; 
    10'b110000000: data <= 24'hFFFE1D; 
    10'b110000001: data <= 24'h0000D3; 
    10'b110000010: data <= 24'h00031F; 
    10'b110000011: data <= 24'h0004E6; 
    10'b110000100: data <= 24'h0002C8; 
    10'b110000101: data <= 24'h000072; 
    10'b110000110: data <= 24'h000000; 
    10'b110000111: data <= 24'h000045; 
    10'b110001000: data <= 24'hFFFFE6; 
    10'b110001001: data <= 24'h000036; 
    10'b110001010: data <= 24'hFFFF74; 
    10'b110001011: data <= 24'hFFFF9B; 
    10'b110001100: data <= 24'hFFFF27; 
    10'b110001101: data <= 24'h00024A; 
    10'b110001110: data <= 24'h0002FA; 
    10'b110001111: data <= 24'h00039D; 
    10'b110010000: data <= 24'h0001BC; 
    10'b110010001: data <= 24'h000215; 
    10'b110010010: data <= 24'h000310; 
    10'b110010011: data <= 24'h0001C2; 
    10'b110010100: data <= 24'h00006E; 
    10'b110010101: data <= 24'hFFFC29; 
    10'b110010110: data <= 24'hFFF771; 
    10'b110010111: data <= 24'hFFF6C0; 
    10'b110011000: data <= 24'hFFF8A4; 
    10'b110011001: data <= 24'hFFFBF9; 
    10'b110011010: data <= 24'hFFFE3A; 
    10'b110011011: data <= 24'hFFFDDB; 
    10'b110011100: data <= 24'h000031; 
    10'b110011101: data <= 24'h0001BE; 
    10'b110011110: data <= 24'h000214; 
    10'b110011111: data <= 24'h0004F3; 
    10'b110100000: data <= 24'h000293; 
    10'b110100001: data <= 24'hFFFF7A; 
    10'b110100010: data <= 24'hFFFFBD; 
    10'b110100011: data <= 24'hFFFF71; 
    10'b110100100: data <= 24'h000049; 
    10'b110100101: data <= 24'h000028; 
    10'b110100110: data <= 24'hFFFF87; 
    10'b110100111: data <= 24'hFFFFE4; 
    10'b110101000: data <= 24'hFFFFF6; 
    10'b110101001: data <= 24'h00033C; 
    10'b110101010: data <= 24'h000259; 
    10'b110101011: data <= 24'h00033B; 
    10'b110101100: data <= 24'h00023B; 
    10'b110101101: data <= 24'h0002F5; 
    10'b110101110: data <= 24'h0003BD; 
    10'b110101111: data <= 24'h000108; 
    10'b110110000: data <= 24'hFFFD2E; 
    10'b110110001: data <= 24'hFFF8D1; 
    10'b110110010: data <= 24'hFFF669; 
    10'b110110011: data <= 24'hFFF6DE; 
    10'b110110100: data <= 24'hFFF9D5; 
    10'b110110101: data <= 24'hFFFCFD; 
    10'b110110110: data <= 24'hFFFEE0; 
    10'b110110111: data <= 24'hFFFEE9; 
    10'b110111000: data <= 24'h0000EF; 
    10'b110111001: data <= 24'h0000D2; 
    10'b110111010: data <= 24'h000325; 
    10'b110111011: data <= 24'h0003B2; 
    10'b110111100: data <= 24'h0001EA; 
    10'b110111101: data <= 24'hFFFFCF; 
    10'b110111110: data <= 24'h00000D; 
    10'b110111111: data <= 24'hFFFF7E; 
    10'b111000000: data <= 24'h000015; 
    10'b111000001: data <= 24'h00005C; 
    10'b111000010: data <= 24'hFFFF44; 
    10'b111000011: data <= 24'hFFFF9A; 
    10'b111000100: data <= 24'h00008B; 
    10'b111000101: data <= 24'h0002EF; 
    10'b111000110: data <= 24'h0003A6; 
    10'b111000111: data <= 24'h0002D2; 
    10'b111001000: data <= 24'h0001F5; 
    10'b111001001: data <= 24'h0001F9; 
    10'b111001010: data <= 24'h000355; 
    10'b111001011: data <= 24'hFFFF8F; 
    10'b111001100: data <= 24'hFFFA87; 
    10'b111001101: data <= 24'hFFF67B; 
    10'b111001110: data <= 24'hFFF6BB; 
    10'b111001111: data <= 24'hFFF8A5; 
    10'b111010000: data <= 24'hFFFC0F; 
    10'b111010001: data <= 24'hFFFE29; 
    10'b111010010: data <= 24'hFFFFF9; 
    10'b111010011: data <= 24'h00009A; 
    10'b111010100: data <= 24'h000162; 
    10'b111010101: data <= 24'h00020F; 
    10'b111010110: data <= 24'h0002D5; 
    10'b111010111: data <= 24'h0002B4; 
    10'b111011000: data <= 24'h000107; 
    10'b111011001: data <= 24'h00000C; 
    10'b111011010: data <= 24'hFFFFAA; 
    10'b111011011: data <= 24'hFFFF8C; 
    10'b111011100: data <= 24'hFFFFBC; 
    10'b111011101: data <= 24'h000016; 
    10'b111011110: data <= 24'hFFFF61; 
    10'b111011111: data <= 24'hFFFECB; 
    10'b111100000: data <= 24'h00001A; 
    10'b111100001: data <= 24'h000216; 
    10'b111100010: data <= 24'h00029E; 
    10'b111100011: data <= 24'h00028B; 
    10'b111100100: data <= 24'h0000CB; 
    10'b111100101: data <= 24'h00020A; 
    10'b111100110: data <= 24'h00033A; 
    10'b111100111: data <= 24'hFFFF81; 
    10'b111101000: data <= 24'hFFF971; 
    10'b111101001: data <= 24'hFFF69C; 
    10'b111101010: data <= 24'hFFF7BC; 
    10'b111101011: data <= 24'hFFFB12; 
    10'b111101100: data <= 24'hFFFF5A; 
    10'b111101101: data <= 24'h000141; 
    10'b111101110: data <= 24'h0001CF; 
    10'b111101111: data <= 24'h0001AB; 
    10'b111110000: data <= 24'h000220; 
    10'b111110001: data <= 24'h00019F; 
    10'b111110010: data <= 24'h000148; 
    10'b111110011: data <= 24'h000174; 
    10'b111110100: data <= 24'hFFFFEB; 
    10'b111110101: data <= 24'hFFFFC8; 
    10'b111110110: data <= 24'h00001C; 
    10'b111110111: data <= 24'hFFFF7D; 
    10'b111111000: data <= 24'hFFFFA6; 
    10'b111111001: data <= 24'h00001D; 
    10'b111111010: data <= 24'hFFFFC1; 
    10'b111111011: data <= 24'hFFFF8A; 
    10'b111111100: data <= 24'hFFFFBF; 
    10'b111111101: data <= 24'h000154; 
    10'b111111110: data <= 24'h0002B6; 
    10'b111111111: data <= 24'h000191; 
    10'b1000000000: data <= 24'h0000F6; 
    10'b1000000001: data <= 24'h0002B2; 
    10'b1000000010: data <= 24'h00052C; 
    10'b1000000011: data <= 24'h000034; 
    10'b1000000100: data <= 24'hFFFBD2; 
    10'b1000000101: data <= 24'hFFF942; 
    10'b1000000110: data <= 24'hFFFB4D; 
    10'b1000000111: data <= 24'hFFFE91; 
    10'b1000001000: data <= 24'h000184; 
    10'b1000001001: data <= 24'h00019E; 
    10'b1000001010: data <= 24'h0001B1; 
    10'b1000001011: data <= 24'h0000E1; 
    10'b1000001100: data <= 24'h000070; 
    10'b1000001101: data <= 24'h0000BB; 
    10'b1000001110: data <= 24'h000169; 
    10'b1000001111: data <= 24'h0000E1; 
    10'b1000010000: data <= 24'hFFFFE4; 
    10'b1000010001: data <= 24'hFFFF91; 
    10'b1000010010: data <= 24'h00000D; 
    10'b1000010011: data <= 24'hFFFFC1; 
    10'b1000010100: data <= 24'hFFFFC8; 
    10'b1000010101: data <= 24'hFFFFB2; 
    10'b1000010110: data <= 24'hFFFFBA; 
    10'b1000010111: data <= 24'hFFFED3; 
    10'b1000011000: data <= 24'h000080; 
    10'b1000011001: data <= 24'h000175; 
    10'b1000011010: data <= 24'h00037C; 
    10'b1000011011: data <= 24'h00032A; 
    10'b1000011100: data <= 24'h00027A; 
    10'b1000011101: data <= 24'h000349; 
    10'b1000011110: data <= 24'h00052F; 
    10'b1000011111: data <= 24'h0003A5; 
    10'b1000100000: data <= 24'h0000C5; 
    10'b1000100001: data <= 24'hFFFE52; 
    10'b1000100010: data <= 24'hFFFF44; 
    10'b1000100011: data <= 24'hFFFF87; 
    10'b1000100100: data <= 24'h0000CA; 
    10'b1000100101: data <= 24'hFFFFA2; 
    10'b1000100110: data <= 24'hFFFF53; 
    10'b1000100111: data <= 24'hFFFF97; 
    10'b1000101000: data <= 24'h0000D0; 
    10'b1000101001: data <= 24'h0000BE; 
    10'b1000101010: data <= 24'h000174; 
    10'b1000101011: data <= 24'hFFFFCE; 
    10'b1000101100: data <= 24'h000035; 
    10'b1000101101: data <= 24'hFFFFAE; 
    10'b1000101110: data <= 24'hFFFF3F; 
    10'b1000101111: data <= 24'h000042; 
    10'b1000110000: data <= 24'h000041; 
    10'b1000110001: data <= 24'h000056; 
    10'b1000110010: data <= 24'hFFFFC1; 
    10'b1000110011: data <= 24'hFFFF71; 
    10'b1000110100: data <= 24'hFFFFAB; 
    10'b1000110101: data <= 24'h00017E; 
    10'b1000110110: data <= 24'h0002CD; 
    10'b1000110111: data <= 24'h000210; 
    10'b1000111000: data <= 24'h00028E; 
    10'b1000111001: data <= 24'h000324; 
    10'b1000111010: data <= 24'h0004E5; 
    10'b1000111011: data <= 24'h0004E4; 
    10'b1000111100: data <= 24'h000273; 
    10'b1000111101: data <= 24'h0000BF; 
    10'b1000111110: data <= 24'hFFFF7D; 
    10'b1000111111: data <= 24'h00005A; 
    10'b1001000000: data <= 24'h000055; 
    10'b1001000001: data <= 24'hFFFF49; 
    10'b1001000010: data <= 24'hFFFF75; 
    10'b1001000011: data <= 24'hFFFF3D; 
    10'b1001000100: data <= 24'h000067; 
    10'b1001000101: data <= 24'h000080; 
    10'b1001000110: data <= 24'h0000C5; 
    10'b1001000111: data <= 24'h000044; 
    10'b1001001000: data <= 24'hFFFF91; 
    10'b1001001001: data <= 24'hFFFFE6; 
    10'b1001001010: data <= 24'hFFFF64; 
    10'b1001001011: data <= 24'hFFFFAF; 
    10'b1001001100: data <= 24'hFFFF8C; 
    10'b1001001101: data <= 24'hFFFF55; 
    10'b1001001110: data <= 24'hFFFFC3; 
    10'b1001001111: data <= 24'hFFFF8F; 
    10'b1001010000: data <= 24'hFFFFB8; 
    10'b1001010001: data <= 24'h000063; 
    10'b1001010010: data <= 24'h0001BB; 
    10'b1001010011: data <= 24'h0002D0; 
    10'b1001010100: data <= 24'h0001F9; 
    10'b1001010101: data <= 24'h000224; 
    10'b1001010110: data <= 24'h000431; 
    10'b1001010111: data <= 24'h0004BD; 
    10'b1001011000: data <= 24'h000324; 
    10'b1001011001: data <= 24'h000130; 
    10'b1001011010: data <= 24'h000071; 
    10'b1001011011: data <= 24'h000017; 
    10'b1001011100: data <= 24'hFFFFEC; 
    10'b1001011101: data <= 24'hFFFEB3; 
    10'b1001011110: data <= 24'hFFFF02; 
    10'b1001011111: data <= 24'hFFFF6E; 
    10'b1001100000: data <= 24'h00007E; 
    10'b1001100001: data <= 24'hFFFFF6; 
    10'b1001100010: data <= 24'hFFFF69; 
    10'b1001100011: data <= 24'hFFFF0F; 
    10'b1001100100: data <= 24'hFFFFC4; 
    10'b1001100101: data <= 24'hFFFFB0; 
    10'b1001100110: data <= 24'hFFFF8B; 
    10'b1001100111: data <= 24'hFFFF9B; 
    10'b1001101000: data <= 24'hFFFF70; 
    10'b1001101001: data <= 24'h000008; 
    10'b1001101010: data <= 24'h00000D; 
    10'b1001101011: data <= 24'hFFFFAB; 
    10'b1001101100: data <= 24'hFFFF68; 
    10'b1001101101: data <= 24'h000037; 
    10'b1001101110: data <= 24'h000142; 
    10'b1001101111: data <= 24'h000117; 
    10'b1001110000: data <= 24'h000328; 
    10'b1001110001: data <= 24'h000291; 
    10'b1001110010: data <= 24'h0002D4; 
    10'b1001110011: data <= 24'h00035E; 
    10'b1001110100: data <= 24'h0002DF; 
    10'b1001110101: data <= 24'h0003B1; 
    10'b1001110110: data <= 24'h000199; 
    10'b1001110111: data <= 24'h0001A2; 
    10'b1001111000: data <= 24'h0000E5; 
    10'b1001111001: data <= 24'hFFFF3D; 
    10'b1001111010: data <= 24'hFFFF65; 
    10'b1001111011: data <= 24'hFFFFF4; 
    10'b1001111100: data <= 24'hFFFF25; 
    10'b1001111101: data <= 24'hFFFF1A; 
    10'b1001111110: data <= 24'hFFFF91; 
    10'b1001111111: data <= 24'hFFFF88; 
    10'b1010000000: data <= 24'hFFFFD5; 
    10'b1010000001: data <= 24'hFFFFB6; 
    10'b1010000010: data <= 24'hFFFFA0; 
    10'b1010000011: data <= 24'hFFFFCD; 
    10'b1010000100: data <= 24'hFFFF70; 
    10'b1010000101: data <= 24'hFFFFD9; 
    10'b1010000110: data <= 24'hFFFFFC; 
    10'b1010000111: data <= 24'hFFFF52; 
    10'b1010001000: data <= 24'hFFFF4E; 
    10'b1010001001: data <= 24'hFFFFCC; 
    10'b1010001010: data <= 24'hFFFFEA; 
    10'b1010001011: data <= 24'h0000DF; 
    10'b1010001100: data <= 24'h00013C; 
    10'b1010001101: data <= 24'h0002ED; 
    10'b1010001110: data <= 24'h000381; 
    10'b1010001111: data <= 24'h000449; 
    10'b1010010000: data <= 24'h00043E; 
    10'b1010010001: data <= 24'h00028B; 
    10'b1010010010: data <= 24'h000212; 
    10'b1010010011: data <= 24'h000125; 
    10'b1010010100: data <= 24'h00007B; 
    10'b1010010101: data <= 24'hFFFFF3; 
    10'b1010010110: data <= 24'hFFFE62; 
    10'b1010010111: data <= 24'hFFFDF9; 
    10'b1010011000: data <= 24'hFFFE6E; 
    10'b1010011001: data <= 24'hFFFF39; 
    10'b1010011010: data <= 24'hFFFF5E; 
    10'b1010011011: data <= 24'hFFFFEB; 
    10'b1010011100: data <= 24'hFFFFC2; 
    10'b1010011101: data <= 24'h000032; 
    10'b1010011110: data <= 24'hFFFFA9; 
    10'b1010011111: data <= 24'hFFFF4B; 
    10'b1010100000: data <= 24'hFFFFAF; 
    10'b1010100001: data <= 24'hFFFFDC; 
    10'b1010100010: data <= 24'hFFFF4E; 
    10'b1010100011: data <= 24'hFFFFF8; 
    10'b1010100100: data <= 24'hFFFFCF; 
    10'b1010100101: data <= 24'hFFFFD1; 
    10'b1010100110: data <= 24'hFFFF2A; 
    10'b1010100111: data <= 24'hFFFEE2; 
    10'b1010101000: data <= 24'hFFFF61; 
    10'b1010101001: data <= 24'hFFFF71; 
    10'b1010101010: data <= 24'h0000A5; 
    10'b1010101011: data <= 24'h00007D; 
    10'b1010101100: data <= 24'h00012F; 
    10'b1010101101: data <= 24'h0001BB; 
    10'b1010101110: data <= 24'h0000EA; 
    10'b1010101111: data <= 24'hFFFF4D; 
    10'b1010110000: data <= 24'hFFFEEB; 
    10'b1010110001: data <= 24'hFFFEB5; 
    10'b1010110010: data <= 24'hFFFEE6; 
    10'b1010110011: data <= 24'hFFFE74; 
    10'b1010110100: data <= 24'hFFFE87; 
    10'b1010110101: data <= 24'hFFFE9C; 
    10'b1010110110: data <= 24'hFFFFBA; 
    10'b1010110111: data <= 24'hFFFFA2; 
    10'b1010111000: data <= 24'hFFFF6A; 
    10'b1010111001: data <= 24'hFFFF91; 
    10'b1010111010: data <= 24'h000008; 
    10'b1010111011: data <= 24'hFFFF7E; 
    10'b1010111100: data <= 24'hFFFF93; 
    10'b1010111101: data <= 24'h000065; 
    10'b1010111110: data <= 24'hFFFFC9; 
    10'b1010111111: data <= 24'h000054; 
    10'b1011000000: data <= 24'h000060; 
    10'b1011000001: data <= 24'hFFFFFB; 
    10'b1011000010: data <= 24'hFFFF3F; 
    10'b1011000011: data <= 24'hFFFFAB; 
    10'b1011000100: data <= 24'hFFFE89; 
    10'b1011000101: data <= 24'hFFFE9D; 
    10'b1011000110: data <= 24'hFFFE46; 
    10'b1011000111: data <= 24'hFFFDC3; 
    10'b1011001000: data <= 24'hFFFD71; 
    10'b1011001001: data <= 24'hFFFDAB; 
    10'b1011001010: data <= 24'hFFFD49; 
    10'b1011001011: data <= 24'hFFFD8D; 
    10'b1011001100: data <= 24'hFFFDAF; 
    10'b1011001101: data <= 24'hFFFE9B; 
    10'b1011001110: data <= 24'hFFFED8; 
    10'b1011001111: data <= 24'hFFFF06; 
    10'b1011010000: data <= 24'hFFFEEB; 
    10'b1011010001: data <= 24'hFFFF00; 
    10'b1011010010: data <= 24'hFFFFAA; 
    10'b1011010011: data <= 24'h00005F; 
    10'b1011010100: data <= 24'h00002E; 
    10'b1011010101: data <= 24'hFFFFBB; 
    10'b1011010110: data <= 24'hFFFFA4; 
    10'b1011010111: data <= 24'hFFFFDD; 
    10'b1011011000: data <= 24'h000050; 
    10'b1011011001: data <= 24'h000048; 
    10'b1011011010: data <= 24'hFFFFB6; 
    10'b1011011011: data <= 24'h000004; 
    10'b1011011100: data <= 24'hFFFF9B; 
    10'b1011011101: data <= 24'hFFFFAF; 
    10'b1011011110: data <= 24'hFFFF52; 
    10'b1011011111: data <= 24'h000022; 
    10'b1011100000: data <= 24'hFFFFA3; 
    10'b1011100001: data <= 24'hFFFEC5; 
    10'b1011100010: data <= 24'hFFFEC4; 
    10'b1011100011: data <= 24'hFFFEE2; 
    10'b1011100100: data <= 24'hFFFF8D; 
    10'b1011100101: data <= 24'hFFFEE3; 
    10'b1011100110: data <= 24'hFFFEF1; 
    10'b1011100111: data <= 24'hFFFF9B; 
    10'b1011101000: data <= 24'hFFFEE0; 
    10'b1011101001: data <= 24'hFFFF16; 
    10'b1011101010: data <= 24'hFFFF51; 
    10'b1011101011: data <= 24'hFFFF24; 
    10'b1011101100: data <= 24'hFFFF92; 
    10'b1011101101: data <= 24'hFFFEF8; 
    10'b1011101110: data <= 24'hFFFF21; 
    10'b1011101111: data <= 24'h000056; 
    10'b1011110000: data <= 24'hFFFF77; 
    10'b1011110001: data <= 24'h000019; 
    10'b1011110010: data <= 24'h000047; 
    10'b1011110011: data <= 24'hFFFFEF; 
    10'b1011110100: data <= 24'hFFFF6B; 
    10'b1011110101: data <= 24'h00003B; 
    10'b1011110110: data <= 24'hFFFFE6; 
    10'b1011110111: data <= 24'hFFFFAF; 
    10'b1011111000: data <= 24'h00004C; 
    10'b1011111001: data <= 24'h00000E; 
    10'b1011111010: data <= 24'h00001A; 
    10'b1011111011: data <= 24'hFFFF4A; 
    10'b1011111100: data <= 24'h000059; 
    10'b1011111101: data <= 24'h000056; 
    10'b1011111110: data <= 24'h00001E; 
    10'b1011111111: data <= 24'h00003E; 
    10'b1100000000: data <= 24'hFFFFD4; 
    10'b1100000001: data <= 24'hFFFF94; 
    10'b1100000010: data <= 24'h00003B; 
    10'b1100000011: data <= 24'hFFFF63; 
    10'b1100000100: data <= 24'hFFFFC6; 
    10'b1100000101: data <= 24'hFFFF92; 
    10'b1100000110: data <= 24'hFFFFE5; 
    10'b1100000111: data <= 24'hFFFF9E; 
    10'b1100001000: data <= 24'hFFFF46; 
    10'b1100001001: data <= 24'hFFFF59; 
    10'b1100001010: data <= 24'hFFFF13; 
    10'b1100001011: data <= 24'hFFFFC9; 
    10'b1100001100: data <= 24'h000026; 
    10'b1100001101: data <= 24'hFFFF69; 
    10'b1100001110: data <= 24'hFFFF42; 
    10'b1100001111: data <= 24'h000031; 
endcase
end

assign dout = data;

endmodule
